magic
tech sky130A
magscale 1 2
timestamp 1636440888
<< metal2 >>
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< metal3 >>
rect 16194 703800 21194 704800
rect 16194 703500 16352 703800
rect 16652 703500 16852 703800
rect 17152 703500 17352 703800
rect 17652 703500 17852 703800
rect 18152 703500 18352 703800
rect 18652 703500 18852 703800
rect 19152 703500 19352 703800
rect 19652 703500 19852 703800
rect 20152 703500 20352 703800
rect 20652 703500 20852 703800
rect 21152 703500 21194 703800
rect 16194 703300 21194 703500
rect 16194 703000 16352 703300
rect 16652 703000 16852 703300
rect 17152 703000 17352 703300
rect 17652 703000 17852 703300
rect 18152 703000 18352 703300
rect 18652 703000 18852 703300
rect 19152 703000 19352 703300
rect 19652 703000 19852 703300
rect 20152 703000 20352 703300
rect 20652 703000 20852 703300
rect 21152 703000 21194 703300
rect 16194 702800 21194 703000
rect 16194 702500 16352 702800
rect 16652 702500 16852 702800
rect 17152 702500 17352 702800
rect 17652 702500 17852 702800
rect 18152 702500 18352 702800
rect 18652 702500 18852 702800
rect 19152 702500 19352 702800
rect 19652 702500 19852 702800
rect 20152 702500 20352 702800
rect 20652 702500 20852 702800
rect 21152 702500 21194 702800
rect 16194 702300 21194 702500
rect 68194 703200 73194 704800
rect 68194 703000 70300 703200
rect 70500 703000 70600 703200
rect 70800 703000 70900 703200
rect 71100 703000 73194 703200
rect 68194 702900 73194 703000
rect 68194 702700 70300 702900
rect 70500 702700 70600 702900
rect 70800 702700 70900 702900
rect 71100 702700 73194 702900
rect 68194 702600 73194 702700
rect 68194 702400 70300 702600
rect 70500 702400 70600 702600
rect 70800 702400 70900 702600
rect 71100 702400 73194 702600
rect 68194 702300 73194 702400
rect 120194 703194 125194 704800
rect 120194 702994 122179 703194
rect 122379 702994 122479 703194
rect 122679 702994 122779 703194
rect 122979 702994 125194 703194
rect 120194 702894 125194 702994
rect 120194 702694 122179 702894
rect 122379 702694 122479 702894
rect 122679 702694 122779 702894
rect 122979 702694 125194 702894
rect 120194 702594 125194 702694
rect 120194 702394 122179 702594
rect 122379 702394 122479 702594
rect 122679 702394 122779 702594
rect 122979 702394 125194 702594
rect 120194 702300 125194 702394
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703110 418394 704800
rect 413394 703040 415760 703110
rect 415830 703040 415850 703110
rect 415920 703040 415940 703110
rect 416010 703040 416030 703110
rect 416100 703040 416120 703110
rect 416190 703040 418394 703110
rect 413394 703020 418394 703040
rect 413394 702950 415760 703020
rect 415830 702950 415850 703020
rect 415920 702950 415940 703020
rect 416010 702950 416030 703020
rect 416100 702950 416120 703020
rect 416190 702950 418394 703020
rect 413394 702930 418394 702950
rect 413394 702860 415760 702930
rect 415830 702860 415850 702930
rect 415920 702860 415940 702930
rect 416010 702860 416030 702930
rect 416100 702860 416120 702930
rect 416190 702860 418394 702930
rect 413394 702840 418394 702860
rect 413394 702770 415760 702840
rect 415830 702770 415850 702840
rect 415920 702770 415940 702840
rect 416010 702770 416030 702840
rect 416100 702770 416120 702840
rect 416190 702770 418394 702840
rect 413394 702750 418394 702770
rect 413394 702680 415760 702750
rect 415830 702680 415850 702750
rect 415920 702680 415940 702750
rect 416010 702680 416030 702750
rect 416100 702680 416120 702750
rect 416190 702680 418394 702750
rect 413394 702300 418394 702680
rect 465394 703310 470394 704800
rect 465394 703240 467220 703310
rect 467290 703240 467320 703310
rect 467390 703240 467420 703310
rect 467490 703240 470394 703310
rect 465394 703220 470394 703240
rect 465394 703150 467220 703220
rect 467290 703150 467320 703220
rect 467390 703150 467420 703220
rect 467490 703150 470394 703220
rect 465394 703130 470394 703150
rect 465394 703060 467220 703130
rect 467290 703060 467320 703130
rect 467390 703060 467420 703130
rect 467490 703060 470394 703130
rect 465394 702300 470394 703060
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702870 571594 704800
rect 566594 702800 569600 702870
rect 569670 702800 569700 702870
rect 569770 702800 569800 702870
rect 569870 702800 571594 702870
rect 566594 702770 571594 702800
rect 566594 702700 569600 702770
rect 569670 702700 569700 702770
rect 569770 702700 569800 702770
rect 569870 702700 571594 702770
rect 566594 702670 571594 702700
rect 566594 702600 569600 702670
rect 569670 702600 569700 702670
rect 569770 702600 569800 702670
rect 569870 702600 571594 702670
rect 566594 702300 571594 702600
rect -800 685200 1700 685242
rect -800 684900 200 685200
rect 500 684900 700 685200
rect 1000 684900 1200 685200
rect 1500 684900 1700 685200
rect -800 684700 1700 684900
rect -800 684400 200 684700
rect 500 684400 700 684700
rect 1000 684400 1200 684700
rect 1500 684400 1700 684700
rect -800 684200 1700 684400
rect -800 683900 200 684200
rect 500 683900 700 684200
rect 1000 683900 1200 684200
rect 1500 683900 1700 684200
rect -800 683700 1700 683900
rect -800 683400 200 683700
rect 500 683400 700 683700
rect 1000 683400 1200 683700
rect 1500 683400 1700 683700
rect -800 683200 1700 683400
rect -800 682900 200 683200
rect 500 682900 700 683200
rect 1000 682900 1200 683200
rect 1500 682900 1700 683200
rect -800 682700 1700 682900
rect -800 682400 200 682700
rect 500 682400 700 682700
rect 1000 682400 1200 682700
rect 1500 682400 1700 682700
rect -800 682200 1700 682400
rect -800 681900 200 682200
rect 500 681900 700 682200
rect 1000 681900 1200 682200
rect 1500 681900 1700 682200
rect -800 681700 1700 681900
rect -800 681400 200 681700
rect 500 681400 700 681700
rect 1000 681400 1200 681700
rect 1500 681400 1700 681700
rect -800 681200 1700 681400
rect -800 680900 200 681200
rect 500 680900 700 681200
rect 1000 680900 1200 681200
rect 1500 680900 1700 681200
rect -800 680700 1700 680900
rect -800 680400 200 680700
rect 500 680400 700 680700
rect 1000 680400 1200 680700
rect 1500 680400 1700 680700
rect -800 680242 1700 680400
rect 110760 683700 155960 694890
rect 110760 683460 110890 683700
rect 111130 683460 111220 683700
rect 111460 683460 111550 683700
rect 111790 683460 111880 683700
rect 112120 683460 112210 683700
rect 112450 683460 112540 683700
rect 112780 683460 112870 683700
rect 113110 683460 113200 683700
rect 113440 683460 113530 683700
rect 113770 683460 113860 683700
rect 114100 683460 114190 683700
rect 114430 683460 114520 683700
rect 114760 683460 114850 683700
rect 115090 683460 115180 683700
rect 115420 683460 115510 683700
rect 115750 683460 115840 683700
rect 116080 683460 116170 683700
rect 116410 683460 116500 683700
rect 116740 683460 116830 683700
rect 117070 683460 117160 683700
rect 117400 683460 117490 683700
rect 117730 683460 117820 683700
rect 118060 683460 118150 683700
rect 118390 683460 118480 683700
rect 118720 683460 118810 683700
rect 119050 683460 119140 683700
rect 119380 683460 119470 683700
rect 119710 683460 119800 683700
rect 120040 683460 120130 683700
rect 120370 683460 120460 683700
rect 120700 683460 120790 683700
rect 121030 683460 121120 683700
rect 121360 683460 121450 683700
rect 121690 683460 122270 683700
rect 122510 683460 122600 683700
rect 122840 683460 122930 683700
rect 123170 683460 123260 683700
rect 123500 683460 123590 683700
rect 123830 683460 123920 683700
rect 124160 683460 124250 683700
rect 124490 683460 124580 683700
rect 124820 683460 124910 683700
rect 125150 683460 125240 683700
rect 125480 683460 125570 683700
rect 125810 683460 125900 683700
rect 126140 683460 126230 683700
rect 126470 683460 126560 683700
rect 126800 683460 126890 683700
rect 127130 683460 127220 683700
rect 127460 683460 127550 683700
rect 127790 683460 127880 683700
rect 128120 683460 128210 683700
rect 128450 683460 128540 683700
rect 128780 683460 128870 683700
rect 129110 683460 129200 683700
rect 129440 683460 129530 683700
rect 129770 683460 129860 683700
rect 130100 683460 130190 683700
rect 130430 683460 130520 683700
rect 130760 683460 130850 683700
rect 131090 683460 131180 683700
rect 131420 683460 131510 683700
rect 131750 683460 131840 683700
rect 132080 683460 132170 683700
rect 132410 683460 132500 683700
rect 132740 683460 132830 683700
rect 133070 683460 133650 683700
rect 133890 683460 133980 683700
rect 134220 683460 134310 683700
rect 134550 683460 134640 683700
rect 134880 683460 134970 683700
rect 135210 683460 135300 683700
rect 135540 683460 135630 683700
rect 135870 683460 135960 683700
rect 136200 683460 136290 683700
rect 136530 683460 136620 683700
rect 136860 683460 136950 683700
rect 137190 683460 137280 683700
rect 137520 683460 137610 683700
rect 137850 683460 137940 683700
rect 138180 683460 138270 683700
rect 138510 683460 138600 683700
rect 138840 683460 138930 683700
rect 139170 683460 139260 683700
rect 139500 683460 139590 683700
rect 139830 683460 139920 683700
rect 140160 683460 140250 683700
rect 140490 683460 140580 683700
rect 140820 683460 140910 683700
rect 141150 683460 141240 683700
rect 141480 683460 141570 683700
rect 141810 683460 141900 683700
rect 142140 683460 142230 683700
rect 142470 683460 142560 683700
rect 142800 683460 142890 683700
rect 143130 683460 143220 683700
rect 143460 683460 143550 683700
rect 143790 683460 143880 683700
rect 144120 683460 144210 683700
rect 144450 683460 145030 683700
rect 145270 683460 145360 683700
rect 145600 683460 145690 683700
rect 145930 683460 146020 683700
rect 146260 683460 146350 683700
rect 146590 683460 146680 683700
rect 146920 683460 147010 683700
rect 147250 683460 147340 683700
rect 147580 683460 147670 683700
rect 147910 683460 148000 683700
rect 148240 683460 148330 683700
rect 148570 683460 148660 683700
rect 148900 683460 148990 683700
rect 149230 683460 149320 683700
rect 149560 683460 149650 683700
rect 149890 683460 149980 683700
rect 150220 683460 150310 683700
rect 150550 683460 150640 683700
rect 150880 683460 150970 683700
rect 151210 683460 151300 683700
rect 151540 683460 151630 683700
rect 151870 683460 151960 683700
rect 152200 683460 152290 683700
rect 152530 683460 152620 683700
rect 152860 683460 152950 683700
rect 153190 683460 153280 683700
rect 153520 683460 153610 683700
rect 153850 683460 153940 683700
rect 154180 683460 154270 683700
rect 154510 683460 154600 683700
rect 154840 683460 154930 683700
rect 155170 683460 155260 683700
rect 155500 683460 155590 683700
rect 155830 683460 155960 683700
rect 110760 660760 155960 683460
rect 582300 679930 584800 682984
rect 582300 679860 582950 679930
rect 583020 679860 583050 679930
rect 583120 679860 583150 679930
rect 583220 679860 584800 679930
rect 582300 679830 584800 679860
rect 582300 679760 582950 679830
rect 583020 679760 583050 679830
rect 583120 679760 583150 679830
rect 583220 679760 584800 679830
rect 582300 679730 584800 679760
rect 582300 679660 582950 679730
rect 583020 679660 583050 679730
rect 583120 679660 583150 679730
rect 583220 679660 584800 679730
rect 582300 677984 584800 679660
rect 110760 660520 110890 660760
rect 111130 660520 111220 660760
rect 111460 660520 111550 660760
rect 111790 660520 111880 660760
rect 112120 660520 112210 660760
rect 112450 660520 112540 660760
rect 112780 660520 112870 660760
rect 113110 660520 113200 660760
rect 113440 660520 113530 660760
rect 113770 660520 113860 660760
rect 114100 660520 114190 660760
rect 114430 660520 114520 660760
rect 114760 660520 114850 660760
rect 115090 660520 115180 660760
rect 115420 660520 115510 660760
rect 115750 660520 115840 660760
rect 116080 660520 116170 660760
rect 116410 660520 116500 660760
rect 116740 660520 116830 660760
rect 117070 660520 117160 660760
rect 117400 660520 117490 660760
rect 117730 660520 117820 660760
rect 118060 660520 118150 660760
rect 118390 660520 118480 660760
rect 118720 660520 118810 660760
rect 119050 660520 119140 660760
rect 119380 660520 119470 660760
rect 119710 660520 119800 660760
rect 120040 660520 120130 660760
rect 120370 660520 120460 660760
rect 120700 660520 120790 660760
rect 121030 660520 121120 660760
rect 121360 660520 121450 660760
rect 121690 660520 122270 660760
rect 122510 660520 122600 660760
rect 122840 660520 122930 660760
rect 123170 660520 123260 660760
rect 123500 660520 123590 660760
rect 123830 660520 123920 660760
rect 124160 660520 124250 660760
rect 124490 660520 124580 660760
rect 124820 660520 124910 660760
rect 125150 660520 125240 660760
rect 125480 660520 125570 660760
rect 125810 660520 125900 660760
rect 126140 660520 126230 660760
rect 126470 660520 126560 660760
rect 126800 660520 126890 660760
rect 127130 660520 127220 660760
rect 127460 660520 127550 660760
rect 127790 660520 127880 660760
rect 128120 660520 128210 660760
rect 128450 660520 128540 660760
rect 128780 660520 128870 660760
rect 129110 660520 129200 660760
rect 129440 660520 129530 660760
rect 129770 660520 129860 660760
rect 130100 660520 130190 660760
rect 130430 660520 130520 660760
rect 130760 660520 130850 660760
rect 131090 660520 131180 660760
rect 131420 660520 131510 660760
rect 131750 660520 131840 660760
rect 132080 660520 132170 660760
rect 132410 660520 132500 660760
rect 132740 660520 132830 660760
rect 133070 660520 133650 660760
rect 133890 660520 133980 660760
rect 134220 660520 134310 660760
rect 134550 660520 134640 660760
rect 134880 660520 134970 660760
rect 135210 660520 135300 660760
rect 135540 660520 135630 660760
rect 135870 660520 135960 660760
rect 136200 660520 136290 660760
rect 136530 660520 136620 660760
rect 136860 660520 136950 660760
rect 137190 660520 137280 660760
rect 137520 660520 137610 660760
rect 137850 660520 137940 660760
rect 138180 660520 138270 660760
rect 138510 660520 138600 660760
rect 138840 660520 138930 660760
rect 139170 660520 139260 660760
rect 139500 660520 139590 660760
rect 139830 660520 139920 660760
rect 140160 660520 140250 660760
rect 140490 660520 140580 660760
rect 140820 660520 140910 660760
rect 141150 660520 141240 660760
rect 141480 660520 141570 660760
rect 141810 660520 141900 660760
rect 142140 660520 142230 660760
rect 142470 660520 142560 660760
rect 142800 660520 142890 660760
rect 143130 660520 143220 660760
rect 143460 660520 143550 660760
rect 143790 660520 143880 660760
rect 144120 660520 144210 660760
rect 144450 660520 145030 660760
rect 145270 660520 145360 660760
rect 145600 660520 145690 660760
rect 145930 660520 146020 660760
rect 146260 660520 146350 660760
rect 146590 660520 146680 660760
rect 146920 660520 147010 660760
rect 147250 660520 147340 660760
rect 147580 660520 147670 660760
rect 147910 660520 148000 660760
rect 148240 660520 148330 660760
rect 148570 660520 148660 660760
rect 148900 660520 148990 660760
rect 149230 660520 149320 660760
rect 149560 660520 149650 660760
rect 149890 660520 149980 660760
rect 150220 660520 150310 660760
rect 150550 660520 150640 660760
rect 150880 660520 150970 660760
rect 151210 660520 151300 660760
rect 151540 660520 151630 660760
rect 151870 660520 151960 660760
rect 152200 660520 152290 660760
rect 152530 660520 152620 660760
rect 152860 660520 152950 660760
rect 153190 660520 153280 660760
rect 153520 660520 153610 660760
rect 153850 660520 153940 660760
rect 154180 660520 154270 660760
rect 154510 660520 154600 660760
rect 154840 660520 154930 660760
rect 155170 660520 155260 660760
rect 155500 660520 155590 660760
rect 155830 660520 155960 660760
rect 110760 649330 155960 660520
rect -800 643842 1660 648642
rect 196654 647380 196974 647600
rect 196654 647310 196680 647380
rect 196750 647310 196780 647380
rect 196850 647310 196880 647380
rect 196950 647310 196974 647380
rect 196654 647290 196974 647310
rect 196654 647220 196680 647290
rect 196750 647220 196780 647290
rect 196850 647220 196880 647290
rect 196950 647220 196974 647290
rect 196654 647190 196974 647220
rect 201214 647380 201534 647600
rect 201214 647310 201238 647380
rect 201308 647310 201338 647380
rect 201408 647310 201438 647380
rect 201508 647310 201534 647380
rect 201214 647290 201534 647310
rect 201214 647220 201238 647290
rect 201308 647220 201338 647290
rect 201408 647220 201438 647290
rect 201508 647220 201534 647290
rect 201214 647190 201534 647220
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 16352 703500 16652 703800
rect 16852 703500 17152 703800
rect 17352 703500 17652 703800
rect 17852 703500 18152 703800
rect 18352 703500 18652 703800
rect 18852 703500 19152 703800
rect 19352 703500 19652 703800
rect 19852 703500 20152 703800
rect 20352 703500 20652 703800
rect 20852 703500 21152 703800
rect 16352 703000 16652 703300
rect 16852 703000 17152 703300
rect 17352 703000 17652 703300
rect 17852 703000 18152 703300
rect 18352 703000 18652 703300
rect 18852 703000 19152 703300
rect 19352 703000 19652 703300
rect 19852 703000 20152 703300
rect 20352 703000 20652 703300
rect 20852 703000 21152 703300
rect 16352 702500 16652 702800
rect 16852 702500 17152 702800
rect 17352 702500 17652 702800
rect 17852 702500 18152 702800
rect 18352 702500 18652 702800
rect 18852 702500 19152 702800
rect 19352 702500 19652 702800
rect 19852 702500 20152 702800
rect 20352 702500 20652 702800
rect 20852 702500 21152 702800
rect 70300 703000 70500 703200
rect 70600 703000 70800 703200
rect 70900 703000 71100 703200
rect 70300 702700 70500 702900
rect 70600 702700 70800 702900
rect 70900 702700 71100 702900
rect 70300 702400 70500 702600
rect 70600 702400 70800 702600
rect 70900 702400 71100 702600
rect 122179 702994 122379 703194
rect 122479 702994 122679 703194
rect 122779 702994 122979 703194
rect 122179 702694 122379 702894
rect 122479 702694 122679 702894
rect 122779 702694 122979 702894
rect 122179 702394 122379 702594
rect 122479 702394 122679 702594
rect 122779 702394 122979 702594
rect 415760 703040 415830 703110
rect 415850 703040 415920 703110
rect 415940 703040 416010 703110
rect 416030 703040 416100 703110
rect 416120 703040 416190 703110
rect 415760 702950 415830 703020
rect 415850 702950 415920 703020
rect 415940 702950 416010 703020
rect 416030 702950 416100 703020
rect 416120 702950 416190 703020
rect 415760 702860 415830 702930
rect 415850 702860 415920 702930
rect 415940 702860 416010 702930
rect 416030 702860 416100 702930
rect 416120 702860 416190 702930
rect 415760 702770 415830 702840
rect 415850 702770 415920 702840
rect 415940 702770 416010 702840
rect 416030 702770 416100 702840
rect 416120 702770 416190 702840
rect 415760 702680 415830 702750
rect 415850 702680 415920 702750
rect 415940 702680 416010 702750
rect 416030 702680 416100 702750
rect 416120 702680 416190 702750
rect 467220 703240 467290 703310
rect 467320 703240 467390 703310
rect 467420 703240 467490 703310
rect 467220 703150 467290 703220
rect 467320 703150 467390 703220
rect 467420 703150 467490 703220
rect 467220 703060 467290 703130
rect 467320 703060 467390 703130
rect 467420 703060 467490 703130
rect 569600 702800 569670 702870
rect 569700 702800 569770 702870
rect 569800 702800 569870 702870
rect 569600 702700 569670 702770
rect 569700 702700 569770 702770
rect 569800 702700 569870 702770
rect 569600 702600 569670 702670
rect 569700 702600 569770 702670
rect 569800 702600 569870 702670
rect 200 684900 500 685200
rect 700 684900 1000 685200
rect 1200 684900 1500 685200
rect 200 684400 500 684700
rect 700 684400 1000 684700
rect 1200 684400 1500 684700
rect 200 683900 500 684200
rect 700 683900 1000 684200
rect 1200 683900 1500 684200
rect 200 683400 500 683700
rect 700 683400 1000 683700
rect 1200 683400 1500 683700
rect 200 682900 500 683200
rect 700 682900 1000 683200
rect 1200 682900 1500 683200
rect 200 682400 500 682700
rect 700 682400 1000 682700
rect 1200 682400 1500 682700
rect 200 681900 500 682200
rect 700 681900 1000 682200
rect 1200 681900 1500 682200
rect 200 681400 500 681700
rect 700 681400 1000 681700
rect 1200 681400 1500 681700
rect 200 680900 500 681200
rect 700 680900 1000 681200
rect 1200 680900 1500 681200
rect 200 680400 500 680700
rect 700 680400 1000 680700
rect 1200 680400 1500 680700
rect 110890 683460 111130 683700
rect 111220 683460 111460 683700
rect 111550 683460 111790 683700
rect 111880 683460 112120 683700
rect 112210 683460 112450 683700
rect 112540 683460 112780 683700
rect 112870 683460 113110 683700
rect 113200 683460 113440 683700
rect 113530 683460 113770 683700
rect 113860 683460 114100 683700
rect 114190 683460 114430 683700
rect 114520 683460 114760 683700
rect 114850 683460 115090 683700
rect 115180 683460 115420 683700
rect 115510 683460 115750 683700
rect 115840 683460 116080 683700
rect 116170 683460 116410 683700
rect 116500 683460 116740 683700
rect 116830 683460 117070 683700
rect 117160 683460 117400 683700
rect 117490 683460 117730 683700
rect 117820 683460 118060 683700
rect 118150 683460 118390 683700
rect 118480 683460 118720 683700
rect 118810 683460 119050 683700
rect 119140 683460 119380 683700
rect 119470 683460 119710 683700
rect 119800 683460 120040 683700
rect 120130 683460 120370 683700
rect 120460 683460 120700 683700
rect 120790 683460 121030 683700
rect 121120 683460 121360 683700
rect 121450 683460 121690 683700
rect 122270 683460 122510 683700
rect 122600 683460 122840 683700
rect 122930 683460 123170 683700
rect 123260 683460 123500 683700
rect 123590 683460 123830 683700
rect 123920 683460 124160 683700
rect 124250 683460 124490 683700
rect 124580 683460 124820 683700
rect 124910 683460 125150 683700
rect 125240 683460 125480 683700
rect 125570 683460 125810 683700
rect 125900 683460 126140 683700
rect 126230 683460 126470 683700
rect 126560 683460 126800 683700
rect 126890 683460 127130 683700
rect 127220 683460 127460 683700
rect 127550 683460 127790 683700
rect 127880 683460 128120 683700
rect 128210 683460 128450 683700
rect 128540 683460 128780 683700
rect 128870 683460 129110 683700
rect 129200 683460 129440 683700
rect 129530 683460 129770 683700
rect 129860 683460 130100 683700
rect 130190 683460 130430 683700
rect 130520 683460 130760 683700
rect 130850 683460 131090 683700
rect 131180 683460 131420 683700
rect 131510 683460 131750 683700
rect 131840 683460 132080 683700
rect 132170 683460 132410 683700
rect 132500 683460 132740 683700
rect 132830 683460 133070 683700
rect 133650 683460 133890 683700
rect 133980 683460 134220 683700
rect 134310 683460 134550 683700
rect 134640 683460 134880 683700
rect 134970 683460 135210 683700
rect 135300 683460 135540 683700
rect 135630 683460 135870 683700
rect 135960 683460 136200 683700
rect 136290 683460 136530 683700
rect 136620 683460 136860 683700
rect 136950 683460 137190 683700
rect 137280 683460 137520 683700
rect 137610 683460 137850 683700
rect 137940 683460 138180 683700
rect 138270 683460 138510 683700
rect 138600 683460 138840 683700
rect 138930 683460 139170 683700
rect 139260 683460 139500 683700
rect 139590 683460 139830 683700
rect 139920 683460 140160 683700
rect 140250 683460 140490 683700
rect 140580 683460 140820 683700
rect 140910 683460 141150 683700
rect 141240 683460 141480 683700
rect 141570 683460 141810 683700
rect 141900 683460 142140 683700
rect 142230 683460 142470 683700
rect 142560 683460 142800 683700
rect 142890 683460 143130 683700
rect 143220 683460 143460 683700
rect 143550 683460 143790 683700
rect 143880 683460 144120 683700
rect 144210 683460 144450 683700
rect 145030 683460 145270 683700
rect 145360 683460 145600 683700
rect 145690 683460 145930 683700
rect 146020 683460 146260 683700
rect 146350 683460 146590 683700
rect 146680 683460 146920 683700
rect 147010 683460 147250 683700
rect 147340 683460 147580 683700
rect 147670 683460 147910 683700
rect 148000 683460 148240 683700
rect 148330 683460 148570 683700
rect 148660 683460 148900 683700
rect 148990 683460 149230 683700
rect 149320 683460 149560 683700
rect 149650 683460 149890 683700
rect 149980 683460 150220 683700
rect 150310 683460 150550 683700
rect 150640 683460 150880 683700
rect 150970 683460 151210 683700
rect 151300 683460 151540 683700
rect 151630 683460 151870 683700
rect 151960 683460 152200 683700
rect 152290 683460 152530 683700
rect 152620 683460 152860 683700
rect 152950 683460 153190 683700
rect 153280 683460 153520 683700
rect 153610 683460 153850 683700
rect 153940 683460 154180 683700
rect 154270 683460 154510 683700
rect 154600 683460 154840 683700
rect 154930 683460 155170 683700
rect 155260 683460 155500 683700
rect 155590 683460 155830 683700
rect 582950 679860 583020 679930
rect 583050 679860 583120 679930
rect 583150 679860 583220 679930
rect 582950 679760 583020 679830
rect 583050 679760 583120 679830
rect 583150 679760 583220 679830
rect 582950 679660 583020 679730
rect 583050 679660 583120 679730
rect 583150 679660 583220 679730
rect 110890 660520 111130 660760
rect 111220 660520 111460 660760
rect 111550 660520 111790 660760
rect 111880 660520 112120 660760
rect 112210 660520 112450 660760
rect 112540 660520 112780 660760
rect 112870 660520 113110 660760
rect 113200 660520 113440 660760
rect 113530 660520 113770 660760
rect 113860 660520 114100 660760
rect 114190 660520 114430 660760
rect 114520 660520 114760 660760
rect 114850 660520 115090 660760
rect 115180 660520 115420 660760
rect 115510 660520 115750 660760
rect 115840 660520 116080 660760
rect 116170 660520 116410 660760
rect 116500 660520 116740 660760
rect 116830 660520 117070 660760
rect 117160 660520 117400 660760
rect 117490 660520 117730 660760
rect 117820 660520 118060 660760
rect 118150 660520 118390 660760
rect 118480 660520 118720 660760
rect 118810 660520 119050 660760
rect 119140 660520 119380 660760
rect 119470 660520 119710 660760
rect 119800 660520 120040 660760
rect 120130 660520 120370 660760
rect 120460 660520 120700 660760
rect 120790 660520 121030 660760
rect 121120 660520 121360 660760
rect 121450 660520 121690 660760
rect 122270 660520 122510 660760
rect 122600 660520 122840 660760
rect 122930 660520 123170 660760
rect 123260 660520 123500 660760
rect 123590 660520 123830 660760
rect 123920 660520 124160 660760
rect 124250 660520 124490 660760
rect 124580 660520 124820 660760
rect 124910 660520 125150 660760
rect 125240 660520 125480 660760
rect 125570 660520 125810 660760
rect 125900 660520 126140 660760
rect 126230 660520 126470 660760
rect 126560 660520 126800 660760
rect 126890 660520 127130 660760
rect 127220 660520 127460 660760
rect 127550 660520 127790 660760
rect 127880 660520 128120 660760
rect 128210 660520 128450 660760
rect 128540 660520 128780 660760
rect 128870 660520 129110 660760
rect 129200 660520 129440 660760
rect 129530 660520 129770 660760
rect 129860 660520 130100 660760
rect 130190 660520 130430 660760
rect 130520 660520 130760 660760
rect 130850 660520 131090 660760
rect 131180 660520 131420 660760
rect 131510 660520 131750 660760
rect 131840 660520 132080 660760
rect 132170 660520 132410 660760
rect 132500 660520 132740 660760
rect 132830 660520 133070 660760
rect 133650 660520 133890 660760
rect 133980 660520 134220 660760
rect 134310 660520 134550 660760
rect 134640 660520 134880 660760
rect 134970 660520 135210 660760
rect 135300 660520 135540 660760
rect 135630 660520 135870 660760
rect 135960 660520 136200 660760
rect 136290 660520 136530 660760
rect 136620 660520 136860 660760
rect 136950 660520 137190 660760
rect 137280 660520 137520 660760
rect 137610 660520 137850 660760
rect 137940 660520 138180 660760
rect 138270 660520 138510 660760
rect 138600 660520 138840 660760
rect 138930 660520 139170 660760
rect 139260 660520 139500 660760
rect 139590 660520 139830 660760
rect 139920 660520 140160 660760
rect 140250 660520 140490 660760
rect 140580 660520 140820 660760
rect 140910 660520 141150 660760
rect 141240 660520 141480 660760
rect 141570 660520 141810 660760
rect 141900 660520 142140 660760
rect 142230 660520 142470 660760
rect 142560 660520 142800 660760
rect 142890 660520 143130 660760
rect 143220 660520 143460 660760
rect 143550 660520 143790 660760
rect 143880 660520 144120 660760
rect 144210 660520 144450 660760
rect 145030 660520 145270 660760
rect 145360 660520 145600 660760
rect 145690 660520 145930 660760
rect 146020 660520 146260 660760
rect 146350 660520 146590 660760
rect 146680 660520 146920 660760
rect 147010 660520 147250 660760
rect 147340 660520 147580 660760
rect 147670 660520 147910 660760
rect 148000 660520 148240 660760
rect 148330 660520 148570 660760
rect 148660 660520 148900 660760
rect 148990 660520 149230 660760
rect 149320 660520 149560 660760
rect 149650 660520 149890 660760
rect 149980 660520 150220 660760
rect 150310 660520 150550 660760
rect 150640 660520 150880 660760
rect 150970 660520 151210 660760
rect 151300 660520 151540 660760
rect 151630 660520 151870 660760
rect 151960 660520 152200 660760
rect 152290 660520 152530 660760
rect 152620 660520 152860 660760
rect 152950 660520 153190 660760
rect 153280 660520 153520 660760
rect 153610 660520 153850 660760
rect 153940 660520 154180 660760
rect 154270 660520 154510 660760
rect 154600 660520 154840 660760
rect 154930 660520 155170 660760
rect 155260 660520 155500 660760
rect 155590 660520 155830 660760
rect 196680 647310 196750 647380
rect 196780 647310 196850 647380
rect 196880 647310 196950 647380
rect 196680 647220 196750 647290
rect 196780 647220 196850 647290
rect 196880 647220 196950 647290
rect 201238 647310 201308 647380
rect 201338 647310 201408 647380
rect 201438 647310 201508 647380
rect 201238 647220 201308 647290
rect 201338 647220 201408 647290
rect 201438 647220 201508 647290
<< mimcap >>
rect 110790 694840 121790 694860
rect 110790 694600 110810 694840
rect 111050 694600 111140 694840
rect 111380 694600 111470 694840
rect 111710 694600 111800 694840
rect 112040 694600 112150 694840
rect 112390 694600 112480 694840
rect 112720 694600 112810 694840
rect 113050 694600 113140 694840
rect 113380 694600 113490 694840
rect 113730 694600 113820 694840
rect 114060 694600 114150 694840
rect 114390 694600 114480 694840
rect 114720 694600 114830 694840
rect 115070 694600 115160 694840
rect 115400 694600 115490 694840
rect 115730 694600 115820 694840
rect 116060 694600 116170 694840
rect 116410 694600 116500 694840
rect 116740 694600 116830 694840
rect 117070 694600 117160 694840
rect 117400 694600 117510 694840
rect 117750 694600 117840 694840
rect 118080 694600 118170 694840
rect 118410 694600 118500 694840
rect 118740 694600 118850 694840
rect 119090 694600 119180 694840
rect 119420 694600 119510 694840
rect 119750 694600 119840 694840
rect 120080 694600 120190 694840
rect 120430 694600 120520 694840
rect 120760 694600 120850 694840
rect 121090 694600 121180 694840
rect 121420 694600 121530 694840
rect 121770 694600 121790 694840
rect 110790 694490 121790 694600
rect 110790 694250 110810 694490
rect 111050 694250 111140 694490
rect 111380 694250 111470 694490
rect 111710 694250 111800 694490
rect 112040 694250 112150 694490
rect 112390 694250 112480 694490
rect 112720 694250 112810 694490
rect 113050 694250 113140 694490
rect 113380 694250 113490 694490
rect 113730 694250 113820 694490
rect 114060 694250 114150 694490
rect 114390 694250 114480 694490
rect 114720 694250 114830 694490
rect 115070 694250 115160 694490
rect 115400 694250 115490 694490
rect 115730 694250 115820 694490
rect 116060 694250 116170 694490
rect 116410 694250 116500 694490
rect 116740 694250 116830 694490
rect 117070 694250 117160 694490
rect 117400 694250 117510 694490
rect 117750 694250 117840 694490
rect 118080 694250 118170 694490
rect 118410 694250 118500 694490
rect 118740 694250 118850 694490
rect 119090 694250 119180 694490
rect 119420 694250 119510 694490
rect 119750 694250 119840 694490
rect 120080 694250 120190 694490
rect 120430 694250 120520 694490
rect 120760 694250 120850 694490
rect 121090 694250 121180 694490
rect 121420 694250 121530 694490
rect 121770 694250 121790 694490
rect 110790 694160 121790 694250
rect 110790 693920 110810 694160
rect 111050 693920 111140 694160
rect 111380 693920 111470 694160
rect 111710 693920 111800 694160
rect 112040 693920 112150 694160
rect 112390 693920 112480 694160
rect 112720 693920 112810 694160
rect 113050 693920 113140 694160
rect 113380 693920 113490 694160
rect 113730 693920 113820 694160
rect 114060 693920 114150 694160
rect 114390 693920 114480 694160
rect 114720 693920 114830 694160
rect 115070 693920 115160 694160
rect 115400 693920 115490 694160
rect 115730 693920 115820 694160
rect 116060 693920 116170 694160
rect 116410 693920 116500 694160
rect 116740 693920 116830 694160
rect 117070 693920 117160 694160
rect 117400 693920 117510 694160
rect 117750 693920 117840 694160
rect 118080 693920 118170 694160
rect 118410 693920 118500 694160
rect 118740 693920 118850 694160
rect 119090 693920 119180 694160
rect 119420 693920 119510 694160
rect 119750 693920 119840 694160
rect 120080 693920 120190 694160
rect 120430 693920 120520 694160
rect 120760 693920 120850 694160
rect 121090 693920 121180 694160
rect 121420 693920 121530 694160
rect 121770 693920 121790 694160
rect 110790 693830 121790 693920
rect 110790 693590 110810 693830
rect 111050 693590 111140 693830
rect 111380 693590 111470 693830
rect 111710 693590 111800 693830
rect 112040 693590 112150 693830
rect 112390 693590 112480 693830
rect 112720 693590 112810 693830
rect 113050 693590 113140 693830
rect 113380 693590 113490 693830
rect 113730 693590 113820 693830
rect 114060 693590 114150 693830
rect 114390 693590 114480 693830
rect 114720 693590 114830 693830
rect 115070 693590 115160 693830
rect 115400 693590 115490 693830
rect 115730 693590 115820 693830
rect 116060 693590 116170 693830
rect 116410 693590 116500 693830
rect 116740 693590 116830 693830
rect 117070 693590 117160 693830
rect 117400 693590 117510 693830
rect 117750 693590 117840 693830
rect 118080 693590 118170 693830
rect 118410 693590 118500 693830
rect 118740 693590 118850 693830
rect 119090 693590 119180 693830
rect 119420 693590 119510 693830
rect 119750 693590 119840 693830
rect 120080 693590 120190 693830
rect 120430 693590 120520 693830
rect 120760 693590 120850 693830
rect 121090 693590 121180 693830
rect 121420 693590 121530 693830
rect 121770 693590 121790 693830
rect 110790 693500 121790 693590
rect 110790 693260 110810 693500
rect 111050 693260 111140 693500
rect 111380 693260 111470 693500
rect 111710 693260 111800 693500
rect 112040 693260 112150 693500
rect 112390 693260 112480 693500
rect 112720 693260 112810 693500
rect 113050 693260 113140 693500
rect 113380 693260 113490 693500
rect 113730 693260 113820 693500
rect 114060 693260 114150 693500
rect 114390 693260 114480 693500
rect 114720 693260 114830 693500
rect 115070 693260 115160 693500
rect 115400 693260 115490 693500
rect 115730 693260 115820 693500
rect 116060 693260 116170 693500
rect 116410 693260 116500 693500
rect 116740 693260 116830 693500
rect 117070 693260 117160 693500
rect 117400 693260 117510 693500
rect 117750 693260 117840 693500
rect 118080 693260 118170 693500
rect 118410 693260 118500 693500
rect 118740 693260 118850 693500
rect 119090 693260 119180 693500
rect 119420 693260 119510 693500
rect 119750 693260 119840 693500
rect 120080 693260 120190 693500
rect 120430 693260 120520 693500
rect 120760 693260 120850 693500
rect 121090 693260 121180 693500
rect 121420 693260 121530 693500
rect 121770 693260 121790 693500
rect 110790 693150 121790 693260
rect 110790 692910 110810 693150
rect 111050 692910 111140 693150
rect 111380 692910 111470 693150
rect 111710 692910 111800 693150
rect 112040 692910 112150 693150
rect 112390 692910 112480 693150
rect 112720 692910 112810 693150
rect 113050 692910 113140 693150
rect 113380 692910 113490 693150
rect 113730 692910 113820 693150
rect 114060 692910 114150 693150
rect 114390 692910 114480 693150
rect 114720 692910 114830 693150
rect 115070 692910 115160 693150
rect 115400 692910 115490 693150
rect 115730 692910 115820 693150
rect 116060 692910 116170 693150
rect 116410 692910 116500 693150
rect 116740 692910 116830 693150
rect 117070 692910 117160 693150
rect 117400 692910 117510 693150
rect 117750 692910 117840 693150
rect 118080 692910 118170 693150
rect 118410 692910 118500 693150
rect 118740 692910 118850 693150
rect 119090 692910 119180 693150
rect 119420 692910 119510 693150
rect 119750 692910 119840 693150
rect 120080 692910 120190 693150
rect 120430 692910 120520 693150
rect 120760 692910 120850 693150
rect 121090 692910 121180 693150
rect 121420 692910 121530 693150
rect 121770 692910 121790 693150
rect 110790 692820 121790 692910
rect 110790 692580 110810 692820
rect 111050 692580 111140 692820
rect 111380 692580 111470 692820
rect 111710 692580 111800 692820
rect 112040 692580 112150 692820
rect 112390 692580 112480 692820
rect 112720 692580 112810 692820
rect 113050 692580 113140 692820
rect 113380 692580 113490 692820
rect 113730 692580 113820 692820
rect 114060 692580 114150 692820
rect 114390 692580 114480 692820
rect 114720 692580 114830 692820
rect 115070 692580 115160 692820
rect 115400 692580 115490 692820
rect 115730 692580 115820 692820
rect 116060 692580 116170 692820
rect 116410 692580 116500 692820
rect 116740 692580 116830 692820
rect 117070 692580 117160 692820
rect 117400 692580 117510 692820
rect 117750 692580 117840 692820
rect 118080 692580 118170 692820
rect 118410 692580 118500 692820
rect 118740 692580 118850 692820
rect 119090 692580 119180 692820
rect 119420 692580 119510 692820
rect 119750 692580 119840 692820
rect 120080 692580 120190 692820
rect 120430 692580 120520 692820
rect 120760 692580 120850 692820
rect 121090 692580 121180 692820
rect 121420 692580 121530 692820
rect 121770 692580 121790 692820
rect 110790 692490 121790 692580
rect 110790 692250 110810 692490
rect 111050 692250 111140 692490
rect 111380 692250 111470 692490
rect 111710 692250 111800 692490
rect 112040 692250 112150 692490
rect 112390 692250 112480 692490
rect 112720 692250 112810 692490
rect 113050 692250 113140 692490
rect 113380 692250 113490 692490
rect 113730 692250 113820 692490
rect 114060 692250 114150 692490
rect 114390 692250 114480 692490
rect 114720 692250 114830 692490
rect 115070 692250 115160 692490
rect 115400 692250 115490 692490
rect 115730 692250 115820 692490
rect 116060 692250 116170 692490
rect 116410 692250 116500 692490
rect 116740 692250 116830 692490
rect 117070 692250 117160 692490
rect 117400 692250 117510 692490
rect 117750 692250 117840 692490
rect 118080 692250 118170 692490
rect 118410 692250 118500 692490
rect 118740 692250 118850 692490
rect 119090 692250 119180 692490
rect 119420 692250 119510 692490
rect 119750 692250 119840 692490
rect 120080 692250 120190 692490
rect 120430 692250 120520 692490
rect 120760 692250 120850 692490
rect 121090 692250 121180 692490
rect 121420 692250 121530 692490
rect 121770 692250 121790 692490
rect 110790 692160 121790 692250
rect 110790 691920 110810 692160
rect 111050 691920 111140 692160
rect 111380 691920 111470 692160
rect 111710 691920 111800 692160
rect 112040 691920 112150 692160
rect 112390 691920 112480 692160
rect 112720 691920 112810 692160
rect 113050 691920 113140 692160
rect 113380 691920 113490 692160
rect 113730 691920 113820 692160
rect 114060 691920 114150 692160
rect 114390 691920 114480 692160
rect 114720 691920 114830 692160
rect 115070 691920 115160 692160
rect 115400 691920 115490 692160
rect 115730 691920 115820 692160
rect 116060 691920 116170 692160
rect 116410 691920 116500 692160
rect 116740 691920 116830 692160
rect 117070 691920 117160 692160
rect 117400 691920 117510 692160
rect 117750 691920 117840 692160
rect 118080 691920 118170 692160
rect 118410 691920 118500 692160
rect 118740 691920 118850 692160
rect 119090 691920 119180 692160
rect 119420 691920 119510 692160
rect 119750 691920 119840 692160
rect 120080 691920 120190 692160
rect 120430 691920 120520 692160
rect 120760 691920 120850 692160
rect 121090 691920 121180 692160
rect 121420 691920 121530 692160
rect 121770 691920 121790 692160
rect 110790 691810 121790 691920
rect 110790 691570 110810 691810
rect 111050 691570 111140 691810
rect 111380 691570 111470 691810
rect 111710 691570 111800 691810
rect 112040 691570 112150 691810
rect 112390 691570 112480 691810
rect 112720 691570 112810 691810
rect 113050 691570 113140 691810
rect 113380 691570 113490 691810
rect 113730 691570 113820 691810
rect 114060 691570 114150 691810
rect 114390 691570 114480 691810
rect 114720 691570 114830 691810
rect 115070 691570 115160 691810
rect 115400 691570 115490 691810
rect 115730 691570 115820 691810
rect 116060 691570 116170 691810
rect 116410 691570 116500 691810
rect 116740 691570 116830 691810
rect 117070 691570 117160 691810
rect 117400 691570 117510 691810
rect 117750 691570 117840 691810
rect 118080 691570 118170 691810
rect 118410 691570 118500 691810
rect 118740 691570 118850 691810
rect 119090 691570 119180 691810
rect 119420 691570 119510 691810
rect 119750 691570 119840 691810
rect 120080 691570 120190 691810
rect 120430 691570 120520 691810
rect 120760 691570 120850 691810
rect 121090 691570 121180 691810
rect 121420 691570 121530 691810
rect 121770 691570 121790 691810
rect 110790 691480 121790 691570
rect 110790 691240 110810 691480
rect 111050 691240 111140 691480
rect 111380 691240 111470 691480
rect 111710 691240 111800 691480
rect 112040 691240 112150 691480
rect 112390 691240 112480 691480
rect 112720 691240 112810 691480
rect 113050 691240 113140 691480
rect 113380 691240 113490 691480
rect 113730 691240 113820 691480
rect 114060 691240 114150 691480
rect 114390 691240 114480 691480
rect 114720 691240 114830 691480
rect 115070 691240 115160 691480
rect 115400 691240 115490 691480
rect 115730 691240 115820 691480
rect 116060 691240 116170 691480
rect 116410 691240 116500 691480
rect 116740 691240 116830 691480
rect 117070 691240 117160 691480
rect 117400 691240 117510 691480
rect 117750 691240 117840 691480
rect 118080 691240 118170 691480
rect 118410 691240 118500 691480
rect 118740 691240 118850 691480
rect 119090 691240 119180 691480
rect 119420 691240 119510 691480
rect 119750 691240 119840 691480
rect 120080 691240 120190 691480
rect 120430 691240 120520 691480
rect 120760 691240 120850 691480
rect 121090 691240 121180 691480
rect 121420 691240 121530 691480
rect 121770 691240 121790 691480
rect 110790 691150 121790 691240
rect 110790 690910 110810 691150
rect 111050 690910 111140 691150
rect 111380 690910 111470 691150
rect 111710 690910 111800 691150
rect 112040 690910 112150 691150
rect 112390 690910 112480 691150
rect 112720 690910 112810 691150
rect 113050 690910 113140 691150
rect 113380 690910 113490 691150
rect 113730 690910 113820 691150
rect 114060 690910 114150 691150
rect 114390 690910 114480 691150
rect 114720 690910 114830 691150
rect 115070 690910 115160 691150
rect 115400 690910 115490 691150
rect 115730 690910 115820 691150
rect 116060 690910 116170 691150
rect 116410 690910 116500 691150
rect 116740 690910 116830 691150
rect 117070 690910 117160 691150
rect 117400 690910 117510 691150
rect 117750 690910 117840 691150
rect 118080 690910 118170 691150
rect 118410 690910 118500 691150
rect 118740 690910 118850 691150
rect 119090 690910 119180 691150
rect 119420 690910 119510 691150
rect 119750 690910 119840 691150
rect 120080 690910 120190 691150
rect 120430 690910 120520 691150
rect 120760 690910 120850 691150
rect 121090 690910 121180 691150
rect 121420 690910 121530 691150
rect 121770 690910 121790 691150
rect 110790 690820 121790 690910
rect 110790 690580 110810 690820
rect 111050 690580 111140 690820
rect 111380 690580 111470 690820
rect 111710 690580 111800 690820
rect 112040 690580 112150 690820
rect 112390 690580 112480 690820
rect 112720 690580 112810 690820
rect 113050 690580 113140 690820
rect 113380 690580 113490 690820
rect 113730 690580 113820 690820
rect 114060 690580 114150 690820
rect 114390 690580 114480 690820
rect 114720 690580 114830 690820
rect 115070 690580 115160 690820
rect 115400 690580 115490 690820
rect 115730 690580 115820 690820
rect 116060 690580 116170 690820
rect 116410 690580 116500 690820
rect 116740 690580 116830 690820
rect 117070 690580 117160 690820
rect 117400 690580 117510 690820
rect 117750 690580 117840 690820
rect 118080 690580 118170 690820
rect 118410 690580 118500 690820
rect 118740 690580 118850 690820
rect 119090 690580 119180 690820
rect 119420 690580 119510 690820
rect 119750 690580 119840 690820
rect 120080 690580 120190 690820
rect 120430 690580 120520 690820
rect 120760 690580 120850 690820
rect 121090 690580 121180 690820
rect 121420 690580 121530 690820
rect 121770 690580 121790 690820
rect 110790 690470 121790 690580
rect 110790 690230 110810 690470
rect 111050 690230 111140 690470
rect 111380 690230 111470 690470
rect 111710 690230 111800 690470
rect 112040 690230 112150 690470
rect 112390 690230 112480 690470
rect 112720 690230 112810 690470
rect 113050 690230 113140 690470
rect 113380 690230 113490 690470
rect 113730 690230 113820 690470
rect 114060 690230 114150 690470
rect 114390 690230 114480 690470
rect 114720 690230 114830 690470
rect 115070 690230 115160 690470
rect 115400 690230 115490 690470
rect 115730 690230 115820 690470
rect 116060 690230 116170 690470
rect 116410 690230 116500 690470
rect 116740 690230 116830 690470
rect 117070 690230 117160 690470
rect 117400 690230 117510 690470
rect 117750 690230 117840 690470
rect 118080 690230 118170 690470
rect 118410 690230 118500 690470
rect 118740 690230 118850 690470
rect 119090 690230 119180 690470
rect 119420 690230 119510 690470
rect 119750 690230 119840 690470
rect 120080 690230 120190 690470
rect 120430 690230 120520 690470
rect 120760 690230 120850 690470
rect 121090 690230 121180 690470
rect 121420 690230 121530 690470
rect 121770 690230 121790 690470
rect 110790 690140 121790 690230
rect 110790 689900 110810 690140
rect 111050 689900 111140 690140
rect 111380 689900 111470 690140
rect 111710 689900 111800 690140
rect 112040 689900 112150 690140
rect 112390 689900 112480 690140
rect 112720 689900 112810 690140
rect 113050 689900 113140 690140
rect 113380 689900 113490 690140
rect 113730 689900 113820 690140
rect 114060 689900 114150 690140
rect 114390 689900 114480 690140
rect 114720 689900 114830 690140
rect 115070 689900 115160 690140
rect 115400 689900 115490 690140
rect 115730 689900 115820 690140
rect 116060 689900 116170 690140
rect 116410 689900 116500 690140
rect 116740 689900 116830 690140
rect 117070 689900 117160 690140
rect 117400 689900 117510 690140
rect 117750 689900 117840 690140
rect 118080 689900 118170 690140
rect 118410 689900 118500 690140
rect 118740 689900 118850 690140
rect 119090 689900 119180 690140
rect 119420 689900 119510 690140
rect 119750 689900 119840 690140
rect 120080 689900 120190 690140
rect 120430 689900 120520 690140
rect 120760 689900 120850 690140
rect 121090 689900 121180 690140
rect 121420 689900 121530 690140
rect 121770 689900 121790 690140
rect 110790 689810 121790 689900
rect 110790 689570 110810 689810
rect 111050 689570 111140 689810
rect 111380 689570 111470 689810
rect 111710 689570 111800 689810
rect 112040 689570 112150 689810
rect 112390 689570 112480 689810
rect 112720 689570 112810 689810
rect 113050 689570 113140 689810
rect 113380 689570 113490 689810
rect 113730 689570 113820 689810
rect 114060 689570 114150 689810
rect 114390 689570 114480 689810
rect 114720 689570 114830 689810
rect 115070 689570 115160 689810
rect 115400 689570 115490 689810
rect 115730 689570 115820 689810
rect 116060 689570 116170 689810
rect 116410 689570 116500 689810
rect 116740 689570 116830 689810
rect 117070 689570 117160 689810
rect 117400 689570 117510 689810
rect 117750 689570 117840 689810
rect 118080 689570 118170 689810
rect 118410 689570 118500 689810
rect 118740 689570 118850 689810
rect 119090 689570 119180 689810
rect 119420 689570 119510 689810
rect 119750 689570 119840 689810
rect 120080 689570 120190 689810
rect 120430 689570 120520 689810
rect 120760 689570 120850 689810
rect 121090 689570 121180 689810
rect 121420 689570 121530 689810
rect 121770 689570 121790 689810
rect 110790 689480 121790 689570
rect 110790 689240 110810 689480
rect 111050 689240 111140 689480
rect 111380 689240 111470 689480
rect 111710 689240 111800 689480
rect 112040 689240 112150 689480
rect 112390 689240 112480 689480
rect 112720 689240 112810 689480
rect 113050 689240 113140 689480
rect 113380 689240 113490 689480
rect 113730 689240 113820 689480
rect 114060 689240 114150 689480
rect 114390 689240 114480 689480
rect 114720 689240 114830 689480
rect 115070 689240 115160 689480
rect 115400 689240 115490 689480
rect 115730 689240 115820 689480
rect 116060 689240 116170 689480
rect 116410 689240 116500 689480
rect 116740 689240 116830 689480
rect 117070 689240 117160 689480
rect 117400 689240 117510 689480
rect 117750 689240 117840 689480
rect 118080 689240 118170 689480
rect 118410 689240 118500 689480
rect 118740 689240 118850 689480
rect 119090 689240 119180 689480
rect 119420 689240 119510 689480
rect 119750 689240 119840 689480
rect 120080 689240 120190 689480
rect 120430 689240 120520 689480
rect 120760 689240 120850 689480
rect 121090 689240 121180 689480
rect 121420 689240 121530 689480
rect 121770 689240 121790 689480
rect 110790 689130 121790 689240
rect 110790 688890 110810 689130
rect 111050 688890 111140 689130
rect 111380 688890 111470 689130
rect 111710 688890 111800 689130
rect 112040 688890 112150 689130
rect 112390 688890 112480 689130
rect 112720 688890 112810 689130
rect 113050 688890 113140 689130
rect 113380 688890 113490 689130
rect 113730 688890 113820 689130
rect 114060 688890 114150 689130
rect 114390 688890 114480 689130
rect 114720 688890 114830 689130
rect 115070 688890 115160 689130
rect 115400 688890 115490 689130
rect 115730 688890 115820 689130
rect 116060 688890 116170 689130
rect 116410 688890 116500 689130
rect 116740 688890 116830 689130
rect 117070 688890 117160 689130
rect 117400 688890 117510 689130
rect 117750 688890 117840 689130
rect 118080 688890 118170 689130
rect 118410 688890 118500 689130
rect 118740 688890 118850 689130
rect 119090 688890 119180 689130
rect 119420 688890 119510 689130
rect 119750 688890 119840 689130
rect 120080 688890 120190 689130
rect 120430 688890 120520 689130
rect 120760 688890 120850 689130
rect 121090 688890 121180 689130
rect 121420 688890 121530 689130
rect 121770 688890 121790 689130
rect 110790 688800 121790 688890
rect 110790 688560 110810 688800
rect 111050 688560 111140 688800
rect 111380 688560 111470 688800
rect 111710 688560 111800 688800
rect 112040 688560 112150 688800
rect 112390 688560 112480 688800
rect 112720 688560 112810 688800
rect 113050 688560 113140 688800
rect 113380 688560 113490 688800
rect 113730 688560 113820 688800
rect 114060 688560 114150 688800
rect 114390 688560 114480 688800
rect 114720 688560 114830 688800
rect 115070 688560 115160 688800
rect 115400 688560 115490 688800
rect 115730 688560 115820 688800
rect 116060 688560 116170 688800
rect 116410 688560 116500 688800
rect 116740 688560 116830 688800
rect 117070 688560 117160 688800
rect 117400 688560 117510 688800
rect 117750 688560 117840 688800
rect 118080 688560 118170 688800
rect 118410 688560 118500 688800
rect 118740 688560 118850 688800
rect 119090 688560 119180 688800
rect 119420 688560 119510 688800
rect 119750 688560 119840 688800
rect 120080 688560 120190 688800
rect 120430 688560 120520 688800
rect 120760 688560 120850 688800
rect 121090 688560 121180 688800
rect 121420 688560 121530 688800
rect 121770 688560 121790 688800
rect 110790 688470 121790 688560
rect 110790 688230 110810 688470
rect 111050 688230 111140 688470
rect 111380 688230 111470 688470
rect 111710 688230 111800 688470
rect 112040 688230 112150 688470
rect 112390 688230 112480 688470
rect 112720 688230 112810 688470
rect 113050 688230 113140 688470
rect 113380 688230 113490 688470
rect 113730 688230 113820 688470
rect 114060 688230 114150 688470
rect 114390 688230 114480 688470
rect 114720 688230 114830 688470
rect 115070 688230 115160 688470
rect 115400 688230 115490 688470
rect 115730 688230 115820 688470
rect 116060 688230 116170 688470
rect 116410 688230 116500 688470
rect 116740 688230 116830 688470
rect 117070 688230 117160 688470
rect 117400 688230 117510 688470
rect 117750 688230 117840 688470
rect 118080 688230 118170 688470
rect 118410 688230 118500 688470
rect 118740 688230 118850 688470
rect 119090 688230 119180 688470
rect 119420 688230 119510 688470
rect 119750 688230 119840 688470
rect 120080 688230 120190 688470
rect 120430 688230 120520 688470
rect 120760 688230 120850 688470
rect 121090 688230 121180 688470
rect 121420 688230 121530 688470
rect 121770 688230 121790 688470
rect 110790 688140 121790 688230
rect 110790 687900 110810 688140
rect 111050 687900 111140 688140
rect 111380 687900 111470 688140
rect 111710 687900 111800 688140
rect 112040 687900 112150 688140
rect 112390 687900 112480 688140
rect 112720 687900 112810 688140
rect 113050 687900 113140 688140
rect 113380 687900 113490 688140
rect 113730 687900 113820 688140
rect 114060 687900 114150 688140
rect 114390 687900 114480 688140
rect 114720 687900 114830 688140
rect 115070 687900 115160 688140
rect 115400 687900 115490 688140
rect 115730 687900 115820 688140
rect 116060 687900 116170 688140
rect 116410 687900 116500 688140
rect 116740 687900 116830 688140
rect 117070 687900 117160 688140
rect 117400 687900 117510 688140
rect 117750 687900 117840 688140
rect 118080 687900 118170 688140
rect 118410 687900 118500 688140
rect 118740 687900 118850 688140
rect 119090 687900 119180 688140
rect 119420 687900 119510 688140
rect 119750 687900 119840 688140
rect 120080 687900 120190 688140
rect 120430 687900 120520 688140
rect 120760 687900 120850 688140
rect 121090 687900 121180 688140
rect 121420 687900 121530 688140
rect 121770 687900 121790 688140
rect 110790 687790 121790 687900
rect 110790 687550 110810 687790
rect 111050 687550 111140 687790
rect 111380 687550 111470 687790
rect 111710 687550 111800 687790
rect 112040 687550 112150 687790
rect 112390 687550 112480 687790
rect 112720 687550 112810 687790
rect 113050 687550 113140 687790
rect 113380 687550 113490 687790
rect 113730 687550 113820 687790
rect 114060 687550 114150 687790
rect 114390 687550 114480 687790
rect 114720 687550 114830 687790
rect 115070 687550 115160 687790
rect 115400 687550 115490 687790
rect 115730 687550 115820 687790
rect 116060 687550 116170 687790
rect 116410 687550 116500 687790
rect 116740 687550 116830 687790
rect 117070 687550 117160 687790
rect 117400 687550 117510 687790
rect 117750 687550 117840 687790
rect 118080 687550 118170 687790
rect 118410 687550 118500 687790
rect 118740 687550 118850 687790
rect 119090 687550 119180 687790
rect 119420 687550 119510 687790
rect 119750 687550 119840 687790
rect 120080 687550 120190 687790
rect 120430 687550 120520 687790
rect 120760 687550 120850 687790
rect 121090 687550 121180 687790
rect 121420 687550 121530 687790
rect 121770 687550 121790 687790
rect 110790 687460 121790 687550
rect 110790 687220 110810 687460
rect 111050 687220 111140 687460
rect 111380 687220 111470 687460
rect 111710 687220 111800 687460
rect 112040 687220 112150 687460
rect 112390 687220 112480 687460
rect 112720 687220 112810 687460
rect 113050 687220 113140 687460
rect 113380 687220 113490 687460
rect 113730 687220 113820 687460
rect 114060 687220 114150 687460
rect 114390 687220 114480 687460
rect 114720 687220 114830 687460
rect 115070 687220 115160 687460
rect 115400 687220 115490 687460
rect 115730 687220 115820 687460
rect 116060 687220 116170 687460
rect 116410 687220 116500 687460
rect 116740 687220 116830 687460
rect 117070 687220 117160 687460
rect 117400 687220 117510 687460
rect 117750 687220 117840 687460
rect 118080 687220 118170 687460
rect 118410 687220 118500 687460
rect 118740 687220 118850 687460
rect 119090 687220 119180 687460
rect 119420 687220 119510 687460
rect 119750 687220 119840 687460
rect 120080 687220 120190 687460
rect 120430 687220 120520 687460
rect 120760 687220 120850 687460
rect 121090 687220 121180 687460
rect 121420 687220 121530 687460
rect 121770 687220 121790 687460
rect 110790 687130 121790 687220
rect 110790 686890 110810 687130
rect 111050 686890 111140 687130
rect 111380 686890 111470 687130
rect 111710 686890 111800 687130
rect 112040 686890 112150 687130
rect 112390 686890 112480 687130
rect 112720 686890 112810 687130
rect 113050 686890 113140 687130
rect 113380 686890 113490 687130
rect 113730 686890 113820 687130
rect 114060 686890 114150 687130
rect 114390 686890 114480 687130
rect 114720 686890 114830 687130
rect 115070 686890 115160 687130
rect 115400 686890 115490 687130
rect 115730 686890 115820 687130
rect 116060 686890 116170 687130
rect 116410 686890 116500 687130
rect 116740 686890 116830 687130
rect 117070 686890 117160 687130
rect 117400 686890 117510 687130
rect 117750 686890 117840 687130
rect 118080 686890 118170 687130
rect 118410 686890 118500 687130
rect 118740 686890 118850 687130
rect 119090 686890 119180 687130
rect 119420 686890 119510 687130
rect 119750 686890 119840 687130
rect 120080 686890 120190 687130
rect 120430 686890 120520 687130
rect 120760 686890 120850 687130
rect 121090 686890 121180 687130
rect 121420 686890 121530 687130
rect 121770 686890 121790 687130
rect 110790 686800 121790 686890
rect 110790 686560 110810 686800
rect 111050 686560 111140 686800
rect 111380 686560 111470 686800
rect 111710 686560 111800 686800
rect 112040 686560 112150 686800
rect 112390 686560 112480 686800
rect 112720 686560 112810 686800
rect 113050 686560 113140 686800
rect 113380 686560 113490 686800
rect 113730 686560 113820 686800
rect 114060 686560 114150 686800
rect 114390 686560 114480 686800
rect 114720 686560 114830 686800
rect 115070 686560 115160 686800
rect 115400 686560 115490 686800
rect 115730 686560 115820 686800
rect 116060 686560 116170 686800
rect 116410 686560 116500 686800
rect 116740 686560 116830 686800
rect 117070 686560 117160 686800
rect 117400 686560 117510 686800
rect 117750 686560 117840 686800
rect 118080 686560 118170 686800
rect 118410 686560 118500 686800
rect 118740 686560 118850 686800
rect 119090 686560 119180 686800
rect 119420 686560 119510 686800
rect 119750 686560 119840 686800
rect 120080 686560 120190 686800
rect 120430 686560 120520 686800
rect 120760 686560 120850 686800
rect 121090 686560 121180 686800
rect 121420 686560 121530 686800
rect 121770 686560 121790 686800
rect 110790 686450 121790 686560
rect 110790 686210 110810 686450
rect 111050 686210 111140 686450
rect 111380 686210 111470 686450
rect 111710 686210 111800 686450
rect 112040 686210 112150 686450
rect 112390 686210 112480 686450
rect 112720 686210 112810 686450
rect 113050 686210 113140 686450
rect 113380 686210 113490 686450
rect 113730 686210 113820 686450
rect 114060 686210 114150 686450
rect 114390 686210 114480 686450
rect 114720 686210 114830 686450
rect 115070 686210 115160 686450
rect 115400 686210 115490 686450
rect 115730 686210 115820 686450
rect 116060 686210 116170 686450
rect 116410 686210 116500 686450
rect 116740 686210 116830 686450
rect 117070 686210 117160 686450
rect 117400 686210 117510 686450
rect 117750 686210 117840 686450
rect 118080 686210 118170 686450
rect 118410 686210 118500 686450
rect 118740 686210 118850 686450
rect 119090 686210 119180 686450
rect 119420 686210 119510 686450
rect 119750 686210 119840 686450
rect 120080 686210 120190 686450
rect 120430 686210 120520 686450
rect 120760 686210 120850 686450
rect 121090 686210 121180 686450
rect 121420 686210 121530 686450
rect 121770 686210 121790 686450
rect 110790 686120 121790 686210
rect 110790 685880 110810 686120
rect 111050 685880 111140 686120
rect 111380 685880 111470 686120
rect 111710 685880 111800 686120
rect 112040 685880 112150 686120
rect 112390 685880 112480 686120
rect 112720 685880 112810 686120
rect 113050 685880 113140 686120
rect 113380 685880 113490 686120
rect 113730 685880 113820 686120
rect 114060 685880 114150 686120
rect 114390 685880 114480 686120
rect 114720 685880 114830 686120
rect 115070 685880 115160 686120
rect 115400 685880 115490 686120
rect 115730 685880 115820 686120
rect 116060 685880 116170 686120
rect 116410 685880 116500 686120
rect 116740 685880 116830 686120
rect 117070 685880 117160 686120
rect 117400 685880 117510 686120
rect 117750 685880 117840 686120
rect 118080 685880 118170 686120
rect 118410 685880 118500 686120
rect 118740 685880 118850 686120
rect 119090 685880 119180 686120
rect 119420 685880 119510 686120
rect 119750 685880 119840 686120
rect 120080 685880 120190 686120
rect 120430 685880 120520 686120
rect 120760 685880 120850 686120
rect 121090 685880 121180 686120
rect 121420 685880 121530 686120
rect 121770 685880 121790 686120
rect 110790 685790 121790 685880
rect 110790 685550 110810 685790
rect 111050 685550 111140 685790
rect 111380 685550 111470 685790
rect 111710 685550 111800 685790
rect 112040 685550 112150 685790
rect 112390 685550 112480 685790
rect 112720 685550 112810 685790
rect 113050 685550 113140 685790
rect 113380 685550 113490 685790
rect 113730 685550 113820 685790
rect 114060 685550 114150 685790
rect 114390 685550 114480 685790
rect 114720 685550 114830 685790
rect 115070 685550 115160 685790
rect 115400 685550 115490 685790
rect 115730 685550 115820 685790
rect 116060 685550 116170 685790
rect 116410 685550 116500 685790
rect 116740 685550 116830 685790
rect 117070 685550 117160 685790
rect 117400 685550 117510 685790
rect 117750 685550 117840 685790
rect 118080 685550 118170 685790
rect 118410 685550 118500 685790
rect 118740 685550 118850 685790
rect 119090 685550 119180 685790
rect 119420 685550 119510 685790
rect 119750 685550 119840 685790
rect 120080 685550 120190 685790
rect 120430 685550 120520 685790
rect 120760 685550 120850 685790
rect 121090 685550 121180 685790
rect 121420 685550 121530 685790
rect 121770 685550 121790 685790
rect 110790 685460 121790 685550
rect 110790 685220 110810 685460
rect 111050 685220 111140 685460
rect 111380 685220 111470 685460
rect 111710 685220 111800 685460
rect 112040 685220 112150 685460
rect 112390 685220 112480 685460
rect 112720 685220 112810 685460
rect 113050 685220 113140 685460
rect 113380 685220 113490 685460
rect 113730 685220 113820 685460
rect 114060 685220 114150 685460
rect 114390 685220 114480 685460
rect 114720 685220 114830 685460
rect 115070 685220 115160 685460
rect 115400 685220 115490 685460
rect 115730 685220 115820 685460
rect 116060 685220 116170 685460
rect 116410 685220 116500 685460
rect 116740 685220 116830 685460
rect 117070 685220 117160 685460
rect 117400 685220 117510 685460
rect 117750 685220 117840 685460
rect 118080 685220 118170 685460
rect 118410 685220 118500 685460
rect 118740 685220 118850 685460
rect 119090 685220 119180 685460
rect 119420 685220 119510 685460
rect 119750 685220 119840 685460
rect 120080 685220 120190 685460
rect 120430 685220 120520 685460
rect 120760 685220 120850 685460
rect 121090 685220 121180 685460
rect 121420 685220 121530 685460
rect 121770 685220 121790 685460
rect 110790 685110 121790 685220
rect 110790 684870 110810 685110
rect 111050 684870 111140 685110
rect 111380 684870 111470 685110
rect 111710 684870 111800 685110
rect 112040 684870 112150 685110
rect 112390 684870 112480 685110
rect 112720 684870 112810 685110
rect 113050 684870 113140 685110
rect 113380 684870 113490 685110
rect 113730 684870 113820 685110
rect 114060 684870 114150 685110
rect 114390 684870 114480 685110
rect 114720 684870 114830 685110
rect 115070 684870 115160 685110
rect 115400 684870 115490 685110
rect 115730 684870 115820 685110
rect 116060 684870 116170 685110
rect 116410 684870 116500 685110
rect 116740 684870 116830 685110
rect 117070 684870 117160 685110
rect 117400 684870 117510 685110
rect 117750 684870 117840 685110
rect 118080 684870 118170 685110
rect 118410 684870 118500 685110
rect 118740 684870 118850 685110
rect 119090 684870 119180 685110
rect 119420 684870 119510 685110
rect 119750 684870 119840 685110
rect 120080 684870 120190 685110
rect 120430 684870 120520 685110
rect 120760 684870 120850 685110
rect 121090 684870 121180 685110
rect 121420 684870 121530 685110
rect 121770 684870 121790 685110
rect 110790 684780 121790 684870
rect 110790 684540 110810 684780
rect 111050 684540 111140 684780
rect 111380 684540 111470 684780
rect 111710 684540 111800 684780
rect 112040 684540 112150 684780
rect 112390 684540 112480 684780
rect 112720 684540 112810 684780
rect 113050 684540 113140 684780
rect 113380 684540 113490 684780
rect 113730 684540 113820 684780
rect 114060 684540 114150 684780
rect 114390 684540 114480 684780
rect 114720 684540 114830 684780
rect 115070 684540 115160 684780
rect 115400 684540 115490 684780
rect 115730 684540 115820 684780
rect 116060 684540 116170 684780
rect 116410 684540 116500 684780
rect 116740 684540 116830 684780
rect 117070 684540 117160 684780
rect 117400 684540 117510 684780
rect 117750 684540 117840 684780
rect 118080 684540 118170 684780
rect 118410 684540 118500 684780
rect 118740 684540 118850 684780
rect 119090 684540 119180 684780
rect 119420 684540 119510 684780
rect 119750 684540 119840 684780
rect 120080 684540 120190 684780
rect 120430 684540 120520 684780
rect 120760 684540 120850 684780
rect 121090 684540 121180 684780
rect 121420 684540 121530 684780
rect 121770 684540 121790 684780
rect 110790 684450 121790 684540
rect 110790 684210 110810 684450
rect 111050 684210 111140 684450
rect 111380 684210 111470 684450
rect 111710 684210 111800 684450
rect 112040 684210 112150 684450
rect 112390 684210 112480 684450
rect 112720 684210 112810 684450
rect 113050 684210 113140 684450
rect 113380 684210 113490 684450
rect 113730 684210 113820 684450
rect 114060 684210 114150 684450
rect 114390 684210 114480 684450
rect 114720 684210 114830 684450
rect 115070 684210 115160 684450
rect 115400 684210 115490 684450
rect 115730 684210 115820 684450
rect 116060 684210 116170 684450
rect 116410 684210 116500 684450
rect 116740 684210 116830 684450
rect 117070 684210 117160 684450
rect 117400 684210 117510 684450
rect 117750 684210 117840 684450
rect 118080 684210 118170 684450
rect 118410 684210 118500 684450
rect 118740 684210 118850 684450
rect 119090 684210 119180 684450
rect 119420 684210 119510 684450
rect 119750 684210 119840 684450
rect 120080 684210 120190 684450
rect 120430 684210 120520 684450
rect 120760 684210 120850 684450
rect 121090 684210 121180 684450
rect 121420 684210 121530 684450
rect 121770 684210 121790 684450
rect 110790 684120 121790 684210
rect 110790 683880 110810 684120
rect 111050 683880 111140 684120
rect 111380 683880 111470 684120
rect 111710 683880 111800 684120
rect 112040 683880 112150 684120
rect 112390 683880 112480 684120
rect 112720 683880 112810 684120
rect 113050 683880 113140 684120
rect 113380 683880 113490 684120
rect 113730 683880 113820 684120
rect 114060 683880 114150 684120
rect 114390 683880 114480 684120
rect 114720 683880 114830 684120
rect 115070 683880 115160 684120
rect 115400 683880 115490 684120
rect 115730 683880 115820 684120
rect 116060 683880 116170 684120
rect 116410 683880 116500 684120
rect 116740 683880 116830 684120
rect 117070 683880 117160 684120
rect 117400 683880 117510 684120
rect 117750 683880 117840 684120
rect 118080 683880 118170 684120
rect 118410 683880 118500 684120
rect 118740 683880 118850 684120
rect 119090 683880 119180 684120
rect 119420 683880 119510 684120
rect 119750 683880 119840 684120
rect 120080 683880 120190 684120
rect 120430 683880 120520 684120
rect 120760 683880 120850 684120
rect 121090 683880 121180 684120
rect 121420 683880 121530 684120
rect 121770 683880 121790 684120
rect 110790 683860 121790 683880
rect 122170 694840 133170 694860
rect 122170 694600 122190 694840
rect 122430 694600 122520 694840
rect 122760 694600 122850 694840
rect 123090 694600 123180 694840
rect 123420 694600 123530 694840
rect 123770 694600 123860 694840
rect 124100 694600 124190 694840
rect 124430 694600 124520 694840
rect 124760 694600 124870 694840
rect 125110 694600 125200 694840
rect 125440 694600 125530 694840
rect 125770 694600 125860 694840
rect 126100 694600 126210 694840
rect 126450 694600 126540 694840
rect 126780 694600 126870 694840
rect 127110 694600 127200 694840
rect 127440 694600 127550 694840
rect 127790 694600 127880 694840
rect 128120 694600 128210 694840
rect 128450 694600 128540 694840
rect 128780 694600 128890 694840
rect 129130 694600 129220 694840
rect 129460 694600 129550 694840
rect 129790 694600 129880 694840
rect 130120 694600 130230 694840
rect 130470 694600 130560 694840
rect 130800 694600 130890 694840
rect 131130 694600 131220 694840
rect 131460 694600 131570 694840
rect 131810 694600 131900 694840
rect 132140 694600 132230 694840
rect 132470 694600 132560 694840
rect 132800 694600 132910 694840
rect 133150 694600 133170 694840
rect 122170 694490 133170 694600
rect 122170 694250 122190 694490
rect 122430 694250 122520 694490
rect 122760 694250 122850 694490
rect 123090 694250 123180 694490
rect 123420 694250 123530 694490
rect 123770 694250 123860 694490
rect 124100 694250 124190 694490
rect 124430 694250 124520 694490
rect 124760 694250 124870 694490
rect 125110 694250 125200 694490
rect 125440 694250 125530 694490
rect 125770 694250 125860 694490
rect 126100 694250 126210 694490
rect 126450 694250 126540 694490
rect 126780 694250 126870 694490
rect 127110 694250 127200 694490
rect 127440 694250 127550 694490
rect 127790 694250 127880 694490
rect 128120 694250 128210 694490
rect 128450 694250 128540 694490
rect 128780 694250 128890 694490
rect 129130 694250 129220 694490
rect 129460 694250 129550 694490
rect 129790 694250 129880 694490
rect 130120 694250 130230 694490
rect 130470 694250 130560 694490
rect 130800 694250 130890 694490
rect 131130 694250 131220 694490
rect 131460 694250 131570 694490
rect 131810 694250 131900 694490
rect 132140 694250 132230 694490
rect 132470 694250 132560 694490
rect 132800 694250 132910 694490
rect 133150 694250 133170 694490
rect 122170 694160 133170 694250
rect 122170 693920 122190 694160
rect 122430 693920 122520 694160
rect 122760 693920 122850 694160
rect 123090 693920 123180 694160
rect 123420 693920 123530 694160
rect 123770 693920 123860 694160
rect 124100 693920 124190 694160
rect 124430 693920 124520 694160
rect 124760 693920 124870 694160
rect 125110 693920 125200 694160
rect 125440 693920 125530 694160
rect 125770 693920 125860 694160
rect 126100 693920 126210 694160
rect 126450 693920 126540 694160
rect 126780 693920 126870 694160
rect 127110 693920 127200 694160
rect 127440 693920 127550 694160
rect 127790 693920 127880 694160
rect 128120 693920 128210 694160
rect 128450 693920 128540 694160
rect 128780 693920 128890 694160
rect 129130 693920 129220 694160
rect 129460 693920 129550 694160
rect 129790 693920 129880 694160
rect 130120 693920 130230 694160
rect 130470 693920 130560 694160
rect 130800 693920 130890 694160
rect 131130 693920 131220 694160
rect 131460 693920 131570 694160
rect 131810 693920 131900 694160
rect 132140 693920 132230 694160
rect 132470 693920 132560 694160
rect 132800 693920 132910 694160
rect 133150 693920 133170 694160
rect 122170 693830 133170 693920
rect 122170 693590 122190 693830
rect 122430 693590 122520 693830
rect 122760 693590 122850 693830
rect 123090 693590 123180 693830
rect 123420 693590 123530 693830
rect 123770 693590 123860 693830
rect 124100 693590 124190 693830
rect 124430 693590 124520 693830
rect 124760 693590 124870 693830
rect 125110 693590 125200 693830
rect 125440 693590 125530 693830
rect 125770 693590 125860 693830
rect 126100 693590 126210 693830
rect 126450 693590 126540 693830
rect 126780 693590 126870 693830
rect 127110 693590 127200 693830
rect 127440 693590 127550 693830
rect 127790 693590 127880 693830
rect 128120 693590 128210 693830
rect 128450 693590 128540 693830
rect 128780 693590 128890 693830
rect 129130 693590 129220 693830
rect 129460 693590 129550 693830
rect 129790 693590 129880 693830
rect 130120 693590 130230 693830
rect 130470 693590 130560 693830
rect 130800 693590 130890 693830
rect 131130 693590 131220 693830
rect 131460 693590 131570 693830
rect 131810 693590 131900 693830
rect 132140 693590 132230 693830
rect 132470 693590 132560 693830
rect 132800 693590 132910 693830
rect 133150 693590 133170 693830
rect 122170 693500 133170 693590
rect 122170 693260 122190 693500
rect 122430 693260 122520 693500
rect 122760 693260 122850 693500
rect 123090 693260 123180 693500
rect 123420 693260 123530 693500
rect 123770 693260 123860 693500
rect 124100 693260 124190 693500
rect 124430 693260 124520 693500
rect 124760 693260 124870 693500
rect 125110 693260 125200 693500
rect 125440 693260 125530 693500
rect 125770 693260 125860 693500
rect 126100 693260 126210 693500
rect 126450 693260 126540 693500
rect 126780 693260 126870 693500
rect 127110 693260 127200 693500
rect 127440 693260 127550 693500
rect 127790 693260 127880 693500
rect 128120 693260 128210 693500
rect 128450 693260 128540 693500
rect 128780 693260 128890 693500
rect 129130 693260 129220 693500
rect 129460 693260 129550 693500
rect 129790 693260 129880 693500
rect 130120 693260 130230 693500
rect 130470 693260 130560 693500
rect 130800 693260 130890 693500
rect 131130 693260 131220 693500
rect 131460 693260 131570 693500
rect 131810 693260 131900 693500
rect 132140 693260 132230 693500
rect 132470 693260 132560 693500
rect 132800 693260 132910 693500
rect 133150 693260 133170 693500
rect 122170 693150 133170 693260
rect 122170 692910 122190 693150
rect 122430 692910 122520 693150
rect 122760 692910 122850 693150
rect 123090 692910 123180 693150
rect 123420 692910 123530 693150
rect 123770 692910 123860 693150
rect 124100 692910 124190 693150
rect 124430 692910 124520 693150
rect 124760 692910 124870 693150
rect 125110 692910 125200 693150
rect 125440 692910 125530 693150
rect 125770 692910 125860 693150
rect 126100 692910 126210 693150
rect 126450 692910 126540 693150
rect 126780 692910 126870 693150
rect 127110 692910 127200 693150
rect 127440 692910 127550 693150
rect 127790 692910 127880 693150
rect 128120 692910 128210 693150
rect 128450 692910 128540 693150
rect 128780 692910 128890 693150
rect 129130 692910 129220 693150
rect 129460 692910 129550 693150
rect 129790 692910 129880 693150
rect 130120 692910 130230 693150
rect 130470 692910 130560 693150
rect 130800 692910 130890 693150
rect 131130 692910 131220 693150
rect 131460 692910 131570 693150
rect 131810 692910 131900 693150
rect 132140 692910 132230 693150
rect 132470 692910 132560 693150
rect 132800 692910 132910 693150
rect 133150 692910 133170 693150
rect 122170 692820 133170 692910
rect 122170 692580 122190 692820
rect 122430 692580 122520 692820
rect 122760 692580 122850 692820
rect 123090 692580 123180 692820
rect 123420 692580 123530 692820
rect 123770 692580 123860 692820
rect 124100 692580 124190 692820
rect 124430 692580 124520 692820
rect 124760 692580 124870 692820
rect 125110 692580 125200 692820
rect 125440 692580 125530 692820
rect 125770 692580 125860 692820
rect 126100 692580 126210 692820
rect 126450 692580 126540 692820
rect 126780 692580 126870 692820
rect 127110 692580 127200 692820
rect 127440 692580 127550 692820
rect 127790 692580 127880 692820
rect 128120 692580 128210 692820
rect 128450 692580 128540 692820
rect 128780 692580 128890 692820
rect 129130 692580 129220 692820
rect 129460 692580 129550 692820
rect 129790 692580 129880 692820
rect 130120 692580 130230 692820
rect 130470 692580 130560 692820
rect 130800 692580 130890 692820
rect 131130 692580 131220 692820
rect 131460 692580 131570 692820
rect 131810 692580 131900 692820
rect 132140 692580 132230 692820
rect 132470 692580 132560 692820
rect 132800 692580 132910 692820
rect 133150 692580 133170 692820
rect 122170 692490 133170 692580
rect 122170 692250 122190 692490
rect 122430 692250 122520 692490
rect 122760 692250 122850 692490
rect 123090 692250 123180 692490
rect 123420 692250 123530 692490
rect 123770 692250 123860 692490
rect 124100 692250 124190 692490
rect 124430 692250 124520 692490
rect 124760 692250 124870 692490
rect 125110 692250 125200 692490
rect 125440 692250 125530 692490
rect 125770 692250 125860 692490
rect 126100 692250 126210 692490
rect 126450 692250 126540 692490
rect 126780 692250 126870 692490
rect 127110 692250 127200 692490
rect 127440 692250 127550 692490
rect 127790 692250 127880 692490
rect 128120 692250 128210 692490
rect 128450 692250 128540 692490
rect 128780 692250 128890 692490
rect 129130 692250 129220 692490
rect 129460 692250 129550 692490
rect 129790 692250 129880 692490
rect 130120 692250 130230 692490
rect 130470 692250 130560 692490
rect 130800 692250 130890 692490
rect 131130 692250 131220 692490
rect 131460 692250 131570 692490
rect 131810 692250 131900 692490
rect 132140 692250 132230 692490
rect 132470 692250 132560 692490
rect 132800 692250 132910 692490
rect 133150 692250 133170 692490
rect 122170 692160 133170 692250
rect 122170 691920 122190 692160
rect 122430 691920 122520 692160
rect 122760 691920 122850 692160
rect 123090 691920 123180 692160
rect 123420 691920 123530 692160
rect 123770 691920 123860 692160
rect 124100 691920 124190 692160
rect 124430 691920 124520 692160
rect 124760 691920 124870 692160
rect 125110 691920 125200 692160
rect 125440 691920 125530 692160
rect 125770 691920 125860 692160
rect 126100 691920 126210 692160
rect 126450 691920 126540 692160
rect 126780 691920 126870 692160
rect 127110 691920 127200 692160
rect 127440 691920 127550 692160
rect 127790 691920 127880 692160
rect 128120 691920 128210 692160
rect 128450 691920 128540 692160
rect 128780 691920 128890 692160
rect 129130 691920 129220 692160
rect 129460 691920 129550 692160
rect 129790 691920 129880 692160
rect 130120 691920 130230 692160
rect 130470 691920 130560 692160
rect 130800 691920 130890 692160
rect 131130 691920 131220 692160
rect 131460 691920 131570 692160
rect 131810 691920 131900 692160
rect 132140 691920 132230 692160
rect 132470 691920 132560 692160
rect 132800 691920 132910 692160
rect 133150 691920 133170 692160
rect 122170 691810 133170 691920
rect 122170 691570 122190 691810
rect 122430 691570 122520 691810
rect 122760 691570 122850 691810
rect 123090 691570 123180 691810
rect 123420 691570 123530 691810
rect 123770 691570 123860 691810
rect 124100 691570 124190 691810
rect 124430 691570 124520 691810
rect 124760 691570 124870 691810
rect 125110 691570 125200 691810
rect 125440 691570 125530 691810
rect 125770 691570 125860 691810
rect 126100 691570 126210 691810
rect 126450 691570 126540 691810
rect 126780 691570 126870 691810
rect 127110 691570 127200 691810
rect 127440 691570 127550 691810
rect 127790 691570 127880 691810
rect 128120 691570 128210 691810
rect 128450 691570 128540 691810
rect 128780 691570 128890 691810
rect 129130 691570 129220 691810
rect 129460 691570 129550 691810
rect 129790 691570 129880 691810
rect 130120 691570 130230 691810
rect 130470 691570 130560 691810
rect 130800 691570 130890 691810
rect 131130 691570 131220 691810
rect 131460 691570 131570 691810
rect 131810 691570 131900 691810
rect 132140 691570 132230 691810
rect 132470 691570 132560 691810
rect 132800 691570 132910 691810
rect 133150 691570 133170 691810
rect 122170 691480 133170 691570
rect 122170 691240 122190 691480
rect 122430 691240 122520 691480
rect 122760 691240 122850 691480
rect 123090 691240 123180 691480
rect 123420 691240 123530 691480
rect 123770 691240 123860 691480
rect 124100 691240 124190 691480
rect 124430 691240 124520 691480
rect 124760 691240 124870 691480
rect 125110 691240 125200 691480
rect 125440 691240 125530 691480
rect 125770 691240 125860 691480
rect 126100 691240 126210 691480
rect 126450 691240 126540 691480
rect 126780 691240 126870 691480
rect 127110 691240 127200 691480
rect 127440 691240 127550 691480
rect 127790 691240 127880 691480
rect 128120 691240 128210 691480
rect 128450 691240 128540 691480
rect 128780 691240 128890 691480
rect 129130 691240 129220 691480
rect 129460 691240 129550 691480
rect 129790 691240 129880 691480
rect 130120 691240 130230 691480
rect 130470 691240 130560 691480
rect 130800 691240 130890 691480
rect 131130 691240 131220 691480
rect 131460 691240 131570 691480
rect 131810 691240 131900 691480
rect 132140 691240 132230 691480
rect 132470 691240 132560 691480
rect 132800 691240 132910 691480
rect 133150 691240 133170 691480
rect 122170 691150 133170 691240
rect 122170 690910 122190 691150
rect 122430 690910 122520 691150
rect 122760 690910 122850 691150
rect 123090 690910 123180 691150
rect 123420 690910 123530 691150
rect 123770 690910 123860 691150
rect 124100 690910 124190 691150
rect 124430 690910 124520 691150
rect 124760 690910 124870 691150
rect 125110 690910 125200 691150
rect 125440 690910 125530 691150
rect 125770 690910 125860 691150
rect 126100 690910 126210 691150
rect 126450 690910 126540 691150
rect 126780 690910 126870 691150
rect 127110 690910 127200 691150
rect 127440 690910 127550 691150
rect 127790 690910 127880 691150
rect 128120 690910 128210 691150
rect 128450 690910 128540 691150
rect 128780 690910 128890 691150
rect 129130 690910 129220 691150
rect 129460 690910 129550 691150
rect 129790 690910 129880 691150
rect 130120 690910 130230 691150
rect 130470 690910 130560 691150
rect 130800 690910 130890 691150
rect 131130 690910 131220 691150
rect 131460 690910 131570 691150
rect 131810 690910 131900 691150
rect 132140 690910 132230 691150
rect 132470 690910 132560 691150
rect 132800 690910 132910 691150
rect 133150 690910 133170 691150
rect 122170 690820 133170 690910
rect 122170 690580 122190 690820
rect 122430 690580 122520 690820
rect 122760 690580 122850 690820
rect 123090 690580 123180 690820
rect 123420 690580 123530 690820
rect 123770 690580 123860 690820
rect 124100 690580 124190 690820
rect 124430 690580 124520 690820
rect 124760 690580 124870 690820
rect 125110 690580 125200 690820
rect 125440 690580 125530 690820
rect 125770 690580 125860 690820
rect 126100 690580 126210 690820
rect 126450 690580 126540 690820
rect 126780 690580 126870 690820
rect 127110 690580 127200 690820
rect 127440 690580 127550 690820
rect 127790 690580 127880 690820
rect 128120 690580 128210 690820
rect 128450 690580 128540 690820
rect 128780 690580 128890 690820
rect 129130 690580 129220 690820
rect 129460 690580 129550 690820
rect 129790 690580 129880 690820
rect 130120 690580 130230 690820
rect 130470 690580 130560 690820
rect 130800 690580 130890 690820
rect 131130 690580 131220 690820
rect 131460 690580 131570 690820
rect 131810 690580 131900 690820
rect 132140 690580 132230 690820
rect 132470 690580 132560 690820
rect 132800 690580 132910 690820
rect 133150 690580 133170 690820
rect 122170 690470 133170 690580
rect 122170 690230 122190 690470
rect 122430 690230 122520 690470
rect 122760 690230 122850 690470
rect 123090 690230 123180 690470
rect 123420 690230 123530 690470
rect 123770 690230 123860 690470
rect 124100 690230 124190 690470
rect 124430 690230 124520 690470
rect 124760 690230 124870 690470
rect 125110 690230 125200 690470
rect 125440 690230 125530 690470
rect 125770 690230 125860 690470
rect 126100 690230 126210 690470
rect 126450 690230 126540 690470
rect 126780 690230 126870 690470
rect 127110 690230 127200 690470
rect 127440 690230 127550 690470
rect 127790 690230 127880 690470
rect 128120 690230 128210 690470
rect 128450 690230 128540 690470
rect 128780 690230 128890 690470
rect 129130 690230 129220 690470
rect 129460 690230 129550 690470
rect 129790 690230 129880 690470
rect 130120 690230 130230 690470
rect 130470 690230 130560 690470
rect 130800 690230 130890 690470
rect 131130 690230 131220 690470
rect 131460 690230 131570 690470
rect 131810 690230 131900 690470
rect 132140 690230 132230 690470
rect 132470 690230 132560 690470
rect 132800 690230 132910 690470
rect 133150 690230 133170 690470
rect 122170 690140 133170 690230
rect 122170 689900 122190 690140
rect 122430 689900 122520 690140
rect 122760 689900 122850 690140
rect 123090 689900 123180 690140
rect 123420 689900 123530 690140
rect 123770 689900 123860 690140
rect 124100 689900 124190 690140
rect 124430 689900 124520 690140
rect 124760 689900 124870 690140
rect 125110 689900 125200 690140
rect 125440 689900 125530 690140
rect 125770 689900 125860 690140
rect 126100 689900 126210 690140
rect 126450 689900 126540 690140
rect 126780 689900 126870 690140
rect 127110 689900 127200 690140
rect 127440 689900 127550 690140
rect 127790 689900 127880 690140
rect 128120 689900 128210 690140
rect 128450 689900 128540 690140
rect 128780 689900 128890 690140
rect 129130 689900 129220 690140
rect 129460 689900 129550 690140
rect 129790 689900 129880 690140
rect 130120 689900 130230 690140
rect 130470 689900 130560 690140
rect 130800 689900 130890 690140
rect 131130 689900 131220 690140
rect 131460 689900 131570 690140
rect 131810 689900 131900 690140
rect 132140 689900 132230 690140
rect 132470 689900 132560 690140
rect 132800 689900 132910 690140
rect 133150 689900 133170 690140
rect 122170 689810 133170 689900
rect 122170 689570 122190 689810
rect 122430 689570 122520 689810
rect 122760 689570 122850 689810
rect 123090 689570 123180 689810
rect 123420 689570 123530 689810
rect 123770 689570 123860 689810
rect 124100 689570 124190 689810
rect 124430 689570 124520 689810
rect 124760 689570 124870 689810
rect 125110 689570 125200 689810
rect 125440 689570 125530 689810
rect 125770 689570 125860 689810
rect 126100 689570 126210 689810
rect 126450 689570 126540 689810
rect 126780 689570 126870 689810
rect 127110 689570 127200 689810
rect 127440 689570 127550 689810
rect 127790 689570 127880 689810
rect 128120 689570 128210 689810
rect 128450 689570 128540 689810
rect 128780 689570 128890 689810
rect 129130 689570 129220 689810
rect 129460 689570 129550 689810
rect 129790 689570 129880 689810
rect 130120 689570 130230 689810
rect 130470 689570 130560 689810
rect 130800 689570 130890 689810
rect 131130 689570 131220 689810
rect 131460 689570 131570 689810
rect 131810 689570 131900 689810
rect 132140 689570 132230 689810
rect 132470 689570 132560 689810
rect 132800 689570 132910 689810
rect 133150 689570 133170 689810
rect 122170 689480 133170 689570
rect 122170 689240 122190 689480
rect 122430 689240 122520 689480
rect 122760 689240 122850 689480
rect 123090 689240 123180 689480
rect 123420 689240 123530 689480
rect 123770 689240 123860 689480
rect 124100 689240 124190 689480
rect 124430 689240 124520 689480
rect 124760 689240 124870 689480
rect 125110 689240 125200 689480
rect 125440 689240 125530 689480
rect 125770 689240 125860 689480
rect 126100 689240 126210 689480
rect 126450 689240 126540 689480
rect 126780 689240 126870 689480
rect 127110 689240 127200 689480
rect 127440 689240 127550 689480
rect 127790 689240 127880 689480
rect 128120 689240 128210 689480
rect 128450 689240 128540 689480
rect 128780 689240 128890 689480
rect 129130 689240 129220 689480
rect 129460 689240 129550 689480
rect 129790 689240 129880 689480
rect 130120 689240 130230 689480
rect 130470 689240 130560 689480
rect 130800 689240 130890 689480
rect 131130 689240 131220 689480
rect 131460 689240 131570 689480
rect 131810 689240 131900 689480
rect 132140 689240 132230 689480
rect 132470 689240 132560 689480
rect 132800 689240 132910 689480
rect 133150 689240 133170 689480
rect 122170 689130 133170 689240
rect 122170 688890 122190 689130
rect 122430 688890 122520 689130
rect 122760 688890 122850 689130
rect 123090 688890 123180 689130
rect 123420 688890 123530 689130
rect 123770 688890 123860 689130
rect 124100 688890 124190 689130
rect 124430 688890 124520 689130
rect 124760 688890 124870 689130
rect 125110 688890 125200 689130
rect 125440 688890 125530 689130
rect 125770 688890 125860 689130
rect 126100 688890 126210 689130
rect 126450 688890 126540 689130
rect 126780 688890 126870 689130
rect 127110 688890 127200 689130
rect 127440 688890 127550 689130
rect 127790 688890 127880 689130
rect 128120 688890 128210 689130
rect 128450 688890 128540 689130
rect 128780 688890 128890 689130
rect 129130 688890 129220 689130
rect 129460 688890 129550 689130
rect 129790 688890 129880 689130
rect 130120 688890 130230 689130
rect 130470 688890 130560 689130
rect 130800 688890 130890 689130
rect 131130 688890 131220 689130
rect 131460 688890 131570 689130
rect 131810 688890 131900 689130
rect 132140 688890 132230 689130
rect 132470 688890 132560 689130
rect 132800 688890 132910 689130
rect 133150 688890 133170 689130
rect 122170 688800 133170 688890
rect 122170 688560 122190 688800
rect 122430 688560 122520 688800
rect 122760 688560 122850 688800
rect 123090 688560 123180 688800
rect 123420 688560 123530 688800
rect 123770 688560 123860 688800
rect 124100 688560 124190 688800
rect 124430 688560 124520 688800
rect 124760 688560 124870 688800
rect 125110 688560 125200 688800
rect 125440 688560 125530 688800
rect 125770 688560 125860 688800
rect 126100 688560 126210 688800
rect 126450 688560 126540 688800
rect 126780 688560 126870 688800
rect 127110 688560 127200 688800
rect 127440 688560 127550 688800
rect 127790 688560 127880 688800
rect 128120 688560 128210 688800
rect 128450 688560 128540 688800
rect 128780 688560 128890 688800
rect 129130 688560 129220 688800
rect 129460 688560 129550 688800
rect 129790 688560 129880 688800
rect 130120 688560 130230 688800
rect 130470 688560 130560 688800
rect 130800 688560 130890 688800
rect 131130 688560 131220 688800
rect 131460 688560 131570 688800
rect 131810 688560 131900 688800
rect 132140 688560 132230 688800
rect 132470 688560 132560 688800
rect 132800 688560 132910 688800
rect 133150 688560 133170 688800
rect 122170 688470 133170 688560
rect 122170 688230 122190 688470
rect 122430 688230 122520 688470
rect 122760 688230 122850 688470
rect 123090 688230 123180 688470
rect 123420 688230 123530 688470
rect 123770 688230 123860 688470
rect 124100 688230 124190 688470
rect 124430 688230 124520 688470
rect 124760 688230 124870 688470
rect 125110 688230 125200 688470
rect 125440 688230 125530 688470
rect 125770 688230 125860 688470
rect 126100 688230 126210 688470
rect 126450 688230 126540 688470
rect 126780 688230 126870 688470
rect 127110 688230 127200 688470
rect 127440 688230 127550 688470
rect 127790 688230 127880 688470
rect 128120 688230 128210 688470
rect 128450 688230 128540 688470
rect 128780 688230 128890 688470
rect 129130 688230 129220 688470
rect 129460 688230 129550 688470
rect 129790 688230 129880 688470
rect 130120 688230 130230 688470
rect 130470 688230 130560 688470
rect 130800 688230 130890 688470
rect 131130 688230 131220 688470
rect 131460 688230 131570 688470
rect 131810 688230 131900 688470
rect 132140 688230 132230 688470
rect 132470 688230 132560 688470
rect 132800 688230 132910 688470
rect 133150 688230 133170 688470
rect 122170 688140 133170 688230
rect 122170 687900 122190 688140
rect 122430 687900 122520 688140
rect 122760 687900 122850 688140
rect 123090 687900 123180 688140
rect 123420 687900 123530 688140
rect 123770 687900 123860 688140
rect 124100 687900 124190 688140
rect 124430 687900 124520 688140
rect 124760 687900 124870 688140
rect 125110 687900 125200 688140
rect 125440 687900 125530 688140
rect 125770 687900 125860 688140
rect 126100 687900 126210 688140
rect 126450 687900 126540 688140
rect 126780 687900 126870 688140
rect 127110 687900 127200 688140
rect 127440 687900 127550 688140
rect 127790 687900 127880 688140
rect 128120 687900 128210 688140
rect 128450 687900 128540 688140
rect 128780 687900 128890 688140
rect 129130 687900 129220 688140
rect 129460 687900 129550 688140
rect 129790 687900 129880 688140
rect 130120 687900 130230 688140
rect 130470 687900 130560 688140
rect 130800 687900 130890 688140
rect 131130 687900 131220 688140
rect 131460 687900 131570 688140
rect 131810 687900 131900 688140
rect 132140 687900 132230 688140
rect 132470 687900 132560 688140
rect 132800 687900 132910 688140
rect 133150 687900 133170 688140
rect 122170 687790 133170 687900
rect 122170 687550 122190 687790
rect 122430 687550 122520 687790
rect 122760 687550 122850 687790
rect 123090 687550 123180 687790
rect 123420 687550 123530 687790
rect 123770 687550 123860 687790
rect 124100 687550 124190 687790
rect 124430 687550 124520 687790
rect 124760 687550 124870 687790
rect 125110 687550 125200 687790
rect 125440 687550 125530 687790
rect 125770 687550 125860 687790
rect 126100 687550 126210 687790
rect 126450 687550 126540 687790
rect 126780 687550 126870 687790
rect 127110 687550 127200 687790
rect 127440 687550 127550 687790
rect 127790 687550 127880 687790
rect 128120 687550 128210 687790
rect 128450 687550 128540 687790
rect 128780 687550 128890 687790
rect 129130 687550 129220 687790
rect 129460 687550 129550 687790
rect 129790 687550 129880 687790
rect 130120 687550 130230 687790
rect 130470 687550 130560 687790
rect 130800 687550 130890 687790
rect 131130 687550 131220 687790
rect 131460 687550 131570 687790
rect 131810 687550 131900 687790
rect 132140 687550 132230 687790
rect 132470 687550 132560 687790
rect 132800 687550 132910 687790
rect 133150 687550 133170 687790
rect 122170 687460 133170 687550
rect 122170 687220 122190 687460
rect 122430 687220 122520 687460
rect 122760 687220 122850 687460
rect 123090 687220 123180 687460
rect 123420 687220 123530 687460
rect 123770 687220 123860 687460
rect 124100 687220 124190 687460
rect 124430 687220 124520 687460
rect 124760 687220 124870 687460
rect 125110 687220 125200 687460
rect 125440 687220 125530 687460
rect 125770 687220 125860 687460
rect 126100 687220 126210 687460
rect 126450 687220 126540 687460
rect 126780 687220 126870 687460
rect 127110 687220 127200 687460
rect 127440 687220 127550 687460
rect 127790 687220 127880 687460
rect 128120 687220 128210 687460
rect 128450 687220 128540 687460
rect 128780 687220 128890 687460
rect 129130 687220 129220 687460
rect 129460 687220 129550 687460
rect 129790 687220 129880 687460
rect 130120 687220 130230 687460
rect 130470 687220 130560 687460
rect 130800 687220 130890 687460
rect 131130 687220 131220 687460
rect 131460 687220 131570 687460
rect 131810 687220 131900 687460
rect 132140 687220 132230 687460
rect 132470 687220 132560 687460
rect 132800 687220 132910 687460
rect 133150 687220 133170 687460
rect 122170 687130 133170 687220
rect 122170 686890 122190 687130
rect 122430 686890 122520 687130
rect 122760 686890 122850 687130
rect 123090 686890 123180 687130
rect 123420 686890 123530 687130
rect 123770 686890 123860 687130
rect 124100 686890 124190 687130
rect 124430 686890 124520 687130
rect 124760 686890 124870 687130
rect 125110 686890 125200 687130
rect 125440 686890 125530 687130
rect 125770 686890 125860 687130
rect 126100 686890 126210 687130
rect 126450 686890 126540 687130
rect 126780 686890 126870 687130
rect 127110 686890 127200 687130
rect 127440 686890 127550 687130
rect 127790 686890 127880 687130
rect 128120 686890 128210 687130
rect 128450 686890 128540 687130
rect 128780 686890 128890 687130
rect 129130 686890 129220 687130
rect 129460 686890 129550 687130
rect 129790 686890 129880 687130
rect 130120 686890 130230 687130
rect 130470 686890 130560 687130
rect 130800 686890 130890 687130
rect 131130 686890 131220 687130
rect 131460 686890 131570 687130
rect 131810 686890 131900 687130
rect 132140 686890 132230 687130
rect 132470 686890 132560 687130
rect 132800 686890 132910 687130
rect 133150 686890 133170 687130
rect 122170 686800 133170 686890
rect 122170 686560 122190 686800
rect 122430 686560 122520 686800
rect 122760 686560 122850 686800
rect 123090 686560 123180 686800
rect 123420 686560 123530 686800
rect 123770 686560 123860 686800
rect 124100 686560 124190 686800
rect 124430 686560 124520 686800
rect 124760 686560 124870 686800
rect 125110 686560 125200 686800
rect 125440 686560 125530 686800
rect 125770 686560 125860 686800
rect 126100 686560 126210 686800
rect 126450 686560 126540 686800
rect 126780 686560 126870 686800
rect 127110 686560 127200 686800
rect 127440 686560 127550 686800
rect 127790 686560 127880 686800
rect 128120 686560 128210 686800
rect 128450 686560 128540 686800
rect 128780 686560 128890 686800
rect 129130 686560 129220 686800
rect 129460 686560 129550 686800
rect 129790 686560 129880 686800
rect 130120 686560 130230 686800
rect 130470 686560 130560 686800
rect 130800 686560 130890 686800
rect 131130 686560 131220 686800
rect 131460 686560 131570 686800
rect 131810 686560 131900 686800
rect 132140 686560 132230 686800
rect 132470 686560 132560 686800
rect 132800 686560 132910 686800
rect 133150 686560 133170 686800
rect 122170 686450 133170 686560
rect 122170 686210 122190 686450
rect 122430 686210 122520 686450
rect 122760 686210 122850 686450
rect 123090 686210 123180 686450
rect 123420 686210 123530 686450
rect 123770 686210 123860 686450
rect 124100 686210 124190 686450
rect 124430 686210 124520 686450
rect 124760 686210 124870 686450
rect 125110 686210 125200 686450
rect 125440 686210 125530 686450
rect 125770 686210 125860 686450
rect 126100 686210 126210 686450
rect 126450 686210 126540 686450
rect 126780 686210 126870 686450
rect 127110 686210 127200 686450
rect 127440 686210 127550 686450
rect 127790 686210 127880 686450
rect 128120 686210 128210 686450
rect 128450 686210 128540 686450
rect 128780 686210 128890 686450
rect 129130 686210 129220 686450
rect 129460 686210 129550 686450
rect 129790 686210 129880 686450
rect 130120 686210 130230 686450
rect 130470 686210 130560 686450
rect 130800 686210 130890 686450
rect 131130 686210 131220 686450
rect 131460 686210 131570 686450
rect 131810 686210 131900 686450
rect 132140 686210 132230 686450
rect 132470 686210 132560 686450
rect 132800 686210 132910 686450
rect 133150 686210 133170 686450
rect 122170 686120 133170 686210
rect 122170 685880 122190 686120
rect 122430 685880 122520 686120
rect 122760 685880 122850 686120
rect 123090 685880 123180 686120
rect 123420 685880 123530 686120
rect 123770 685880 123860 686120
rect 124100 685880 124190 686120
rect 124430 685880 124520 686120
rect 124760 685880 124870 686120
rect 125110 685880 125200 686120
rect 125440 685880 125530 686120
rect 125770 685880 125860 686120
rect 126100 685880 126210 686120
rect 126450 685880 126540 686120
rect 126780 685880 126870 686120
rect 127110 685880 127200 686120
rect 127440 685880 127550 686120
rect 127790 685880 127880 686120
rect 128120 685880 128210 686120
rect 128450 685880 128540 686120
rect 128780 685880 128890 686120
rect 129130 685880 129220 686120
rect 129460 685880 129550 686120
rect 129790 685880 129880 686120
rect 130120 685880 130230 686120
rect 130470 685880 130560 686120
rect 130800 685880 130890 686120
rect 131130 685880 131220 686120
rect 131460 685880 131570 686120
rect 131810 685880 131900 686120
rect 132140 685880 132230 686120
rect 132470 685880 132560 686120
rect 132800 685880 132910 686120
rect 133150 685880 133170 686120
rect 122170 685790 133170 685880
rect 122170 685550 122190 685790
rect 122430 685550 122520 685790
rect 122760 685550 122850 685790
rect 123090 685550 123180 685790
rect 123420 685550 123530 685790
rect 123770 685550 123860 685790
rect 124100 685550 124190 685790
rect 124430 685550 124520 685790
rect 124760 685550 124870 685790
rect 125110 685550 125200 685790
rect 125440 685550 125530 685790
rect 125770 685550 125860 685790
rect 126100 685550 126210 685790
rect 126450 685550 126540 685790
rect 126780 685550 126870 685790
rect 127110 685550 127200 685790
rect 127440 685550 127550 685790
rect 127790 685550 127880 685790
rect 128120 685550 128210 685790
rect 128450 685550 128540 685790
rect 128780 685550 128890 685790
rect 129130 685550 129220 685790
rect 129460 685550 129550 685790
rect 129790 685550 129880 685790
rect 130120 685550 130230 685790
rect 130470 685550 130560 685790
rect 130800 685550 130890 685790
rect 131130 685550 131220 685790
rect 131460 685550 131570 685790
rect 131810 685550 131900 685790
rect 132140 685550 132230 685790
rect 132470 685550 132560 685790
rect 132800 685550 132910 685790
rect 133150 685550 133170 685790
rect 122170 685460 133170 685550
rect 122170 685220 122190 685460
rect 122430 685220 122520 685460
rect 122760 685220 122850 685460
rect 123090 685220 123180 685460
rect 123420 685220 123530 685460
rect 123770 685220 123860 685460
rect 124100 685220 124190 685460
rect 124430 685220 124520 685460
rect 124760 685220 124870 685460
rect 125110 685220 125200 685460
rect 125440 685220 125530 685460
rect 125770 685220 125860 685460
rect 126100 685220 126210 685460
rect 126450 685220 126540 685460
rect 126780 685220 126870 685460
rect 127110 685220 127200 685460
rect 127440 685220 127550 685460
rect 127790 685220 127880 685460
rect 128120 685220 128210 685460
rect 128450 685220 128540 685460
rect 128780 685220 128890 685460
rect 129130 685220 129220 685460
rect 129460 685220 129550 685460
rect 129790 685220 129880 685460
rect 130120 685220 130230 685460
rect 130470 685220 130560 685460
rect 130800 685220 130890 685460
rect 131130 685220 131220 685460
rect 131460 685220 131570 685460
rect 131810 685220 131900 685460
rect 132140 685220 132230 685460
rect 132470 685220 132560 685460
rect 132800 685220 132910 685460
rect 133150 685220 133170 685460
rect 122170 685110 133170 685220
rect 122170 684870 122190 685110
rect 122430 684870 122520 685110
rect 122760 684870 122850 685110
rect 123090 684870 123180 685110
rect 123420 684870 123530 685110
rect 123770 684870 123860 685110
rect 124100 684870 124190 685110
rect 124430 684870 124520 685110
rect 124760 684870 124870 685110
rect 125110 684870 125200 685110
rect 125440 684870 125530 685110
rect 125770 684870 125860 685110
rect 126100 684870 126210 685110
rect 126450 684870 126540 685110
rect 126780 684870 126870 685110
rect 127110 684870 127200 685110
rect 127440 684870 127550 685110
rect 127790 684870 127880 685110
rect 128120 684870 128210 685110
rect 128450 684870 128540 685110
rect 128780 684870 128890 685110
rect 129130 684870 129220 685110
rect 129460 684870 129550 685110
rect 129790 684870 129880 685110
rect 130120 684870 130230 685110
rect 130470 684870 130560 685110
rect 130800 684870 130890 685110
rect 131130 684870 131220 685110
rect 131460 684870 131570 685110
rect 131810 684870 131900 685110
rect 132140 684870 132230 685110
rect 132470 684870 132560 685110
rect 132800 684870 132910 685110
rect 133150 684870 133170 685110
rect 122170 684780 133170 684870
rect 122170 684540 122190 684780
rect 122430 684540 122520 684780
rect 122760 684540 122850 684780
rect 123090 684540 123180 684780
rect 123420 684540 123530 684780
rect 123770 684540 123860 684780
rect 124100 684540 124190 684780
rect 124430 684540 124520 684780
rect 124760 684540 124870 684780
rect 125110 684540 125200 684780
rect 125440 684540 125530 684780
rect 125770 684540 125860 684780
rect 126100 684540 126210 684780
rect 126450 684540 126540 684780
rect 126780 684540 126870 684780
rect 127110 684540 127200 684780
rect 127440 684540 127550 684780
rect 127790 684540 127880 684780
rect 128120 684540 128210 684780
rect 128450 684540 128540 684780
rect 128780 684540 128890 684780
rect 129130 684540 129220 684780
rect 129460 684540 129550 684780
rect 129790 684540 129880 684780
rect 130120 684540 130230 684780
rect 130470 684540 130560 684780
rect 130800 684540 130890 684780
rect 131130 684540 131220 684780
rect 131460 684540 131570 684780
rect 131810 684540 131900 684780
rect 132140 684540 132230 684780
rect 132470 684540 132560 684780
rect 132800 684540 132910 684780
rect 133150 684540 133170 684780
rect 122170 684450 133170 684540
rect 122170 684210 122190 684450
rect 122430 684210 122520 684450
rect 122760 684210 122850 684450
rect 123090 684210 123180 684450
rect 123420 684210 123530 684450
rect 123770 684210 123860 684450
rect 124100 684210 124190 684450
rect 124430 684210 124520 684450
rect 124760 684210 124870 684450
rect 125110 684210 125200 684450
rect 125440 684210 125530 684450
rect 125770 684210 125860 684450
rect 126100 684210 126210 684450
rect 126450 684210 126540 684450
rect 126780 684210 126870 684450
rect 127110 684210 127200 684450
rect 127440 684210 127550 684450
rect 127790 684210 127880 684450
rect 128120 684210 128210 684450
rect 128450 684210 128540 684450
rect 128780 684210 128890 684450
rect 129130 684210 129220 684450
rect 129460 684210 129550 684450
rect 129790 684210 129880 684450
rect 130120 684210 130230 684450
rect 130470 684210 130560 684450
rect 130800 684210 130890 684450
rect 131130 684210 131220 684450
rect 131460 684210 131570 684450
rect 131810 684210 131900 684450
rect 132140 684210 132230 684450
rect 132470 684210 132560 684450
rect 132800 684210 132910 684450
rect 133150 684210 133170 684450
rect 122170 684120 133170 684210
rect 122170 683880 122190 684120
rect 122430 683880 122520 684120
rect 122760 683880 122850 684120
rect 123090 683880 123180 684120
rect 123420 683880 123530 684120
rect 123770 683880 123860 684120
rect 124100 683880 124190 684120
rect 124430 683880 124520 684120
rect 124760 683880 124870 684120
rect 125110 683880 125200 684120
rect 125440 683880 125530 684120
rect 125770 683880 125860 684120
rect 126100 683880 126210 684120
rect 126450 683880 126540 684120
rect 126780 683880 126870 684120
rect 127110 683880 127200 684120
rect 127440 683880 127550 684120
rect 127790 683880 127880 684120
rect 128120 683880 128210 684120
rect 128450 683880 128540 684120
rect 128780 683880 128890 684120
rect 129130 683880 129220 684120
rect 129460 683880 129550 684120
rect 129790 683880 129880 684120
rect 130120 683880 130230 684120
rect 130470 683880 130560 684120
rect 130800 683880 130890 684120
rect 131130 683880 131220 684120
rect 131460 683880 131570 684120
rect 131810 683880 131900 684120
rect 132140 683880 132230 684120
rect 132470 683880 132560 684120
rect 132800 683880 132910 684120
rect 133150 683880 133170 684120
rect 122170 683860 133170 683880
rect 133550 694840 144550 694860
rect 133550 694600 133570 694840
rect 133810 694600 133900 694840
rect 134140 694600 134230 694840
rect 134470 694600 134560 694840
rect 134800 694600 134910 694840
rect 135150 694600 135240 694840
rect 135480 694600 135570 694840
rect 135810 694600 135900 694840
rect 136140 694600 136250 694840
rect 136490 694600 136580 694840
rect 136820 694600 136910 694840
rect 137150 694600 137240 694840
rect 137480 694600 137590 694840
rect 137830 694600 137920 694840
rect 138160 694600 138250 694840
rect 138490 694600 138580 694840
rect 138820 694600 138930 694840
rect 139170 694600 139260 694840
rect 139500 694600 139590 694840
rect 139830 694600 139920 694840
rect 140160 694600 140270 694840
rect 140510 694600 140600 694840
rect 140840 694600 140930 694840
rect 141170 694600 141260 694840
rect 141500 694600 141610 694840
rect 141850 694600 141940 694840
rect 142180 694600 142270 694840
rect 142510 694600 142600 694840
rect 142840 694600 142950 694840
rect 143190 694600 143280 694840
rect 143520 694600 143610 694840
rect 143850 694600 143940 694840
rect 144180 694600 144290 694840
rect 144530 694600 144550 694840
rect 133550 694490 144550 694600
rect 133550 694250 133570 694490
rect 133810 694250 133900 694490
rect 134140 694250 134230 694490
rect 134470 694250 134560 694490
rect 134800 694250 134910 694490
rect 135150 694250 135240 694490
rect 135480 694250 135570 694490
rect 135810 694250 135900 694490
rect 136140 694250 136250 694490
rect 136490 694250 136580 694490
rect 136820 694250 136910 694490
rect 137150 694250 137240 694490
rect 137480 694250 137590 694490
rect 137830 694250 137920 694490
rect 138160 694250 138250 694490
rect 138490 694250 138580 694490
rect 138820 694250 138930 694490
rect 139170 694250 139260 694490
rect 139500 694250 139590 694490
rect 139830 694250 139920 694490
rect 140160 694250 140270 694490
rect 140510 694250 140600 694490
rect 140840 694250 140930 694490
rect 141170 694250 141260 694490
rect 141500 694250 141610 694490
rect 141850 694250 141940 694490
rect 142180 694250 142270 694490
rect 142510 694250 142600 694490
rect 142840 694250 142950 694490
rect 143190 694250 143280 694490
rect 143520 694250 143610 694490
rect 143850 694250 143940 694490
rect 144180 694250 144290 694490
rect 144530 694250 144550 694490
rect 133550 694160 144550 694250
rect 133550 693920 133570 694160
rect 133810 693920 133900 694160
rect 134140 693920 134230 694160
rect 134470 693920 134560 694160
rect 134800 693920 134910 694160
rect 135150 693920 135240 694160
rect 135480 693920 135570 694160
rect 135810 693920 135900 694160
rect 136140 693920 136250 694160
rect 136490 693920 136580 694160
rect 136820 693920 136910 694160
rect 137150 693920 137240 694160
rect 137480 693920 137590 694160
rect 137830 693920 137920 694160
rect 138160 693920 138250 694160
rect 138490 693920 138580 694160
rect 138820 693920 138930 694160
rect 139170 693920 139260 694160
rect 139500 693920 139590 694160
rect 139830 693920 139920 694160
rect 140160 693920 140270 694160
rect 140510 693920 140600 694160
rect 140840 693920 140930 694160
rect 141170 693920 141260 694160
rect 141500 693920 141610 694160
rect 141850 693920 141940 694160
rect 142180 693920 142270 694160
rect 142510 693920 142600 694160
rect 142840 693920 142950 694160
rect 143190 693920 143280 694160
rect 143520 693920 143610 694160
rect 143850 693920 143940 694160
rect 144180 693920 144290 694160
rect 144530 693920 144550 694160
rect 133550 693830 144550 693920
rect 133550 693590 133570 693830
rect 133810 693590 133900 693830
rect 134140 693590 134230 693830
rect 134470 693590 134560 693830
rect 134800 693590 134910 693830
rect 135150 693590 135240 693830
rect 135480 693590 135570 693830
rect 135810 693590 135900 693830
rect 136140 693590 136250 693830
rect 136490 693590 136580 693830
rect 136820 693590 136910 693830
rect 137150 693590 137240 693830
rect 137480 693590 137590 693830
rect 137830 693590 137920 693830
rect 138160 693590 138250 693830
rect 138490 693590 138580 693830
rect 138820 693590 138930 693830
rect 139170 693590 139260 693830
rect 139500 693590 139590 693830
rect 139830 693590 139920 693830
rect 140160 693590 140270 693830
rect 140510 693590 140600 693830
rect 140840 693590 140930 693830
rect 141170 693590 141260 693830
rect 141500 693590 141610 693830
rect 141850 693590 141940 693830
rect 142180 693590 142270 693830
rect 142510 693590 142600 693830
rect 142840 693590 142950 693830
rect 143190 693590 143280 693830
rect 143520 693590 143610 693830
rect 143850 693590 143940 693830
rect 144180 693590 144290 693830
rect 144530 693590 144550 693830
rect 133550 693500 144550 693590
rect 133550 693260 133570 693500
rect 133810 693260 133900 693500
rect 134140 693260 134230 693500
rect 134470 693260 134560 693500
rect 134800 693260 134910 693500
rect 135150 693260 135240 693500
rect 135480 693260 135570 693500
rect 135810 693260 135900 693500
rect 136140 693260 136250 693500
rect 136490 693260 136580 693500
rect 136820 693260 136910 693500
rect 137150 693260 137240 693500
rect 137480 693260 137590 693500
rect 137830 693260 137920 693500
rect 138160 693260 138250 693500
rect 138490 693260 138580 693500
rect 138820 693260 138930 693500
rect 139170 693260 139260 693500
rect 139500 693260 139590 693500
rect 139830 693260 139920 693500
rect 140160 693260 140270 693500
rect 140510 693260 140600 693500
rect 140840 693260 140930 693500
rect 141170 693260 141260 693500
rect 141500 693260 141610 693500
rect 141850 693260 141940 693500
rect 142180 693260 142270 693500
rect 142510 693260 142600 693500
rect 142840 693260 142950 693500
rect 143190 693260 143280 693500
rect 143520 693260 143610 693500
rect 143850 693260 143940 693500
rect 144180 693260 144290 693500
rect 144530 693260 144550 693500
rect 133550 693150 144550 693260
rect 133550 692910 133570 693150
rect 133810 692910 133900 693150
rect 134140 692910 134230 693150
rect 134470 692910 134560 693150
rect 134800 692910 134910 693150
rect 135150 692910 135240 693150
rect 135480 692910 135570 693150
rect 135810 692910 135900 693150
rect 136140 692910 136250 693150
rect 136490 692910 136580 693150
rect 136820 692910 136910 693150
rect 137150 692910 137240 693150
rect 137480 692910 137590 693150
rect 137830 692910 137920 693150
rect 138160 692910 138250 693150
rect 138490 692910 138580 693150
rect 138820 692910 138930 693150
rect 139170 692910 139260 693150
rect 139500 692910 139590 693150
rect 139830 692910 139920 693150
rect 140160 692910 140270 693150
rect 140510 692910 140600 693150
rect 140840 692910 140930 693150
rect 141170 692910 141260 693150
rect 141500 692910 141610 693150
rect 141850 692910 141940 693150
rect 142180 692910 142270 693150
rect 142510 692910 142600 693150
rect 142840 692910 142950 693150
rect 143190 692910 143280 693150
rect 143520 692910 143610 693150
rect 143850 692910 143940 693150
rect 144180 692910 144290 693150
rect 144530 692910 144550 693150
rect 133550 692820 144550 692910
rect 133550 692580 133570 692820
rect 133810 692580 133900 692820
rect 134140 692580 134230 692820
rect 134470 692580 134560 692820
rect 134800 692580 134910 692820
rect 135150 692580 135240 692820
rect 135480 692580 135570 692820
rect 135810 692580 135900 692820
rect 136140 692580 136250 692820
rect 136490 692580 136580 692820
rect 136820 692580 136910 692820
rect 137150 692580 137240 692820
rect 137480 692580 137590 692820
rect 137830 692580 137920 692820
rect 138160 692580 138250 692820
rect 138490 692580 138580 692820
rect 138820 692580 138930 692820
rect 139170 692580 139260 692820
rect 139500 692580 139590 692820
rect 139830 692580 139920 692820
rect 140160 692580 140270 692820
rect 140510 692580 140600 692820
rect 140840 692580 140930 692820
rect 141170 692580 141260 692820
rect 141500 692580 141610 692820
rect 141850 692580 141940 692820
rect 142180 692580 142270 692820
rect 142510 692580 142600 692820
rect 142840 692580 142950 692820
rect 143190 692580 143280 692820
rect 143520 692580 143610 692820
rect 143850 692580 143940 692820
rect 144180 692580 144290 692820
rect 144530 692580 144550 692820
rect 133550 692490 144550 692580
rect 133550 692250 133570 692490
rect 133810 692250 133900 692490
rect 134140 692250 134230 692490
rect 134470 692250 134560 692490
rect 134800 692250 134910 692490
rect 135150 692250 135240 692490
rect 135480 692250 135570 692490
rect 135810 692250 135900 692490
rect 136140 692250 136250 692490
rect 136490 692250 136580 692490
rect 136820 692250 136910 692490
rect 137150 692250 137240 692490
rect 137480 692250 137590 692490
rect 137830 692250 137920 692490
rect 138160 692250 138250 692490
rect 138490 692250 138580 692490
rect 138820 692250 138930 692490
rect 139170 692250 139260 692490
rect 139500 692250 139590 692490
rect 139830 692250 139920 692490
rect 140160 692250 140270 692490
rect 140510 692250 140600 692490
rect 140840 692250 140930 692490
rect 141170 692250 141260 692490
rect 141500 692250 141610 692490
rect 141850 692250 141940 692490
rect 142180 692250 142270 692490
rect 142510 692250 142600 692490
rect 142840 692250 142950 692490
rect 143190 692250 143280 692490
rect 143520 692250 143610 692490
rect 143850 692250 143940 692490
rect 144180 692250 144290 692490
rect 144530 692250 144550 692490
rect 133550 692160 144550 692250
rect 133550 691920 133570 692160
rect 133810 691920 133900 692160
rect 134140 691920 134230 692160
rect 134470 691920 134560 692160
rect 134800 691920 134910 692160
rect 135150 691920 135240 692160
rect 135480 691920 135570 692160
rect 135810 691920 135900 692160
rect 136140 691920 136250 692160
rect 136490 691920 136580 692160
rect 136820 691920 136910 692160
rect 137150 691920 137240 692160
rect 137480 691920 137590 692160
rect 137830 691920 137920 692160
rect 138160 691920 138250 692160
rect 138490 691920 138580 692160
rect 138820 691920 138930 692160
rect 139170 691920 139260 692160
rect 139500 691920 139590 692160
rect 139830 691920 139920 692160
rect 140160 691920 140270 692160
rect 140510 691920 140600 692160
rect 140840 691920 140930 692160
rect 141170 691920 141260 692160
rect 141500 691920 141610 692160
rect 141850 691920 141940 692160
rect 142180 691920 142270 692160
rect 142510 691920 142600 692160
rect 142840 691920 142950 692160
rect 143190 691920 143280 692160
rect 143520 691920 143610 692160
rect 143850 691920 143940 692160
rect 144180 691920 144290 692160
rect 144530 691920 144550 692160
rect 133550 691810 144550 691920
rect 133550 691570 133570 691810
rect 133810 691570 133900 691810
rect 134140 691570 134230 691810
rect 134470 691570 134560 691810
rect 134800 691570 134910 691810
rect 135150 691570 135240 691810
rect 135480 691570 135570 691810
rect 135810 691570 135900 691810
rect 136140 691570 136250 691810
rect 136490 691570 136580 691810
rect 136820 691570 136910 691810
rect 137150 691570 137240 691810
rect 137480 691570 137590 691810
rect 137830 691570 137920 691810
rect 138160 691570 138250 691810
rect 138490 691570 138580 691810
rect 138820 691570 138930 691810
rect 139170 691570 139260 691810
rect 139500 691570 139590 691810
rect 139830 691570 139920 691810
rect 140160 691570 140270 691810
rect 140510 691570 140600 691810
rect 140840 691570 140930 691810
rect 141170 691570 141260 691810
rect 141500 691570 141610 691810
rect 141850 691570 141940 691810
rect 142180 691570 142270 691810
rect 142510 691570 142600 691810
rect 142840 691570 142950 691810
rect 143190 691570 143280 691810
rect 143520 691570 143610 691810
rect 143850 691570 143940 691810
rect 144180 691570 144290 691810
rect 144530 691570 144550 691810
rect 133550 691480 144550 691570
rect 133550 691240 133570 691480
rect 133810 691240 133900 691480
rect 134140 691240 134230 691480
rect 134470 691240 134560 691480
rect 134800 691240 134910 691480
rect 135150 691240 135240 691480
rect 135480 691240 135570 691480
rect 135810 691240 135900 691480
rect 136140 691240 136250 691480
rect 136490 691240 136580 691480
rect 136820 691240 136910 691480
rect 137150 691240 137240 691480
rect 137480 691240 137590 691480
rect 137830 691240 137920 691480
rect 138160 691240 138250 691480
rect 138490 691240 138580 691480
rect 138820 691240 138930 691480
rect 139170 691240 139260 691480
rect 139500 691240 139590 691480
rect 139830 691240 139920 691480
rect 140160 691240 140270 691480
rect 140510 691240 140600 691480
rect 140840 691240 140930 691480
rect 141170 691240 141260 691480
rect 141500 691240 141610 691480
rect 141850 691240 141940 691480
rect 142180 691240 142270 691480
rect 142510 691240 142600 691480
rect 142840 691240 142950 691480
rect 143190 691240 143280 691480
rect 143520 691240 143610 691480
rect 143850 691240 143940 691480
rect 144180 691240 144290 691480
rect 144530 691240 144550 691480
rect 133550 691150 144550 691240
rect 133550 690910 133570 691150
rect 133810 690910 133900 691150
rect 134140 690910 134230 691150
rect 134470 690910 134560 691150
rect 134800 690910 134910 691150
rect 135150 690910 135240 691150
rect 135480 690910 135570 691150
rect 135810 690910 135900 691150
rect 136140 690910 136250 691150
rect 136490 690910 136580 691150
rect 136820 690910 136910 691150
rect 137150 690910 137240 691150
rect 137480 690910 137590 691150
rect 137830 690910 137920 691150
rect 138160 690910 138250 691150
rect 138490 690910 138580 691150
rect 138820 690910 138930 691150
rect 139170 690910 139260 691150
rect 139500 690910 139590 691150
rect 139830 690910 139920 691150
rect 140160 690910 140270 691150
rect 140510 690910 140600 691150
rect 140840 690910 140930 691150
rect 141170 690910 141260 691150
rect 141500 690910 141610 691150
rect 141850 690910 141940 691150
rect 142180 690910 142270 691150
rect 142510 690910 142600 691150
rect 142840 690910 142950 691150
rect 143190 690910 143280 691150
rect 143520 690910 143610 691150
rect 143850 690910 143940 691150
rect 144180 690910 144290 691150
rect 144530 690910 144550 691150
rect 133550 690820 144550 690910
rect 133550 690580 133570 690820
rect 133810 690580 133900 690820
rect 134140 690580 134230 690820
rect 134470 690580 134560 690820
rect 134800 690580 134910 690820
rect 135150 690580 135240 690820
rect 135480 690580 135570 690820
rect 135810 690580 135900 690820
rect 136140 690580 136250 690820
rect 136490 690580 136580 690820
rect 136820 690580 136910 690820
rect 137150 690580 137240 690820
rect 137480 690580 137590 690820
rect 137830 690580 137920 690820
rect 138160 690580 138250 690820
rect 138490 690580 138580 690820
rect 138820 690580 138930 690820
rect 139170 690580 139260 690820
rect 139500 690580 139590 690820
rect 139830 690580 139920 690820
rect 140160 690580 140270 690820
rect 140510 690580 140600 690820
rect 140840 690580 140930 690820
rect 141170 690580 141260 690820
rect 141500 690580 141610 690820
rect 141850 690580 141940 690820
rect 142180 690580 142270 690820
rect 142510 690580 142600 690820
rect 142840 690580 142950 690820
rect 143190 690580 143280 690820
rect 143520 690580 143610 690820
rect 143850 690580 143940 690820
rect 144180 690580 144290 690820
rect 144530 690580 144550 690820
rect 133550 690470 144550 690580
rect 133550 690230 133570 690470
rect 133810 690230 133900 690470
rect 134140 690230 134230 690470
rect 134470 690230 134560 690470
rect 134800 690230 134910 690470
rect 135150 690230 135240 690470
rect 135480 690230 135570 690470
rect 135810 690230 135900 690470
rect 136140 690230 136250 690470
rect 136490 690230 136580 690470
rect 136820 690230 136910 690470
rect 137150 690230 137240 690470
rect 137480 690230 137590 690470
rect 137830 690230 137920 690470
rect 138160 690230 138250 690470
rect 138490 690230 138580 690470
rect 138820 690230 138930 690470
rect 139170 690230 139260 690470
rect 139500 690230 139590 690470
rect 139830 690230 139920 690470
rect 140160 690230 140270 690470
rect 140510 690230 140600 690470
rect 140840 690230 140930 690470
rect 141170 690230 141260 690470
rect 141500 690230 141610 690470
rect 141850 690230 141940 690470
rect 142180 690230 142270 690470
rect 142510 690230 142600 690470
rect 142840 690230 142950 690470
rect 143190 690230 143280 690470
rect 143520 690230 143610 690470
rect 143850 690230 143940 690470
rect 144180 690230 144290 690470
rect 144530 690230 144550 690470
rect 133550 690140 144550 690230
rect 133550 689900 133570 690140
rect 133810 689900 133900 690140
rect 134140 689900 134230 690140
rect 134470 689900 134560 690140
rect 134800 689900 134910 690140
rect 135150 689900 135240 690140
rect 135480 689900 135570 690140
rect 135810 689900 135900 690140
rect 136140 689900 136250 690140
rect 136490 689900 136580 690140
rect 136820 689900 136910 690140
rect 137150 689900 137240 690140
rect 137480 689900 137590 690140
rect 137830 689900 137920 690140
rect 138160 689900 138250 690140
rect 138490 689900 138580 690140
rect 138820 689900 138930 690140
rect 139170 689900 139260 690140
rect 139500 689900 139590 690140
rect 139830 689900 139920 690140
rect 140160 689900 140270 690140
rect 140510 689900 140600 690140
rect 140840 689900 140930 690140
rect 141170 689900 141260 690140
rect 141500 689900 141610 690140
rect 141850 689900 141940 690140
rect 142180 689900 142270 690140
rect 142510 689900 142600 690140
rect 142840 689900 142950 690140
rect 143190 689900 143280 690140
rect 143520 689900 143610 690140
rect 143850 689900 143940 690140
rect 144180 689900 144290 690140
rect 144530 689900 144550 690140
rect 133550 689810 144550 689900
rect 133550 689570 133570 689810
rect 133810 689570 133900 689810
rect 134140 689570 134230 689810
rect 134470 689570 134560 689810
rect 134800 689570 134910 689810
rect 135150 689570 135240 689810
rect 135480 689570 135570 689810
rect 135810 689570 135900 689810
rect 136140 689570 136250 689810
rect 136490 689570 136580 689810
rect 136820 689570 136910 689810
rect 137150 689570 137240 689810
rect 137480 689570 137590 689810
rect 137830 689570 137920 689810
rect 138160 689570 138250 689810
rect 138490 689570 138580 689810
rect 138820 689570 138930 689810
rect 139170 689570 139260 689810
rect 139500 689570 139590 689810
rect 139830 689570 139920 689810
rect 140160 689570 140270 689810
rect 140510 689570 140600 689810
rect 140840 689570 140930 689810
rect 141170 689570 141260 689810
rect 141500 689570 141610 689810
rect 141850 689570 141940 689810
rect 142180 689570 142270 689810
rect 142510 689570 142600 689810
rect 142840 689570 142950 689810
rect 143190 689570 143280 689810
rect 143520 689570 143610 689810
rect 143850 689570 143940 689810
rect 144180 689570 144290 689810
rect 144530 689570 144550 689810
rect 133550 689480 144550 689570
rect 133550 689240 133570 689480
rect 133810 689240 133900 689480
rect 134140 689240 134230 689480
rect 134470 689240 134560 689480
rect 134800 689240 134910 689480
rect 135150 689240 135240 689480
rect 135480 689240 135570 689480
rect 135810 689240 135900 689480
rect 136140 689240 136250 689480
rect 136490 689240 136580 689480
rect 136820 689240 136910 689480
rect 137150 689240 137240 689480
rect 137480 689240 137590 689480
rect 137830 689240 137920 689480
rect 138160 689240 138250 689480
rect 138490 689240 138580 689480
rect 138820 689240 138930 689480
rect 139170 689240 139260 689480
rect 139500 689240 139590 689480
rect 139830 689240 139920 689480
rect 140160 689240 140270 689480
rect 140510 689240 140600 689480
rect 140840 689240 140930 689480
rect 141170 689240 141260 689480
rect 141500 689240 141610 689480
rect 141850 689240 141940 689480
rect 142180 689240 142270 689480
rect 142510 689240 142600 689480
rect 142840 689240 142950 689480
rect 143190 689240 143280 689480
rect 143520 689240 143610 689480
rect 143850 689240 143940 689480
rect 144180 689240 144290 689480
rect 144530 689240 144550 689480
rect 133550 689130 144550 689240
rect 133550 688890 133570 689130
rect 133810 688890 133900 689130
rect 134140 688890 134230 689130
rect 134470 688890 134560 689130
rect 134800 688890 134910 689130
rect 135150 688890 135240 689130
rect 135480 688890 135570 689130
rect 135810 688890 135900 689130
rect 136140 688890 136250 689130
rect 136490 688890 136580 689130
rect 136820 688890 136910 689130
rect 137150 688890 137240 689130
rect 137480 688890 137590 689130
rect 137830 688890 137920 689130
rect 138160 688890 138250 689130
rect 138490 688890 138580 689130
rect 138820 688890 138930 689130
rect 139170 688890 139260 689130
rect 139500 688890 139590 689130
rect 139830 688890 139920 689130
rect 140160 688890 140270 689130
rect 140510 688890 140600 689130
rect 140840 688890 140930 689130
rect 141170 688890 141260 689130
rect 141500 688890 141610 689130
rect 141850 688890 141940 689130
rect 142180 688890 142270 689130
rect 142510 688890 142600 689130
rect 142840 688890 142950 689130
rect 143190 688890 143280 689130
rect 143520 688890 143610 689130
rect 143850 688890 143940 689130
rect 144180 688890 144290 689130
rect 144530 688890 144550 689130
rect 133550 688800 144550 688890
rect 133550 688560 133570 688800
rect 133810 688560 133900 688800
rect 134140 688560 134230 688800
rect 134470 688560 134560 688800
rect 134800 688560 134910 688800
rect 135150 688560 135240 688800
rect 135480 688560 135570 688800
rect 135810 688560 135900 688800
rect 136140 688560 136250 688800
rect 136490 688560 136580 688800
rect 136820 688560 136910 688800
rect 137150 688560 137240 688800
rect 137480 688560 137590 688800
rect 137830 688560 137920 688800
rect 138160 688560 138250 688800
rect 138490 688560 138580 688800
rect 138820 688560 138930 688800
rect 139170 688560 139260 688800
rect 139500 688560 139590 688800
rect 139830 688560 139920 688800
rect 140160 688560 140270 688800
rect 140510 688560 140600 688800
rect 140840 688560 140930 688800
rect 141170 688560 141260 688800
rect 141500 688560 141610 688800
rect 141850 688560 141940 688800
rect 142180 688560 142270 688800
rect 142510 688560 142600 688800
rect 142840 688560 142950 688800
rect 143190 688560 143280 688800
rect 143520 688560 143610 688800
rect 143850 688560 143940 688800
rect 144180 688560 144290 688800
rect 144530 688560 144550 688800
rect 133550 688470 144550 688560
rect 133550 688230 133570 688470
rect 133810 688230 133900 688470
rect 134140 688230 134230 688470
rect 134470 688230 134560 688470
rect 134800 688230 134910 688470
rect 135150 688230 135240 688470
rect 135480 688230 135570 688470
rect 135810 688230 135900 688470
rect 136140 688230 136250 688470
rect 136490 688230 136580 688470
rect 136820 688230 136910 688470
rect 137150 688230 137240 688470
rect 137480 688230 137590 688470
rect 137830 688230 137920 688470
rect 138160 688230 138250 688470
rect 138490 688230 138580 688470
rect 138820 688230 138930 688470
rect 139170 688230 139260 688470
rect 139500 688230 139590 688470
rect 139830 688230 139920 688470
rect 140160 688230 140270 688470
rect 140510 688230 140600 688470
rect 140840 688230 140930 688470
rect 141170 688230 141260 688470
rect 141500 688230 141610 688470
rect 141850 688230 141940 688470
rect 142180 688230 142270 688470
rect 142510 688230 142600 688470
rect 142840 688230 142950 688470
rect 143190 688230 143280 688470
rect 143520 688230 143610 688470
rect 143850 688230 143940 688470
rect 144180 688230 144290 688470
rect 144530 688230 144550 688470
rect 133550 688140 144550 688230
rect 133550 687900 133570 688140
rect 133810 687900 133900 688140
rect 134140 687900 134230 688140
rect 134470 687900 134560 688140
rect 134800 687900 134910 688140
rect 135150 687900 135240 688140
rect 135480 687900 135570 688140
rect 135810 687900 135900 688140
rect 136140 687900 136250 688140
rect 136490 687900 136580 688140
rect 136820 687900 136910 688140
rect 137150 687900 137240 688140
rect 137480 687900 137590 688140
rect 137830 687900 137920 688140
rect 138160 687900 138250 688140
rect 138490 687900 138580 688140
rect 138820 687900 138930 688140
rect 139170 687900 139260 688140
rect 139500 687900 139590 688140
rect 139830 687900 139920 688140
rect 140160 687900 140270 688140
rect 140510 687900 140600 688140
rect 140840 687900 140930 688140
rect 141170 687900 141260 688140
rect 141500 687900 141610 688140
rect 141850 687900 141940 688140
rect 142180 687900 142270 688140
rect 142510 687900 142600 688140
rect 142840 687900 142950 688140
rect 143190 687900 143280 688140
rect 143520 687900 143610 688140
rect 143850 687900 143940 688140
rect 144180 687900 144290 688140
rect 144530 687900 144550 688140
rect 133550 687790 144550 687900
rect 133550 687550 133570 687790
rect 133810 687550 133900 687790
rect 134140 687550 134230 687790
rect 134470 687550 134560 687790
rect 134800 687550 134910 687790
rect 135150 687550 135240 687790
rect 135480 687550 135570 687790
rect 135810 687550 135900 687790
rect 136140 687550 136250 687790
rect 136490 687550 136580 687790
rect 136820 687550 136910 687790
rect 137150 687550 137240 687790
rect 137480 687550 137590 687790
rect 137830 687550 137920 687790
rect 138160 687550 138250 687790
rect 138490 687550 138580 687790
rect 138820 687550 138930 687790
rect 139170 687550 139260 687790
rect 139500 687550 139590 687790
rect 139830 687550 139920 687790
rect 140160 687550 140270 687790
rect 140510 687550 140600 687790
rect 140840 687550 140930 687790
rect 141170 687550 141260 687790
rect 141500 687550 141610 687790
rect 141850 687550 141940 687790
rect 142180 687550 142270 687790
rect 142510 687550 142600 687790
rect 142840 687550 142950 687790
rect 143190 687550 143280 687790
rect 143520 687550 143610 687790
rect 143850 687550 143940 687790
rect 144180 687550 144290 687790
rect 144530 687550 144550 687790
rect 133550 687460 144550 687550
rect 133550 687220 133570 687460
rect 133810 687220 133900 687460
rect 134140 687220 134230 687460
rect 134470 687220 134560 687460
rect 134800 687220 134910 687460
rect 135150 687220 135240 687460
rect 135480 687220 135570 687460
rect 135810 687220 135900 687460
rect 136140 687220 136250 687460
rect 136490 687220 136580 687460
rect 136820 687220 136910 687460
rect 137150 687220 137240 687460
rect 137480 687220 137590 687460
rect 137830 687220 137920 687460
rect 138160 687220 138250 687460
rect 138490 687220 138580 687460
rect 138820 687220 138930 687460
rect 139170 687220 139260 687460
rect 139500 687220 139590 687460
rect 139830 687220 139920 687460
rect 140160 687220 140270 687460
rect 140510 687220 140600 687460
rect 140840 687220 140930 687460
rect 141170 687220 141260 687460
rect 141500 687220 141610 687460
rect 141850 687220 141940 687460
rect 142180 687220 142270 687460
rect 142510 687220 142600 687460
rect 142840 687220 142950 687460
rect 143190 687220 143280 687460
rect 143520 687220 143610 687460
rect 143850 687220 143940 687460
rect 144180 687220 144290 687460
rect 144530 687220 144550 687460
rect 133550 687130 144550 687220
rect 133550 686890 133570 687130
rect 133810 686890 133900 687130
rect 134140 686890 134230 687130
rect 134470 686890 134560 687130
rect 134800 686890 134910 687130
rect 135150 686890 135240 687130
rect 135480 686890 135570 687130
rect 135810 686890 135900 687130
rect 136140 686890 136250 687130
rect 136490 686890 136580 687130
rect 136820 686890 136910 687130
rect 137150 686890 137240 687130
rect 137480 686890 137590 687130
rect 137830 686890 137920 687130
rect 138160 686890 138250 687130
rect 138490 686890 138580 687130
rect 138820 686890 138930 687130
rect 139170 686890 139260 687130
rect 139500 686890 139590 687130
rect 139830 686890 139920 687130
rect 140160 686890 140270 687130
rect 140510 686890 140600 687130
rect 140840 686890 140930 687130
rect 141170 686890 141260 687130
rect 141500 686890 141610 687130
rect 141850 686890 141940 687130
rect 142180 686890 142270 687130
rect 142510 686890 142600 687130
rect 142840 686890 142950 687130
rect 143190 686890 143280 687130
rect 143520 686890 143610 687130
rect 143850 686890 143940 687130
rect 144180 686890 144290 687130
rect 144530 686890 144550 687130
rect 133550 686800 144550 686890
rect 133550 686560 133570 686800
rect 133810 686560 133900 686800
rect 134140 686560 134230 686800
rect 134470 686560 134560 686800
rect 134800 686560 134910 686800
rect 135150 686560 135240 686800
rect 135480 686560 135570 686800
rect 135810 686560 135900 686800
rect 136140 686560 136250 686800
rect 136490 686560 136580 686800
rect 136820 686560 136910 686800
rect 137150 686560 137240 686800
rect 137480 686560 137590 686800
rect 137830 686560 137920 686800
rect 138160 686560 138250 686800
rect 138490 686560 138580 686800
rect 138820 686560 138930 686800
rect 139170 686560 139260 686800
rect 139500 686560 139590 686800
rect 139830 686560 139920 686800
rect 140160 686560 140270 686800
rect 140510 686560 140600 686800
rect 140840 686560 140930 686800
rect 141170 686560 141260 686800
rect 141500 686560 141610 686800
rect 141850 686560 141940 686800
rect 142180 686560 142270 686800
rect 142510 686560 142600 686800
rect 142840 686560 142950 686800
rect 143190 686560 143280 686800
rect 143520 686560 143610 686800
rect 143850 686560 143940 686800
rect 144180 686560 144290 686800
rect 144530 686560 144550 686800
rect 133550 686450 144550 686560
rect 133550 686210 133570 686450
rect 133810 686210 133900 686450
rect 134140 686210 134230 686450
rect 134470 686210 134560 686450
rect 134800 686210 134910 686450
rect 135150 686210 135240 686450
rect 135480 686210 135570 686450
rect 135810 686210 135900 686450
rect 136140 686210 136250 686450
rect 136490 686210 136580 686450
rect 136820 686210 136910 686450
rect 137150 686210 137240 686450
rect 137480 686210 137590 686450
rect 137830 686210 137920 686450
rect 138160 686210 138250 686450
rect 138490 686210 138580 686450
rect 138820 686210 138930 686450
rect 139170 686210 139260 686450
rect 139500 686210 139590 686450
rect 139830 686210 139920 686450
rect 140160 686210 140270 686450
rect 140510 686210 140600 686450
rect 140840 686210 140930 686450
rect 141170 686210 141260 686450
rect 141500 686210 141610 686450
rect 141850 686210 141940 686450
rect 142180 686210 142270 686450
rect 142510 686210 142600 686450
rect 142840 686210 142950 686450
rect 143190 686210 143280 686450
rect 143520 686210 143610 686450
rect 143850 686210 143940 686450
rect 144180 686210 144290 686450
rect 144530 686210 144550 686450
rect 133550 686120 144550 686210
rect 133550 685880 133570 686120
rect 133810 685880 133900 686120
rect 134140 685880 134230 686120
rect 134470 685880 134560 686120
rect 134800 685880 134910 686120
rect 135150 685880 135240 686120
rect 135480 685880 135570 686120
rect 135810 685880 135900 686120
rect 136140 685880 136250 686120
rect 136490 685880 136580 686120
rect 136820 685880 136910 686120
rect 137150 685880 137240 686120
rect 137480 685880 137590 686120
rect 137830 685880 137920 686120
rect 138160 685880 138250 686120
rect 138490 685880 138580 686120
rect 138820 685880 138930 686120
rect 139170 685880 139260 686120
rect 139500 685880 139590 686120
rect 139830 685880 139920 686120
rect 140160 685880 140270 686120
rect 140510 685880 140600 686120
rect 140840 685880 140930 686120
rect 141170 685880 141260 686120
rect 141500 685880 141610 686120
rect 141850 685880 141940 686120
rect 142180 685880 142270 686120
rect 142510 685880 142600 686120
rect 142840 685880 142950 686120
rect 143190 685880 143280 686120
rect 143520 685880 143610 686120
rect 143850 685880 143940 686120
rect 144180 685880 144290 686120
rect 144530 685880 144550 686120
rect 133550 685790 144550 685880
rect 133550 685550 133570 685790
rect 133810 685550 133900 685790
rect 134140 685550 134230 685790
rect 134470 685550 134560 685790
rect 134800 685550 134910 685790
rect 135150 685550 135240 685790
rect 135480 685550 135570 685790
rect 135810 685550 135900 685790
rect 136140 685550 136250 685790
rect 136490 685550 136580 685790
rect 136820 685550 136910 685790
rect 137150 685550 137240 685790
rect 137480 685550 137590 685790
rect 137830 685550 137920 685790
rect 138160 685550 138250 685790
rect 138490 685550 138580 685790
rect 138820 685550 138930 685790
rect 139170 685550 139260 685790
rect 139500 685550 139590 685790
rect 139830 685550 139920 685790
rect 140160 685550 140270 685790
rect 140510 685550 140600 685790
rect 140840 685550 140930 685790
rect 141170 685550 141260 685790
rect 141500 685550 141610 685790
rect 141850 685550 141940 685790
rect 142180 685550 142270 685790
rect 142510 685550 142600 685790
rect 142840 685550 142950 685790
rect 143190 685550 143280 685790
rect 143520 685550 143610 685790
rect 143850 685550 143940 685790
rect 144180 685550 144290 685790
rect 144530 685550 144550 685790
rect 133550 685460 144550 685550
rect 133550 685220 133570 685460
rect 133810 685220 133900 685460
rect 134140 685220 134230 685460
rect 134470 685220 134560 685460
rect 134800 685220 134910 685460
rect 135150 685220 135240 685460
rect 135480 685220 135570 685460
rect 135810 685220 135900 685460
rect 136140 685220 136250 685460
rect 136490 685220 136580 685460
rect 136820 685220 136910 685460
rect 137150 685220 137240 685460
rect 137480 685220 137590 685460
rect 137830 685220 137920 685460
rect 138160 685220 138250 685460
rect 138490 685220 138580 685460
rect 138820 685220 138930 685460
rect 139170 685220 139260 685460
rect 139500 685220 139590 685460
rect 139830 685220 139920 685460
rect 140160 685220 140270 685460
rect 140510 685220 140600 685460
rect 140840 685220 140930 685460
rect 141170 685220 141260 685460
rect 141500 685220 141610 685460
rect 141850 685220 141940 685460
rect 142180 685220 142270 685460
rect 142510 685220 142600 685460
rect 142840 685220 142950 685460
rect 143190 685220 143280 685460
rect 143520 685220 143610 685460
rect 143850 685220 143940 685460
rect 144180 685220 144290 685460
rect 144530 685220 144550 685460
rect 133550 685110 144550 685220
rect 133550 684870 133570 685110
rect 133810 684870 133900 685110
rect 134140 684870 134230 685110
rect 134470 684870 134560 685110
rect 134800 684870 134910 685110
rect 135150 684870 135240 685110
rect 135480 684870 135570 685110
rect 135810 684870 135900 685110
rect 136140 684870 136250 685110
rect 136490 684870 136580 685110
rect 136820 684870 136910 685110
rect 137150 684870 137240 685110
rect 137480 684870 137590 685110
rect 137830 684870 137920 685110
rect 138160 684870 138250 685110
rect 138490 684870 138580 685110
rect 138820 684870 138930 685110
rect 139170 684870 139260 685110
rect 139500 684870 139590 685110
rect 139830 684870 139920 685110
rect 140160 684870 140270 685110
rect 140510 684870 140600 685110
rect 140840 684870 140930 685110
rect 141170 684870 141260 685110
rect 141500 684870 141610 685110
rect 141850 684870 141940 685110
rect 142180 684870 142270 685110
rect 142510 684870 142600 685110
rect 142840 684870 142950 685110
rect 143190 684870 143280 685110
rect 143520 684870 143610 685110
rect 143850 684870 143940 685110
rect 144180 684870 144290 685110
rect 144530 684870 144550 685110
rect 133550 684780 144550 684870
rect 133550 684540 133570 684780
rect 133810 684540 133900 684780
rect 134140 684540 134230 684780
rect 134470 684540 134560 684780
rect 134800 684540 134910 684780
rect 135150 684540 135240 684780
rect 135480 684540 135570 684780
rect 135810 684540 135900 684780
rect 136140 684540 136250 684780
rect 136490 684540 136580 684780
rect 136820 684540 136910 684780
rect 137150 684540 137240 684780
rect 137480 684540 137590 684780
rect 137830 684540 137920 684780
rect 138160 684540 138250 684780
rect 138490 684540 138580 684780
rect 138820 684540 138930 684780
rect 139170 684540 139260 684780
rect 139500 684540 139590 684780
rect 139830 684540 139920 684780
rect 140160 684540 140270 684780
rect 140510 684540 140600 684780
rect 140840 684540 140930 684780
rect 141170 684540 141260 684780
rect 141500 684540 141610 684780
rect 141850 684540 141940 684780
rect 142180 684540 142270 684780
rect 142510 684540 142600 684780
rect 142840 684540 142950 684780
rect 143190 684540 143280 684780
rect 143520 684540 143610 684780
rect 143850 684540 143940 684780
rect 144180 684540 144290 684780
rect 144530 684540 144550 684780
rect 133550 684450 144550 684540
rect 133550 684210 133570 684450
rect 133810 684210 133900 684450
rect 134140 684210 134230 684450
rect 134470 684210 134560 684450
rect 134800 684210 134910 684450
rect 135150 684210 135240 684450
rect 135480 684210 135570 684450
rect 135810 684210 135900 684450
rect 136140 684210 136250 684450
rect 136490 684210 136580 684450
rect 136820 684210 136910 684450
rect 137150 684210 137240 684450
rect 137480 684210 137590 684450
rect 137830 684210 137920 684450
rect 138160 684210 138250 684450
rect 138490 684210 138580 684450
rect 138820 684210 138930 684450
rect 139170 684210 139260 684450
rect 139500 684210 139590 684450
rect 139830 684210 139920 684450
rect 140160 684210 140270 684450
rect 140510 684210 140600 684450
rect 140840 684210 140930 684450
rect 141170 684210 141260 684450
rect 141500 684210 141610 684450
rect 141850 684210 141940 684450
rect 142180 684210 142270 684450
rect 142510 684210 142600 684450
rect 142840 684210 142950 684450
rect 143190 684210 143280 684450
rect 143520 684210 143610 684450
rect 143850 684210 143940 684450
rect 144180 684210 144290 684450
rect 144530 684210 144550 684450
rect 133550 684120 144550 684210
rect 133550 683880 133570 684120
rect 133810 683880 133900 684120
rect 134140 683880 134230 684120
rect 134470 683880 134560 684120
rect 134800 683880 134910 684120
rect 135150 683880 135240 684120
rect 135480 683880 135570 684120
rect 135810 683880 135900 684120
rect 136140 683880 136250 684120
rect 136490 683880 136580 684120
rect 136820 683880 136910 684120
rect 137150 683880 137240 684120
rect 137480 683880 137590 684120
rect 137830 683880 137920 684120
rect 138160 683880 138250 684120
rect 138490 683880 138580 684120
rect 138820 683880 138930 684120
rect 139170 683880 139260 684120
rect 139500 683880 139590 684120
rect 139830 683880 139920 684120
rect 140160 683880 140270 684120
rect 140510 683880 140600 684120
rect 140840 683880 140930 684120
rect 141170 683880 141260 684120
rect 141500 683880 141610 684120
rect 141850 683880 141940 684120
rect 142180 683880 142270 684120
rect 142510 683880 142600 684120
rect 142840 683880 142950 684120
rect 143190 683880 143280 684120
rect 143520 683880 143610 684120
rect 143850 683880 143940 684120
rect 144180 683880 144290 684120
rect 144530 683880 144550 684120
rect 133550 683860 144550 683880
rect 144930 694840 155930 694860
rect 144930 694600 144950 694840
rect 145190 694600 145280 694840
rect 145520 694600 145610 694840
rect 145850 694600 145940 694840
rect 146180 694600 146290 694840
rect 146530 694600 146620 694840
rect 146860 694600 146950 694840
rect 147190 694600 147280 694840
rect 147520 694600 147630 694840
rect 147870 694600 147960 694840
rect 148200 694600 148290 694840
rect 148530 694600 148620 694840
rect 148860 694600 148970 694840
rect 149210 694600 149300 694840
rect 149540 694600 149630 694840
rect 149870 694600 149960 694840
rect 150200 694600 150310 694840
rect 150550 694600 150640 694840
rect 150880 694600 150970 694840
rect 151210 694600 151300 694840
rect 151540 694600 151650 694840
rect 151890 694600 151980 694840
rect 152220 694600 152310 694840
rect 152550 694600 152640 694840
rect 152880 694600 152990 694840
rect 153230 694600 153320 694840
rect 153560 694600 153650 694840
rect 153890 694600 153980 694840
rect 154220 694600 154330 694840
rect 154570 694600 154660 694840
rect 154900 694600 154990 694840
rect 155230 694600 155320 694840
rect 155560 694600 155670 694840
rect 155910 694600 155930 694840
rect 144930 694490 155930 694600
rect 144930 694250 144950 694490
rect 145190 694250 145280 694490
rect 145520 694250 145610 694490
rect 145850 694250 145940 694490
rect 146180 694250 146290 694490
rect 146530 694250 146620 694490
rect 146860 694250 146950 694490
rect 147190 694250 147280 694490
rect 147520 694250 147630 694490
rect 147870 694250 147960 694490
rect 148200 694250 148290 694490
rect 148530 694250 148620 694490
rect 148860 694250 148970 694490
rect 149210 694250 149300 694490
rect 149540 694250 149630 694490
rect 149870 694250 149960 694490
rect 150200 694250 150310 694490
rect 150550 694250 150640 694490
rect 150880 694250 150970 694490
rect 151210 694250 151300 694490
rect 151540 694250 151650 694490
rect 151890 694250 151980 694490
rect 152220 694250 152310 694490
rect 152550 694250 152640 694490
rect 152880 694250 152990 694490
rect 153230 694250 153320 694490
rect 153560 694250 153650 694490
rect 153890 694250 153980 694490
rect 154220 694250 154330 694490
rect 154570 694250 154660 694490
rect 154900 694250 154990 694490
rect 155230 694250 155320 694490
rect 155560 694250 155670 694490
rect 155910 694250 155930 694490
rect 144930 694160 155930 694250
rect 144930 693920 144950 694160
rect 145190 693920 145280 694160
rect 145520 693920 145610 694160
rect 145850 693920 145940 694160
rect 146180 693920 146290 694160
rect 146530 693920 146620 694160
rect 146860 693920 146950 694160
rect 147190 693920 147280 694160
rect 147520 693920 147630 694160
rect 147870 693920 147960 694160
rect 148200 693920 148290 694160
rect 148530 693920 148620 694160
rect 148860 693920 148970 694160
rect 149210 693920 149300 694160
rect 149540 693920 149630 694160
rect 149870 693920 149960 694160
rect 150200 693920 150310 694160
rect 150550 693920 150640 694160
rect 150880 693920 150970 694160
rect 151210 693920 151300 694160
rect 151540 693920 151650 694160
rect 151890 693920 151980 694160
rect 152220 693920 152310 694160
rect 152550 693920 152640 694160
rect 152880 693920 152990 694160
rect 153230 693920 153320 694160
rect 153560 693920 153650 694160
rect 153890 693920 153980 694160
rect 154220 693920 154330 694160
rect 154570 693920 154660 694160
rect 154900 693920 154990 694160
rect 155230 693920 155320 694160
rect 155560 693920 155670 694160
rect 155910 693920 155930 694160
rect 144930 693830 155930 693920
rect 144930 693590 144950 693830
rect 145190 693590 145280 693830
rect 145520 693590 145610 693830
rect 145850 693590 145940 693830
rect 146180 693590 146290 693830
rect 146530 693590 146620 693830
rect 146860 693590 146950 693830
rect 147190 693590 147280 693830
rect 147520 693590 147630 693830
rect 147870 693590 147960 693830
rect 148200 693590 148290 693830
rect 148530 693590 148620 693830
rect 148860 693590 148970 693830
rect 149210 693590 149300 693830
rect 149540 693590 149630 693830
rect 149870 693590 149960 693830
rect 150200 693590 150310 693830
rect 150550 693590 150640 693830
rect 150880 693590 150970 693830
rect 151210 693590 151300 693830
rect 151540 693590 151650 693830
rect 151890 693590 151980 693830
rect 152220 693590 152310 693830
rect 152550 693590 152640 693830
rect 152880 693590 152990 693830
rect 153230 693590 153320 693830
rect 153560 693590 153650 693830
rect 153890 693590 153980 693830
rect 154220 693590 154330 693830
rect 154570 693590 154660 693830
rect 154900 693590 154990 693830
rect 155230 693590 155320 693830
rect 155560 693590 155670 693830
rect 155910 693590 155930 693830
rect 144930 693500 155930 693590
rect 144930 693260 144950 693500
rect 145190 693260 145280 693500
rect 145520 693260 145610 693500
rect 145850 693260 145940 693500
rect 146180 693260 146290 693500
rect 146530 693260 146620 693500
rect 146860 693260 146950 693500
rect 147190 693260 147280 693500
rect 147520 693260 147630 693500
rect 147870 693260 147960 693500
rect 148200 693260 148290 693500
rect 148530 693260 148620 693500
rect 148860 693260 148970 693500
rect 149210 693260 149300 693500
rect 149540 693260 149630 693500
rect 149870 693260 149960 693500
rect 150200 693260 150310 693500
rect 150550 693260 150640 693500
rect 150880 693260 150970 693500
rect 151210 693260 151300 693500
rect 151540 693260 151650 693500
rect 151890 693260 151980 693500
rect 152220 693260 152310 693500
rect 152550 693260 152640 693500
rect 152880 693260 152990 693500
rect 153230 693260 153320 693500
rect 153560 693260 153650 693500
rect 153890 693260 153980 693500
rect 154220 693260 154330 693500
rect 154570 693260 154660 693500
rect 154900 693260 154990 693500
rect 155230 693260 155320 693500
rect 155560 693260 155670 693500
rect 155910 693260 155930 693500
rect 144930 693150 155930 693260
rect 144930 692910 144950 693150
rect 145190 692910 145280 693150
rect 145520 692910 145610 693150
rect 145850 692910 145940 693150
rect 146180 692910 146290 693150
rect 146530 692910 146620 693150
rect 146860 692910 146950 693150
rect 147190 692910 147280 693150
rect 147520 692910 147630 693150
rect 147870 692910 147960 693150
rect 148200 692910 148290 693150
rect 148530 692910 148620 693150
rect 148860 692910 148970 693150
rect 149210 692910 149300 693150
rect 149540 692910 149630 693150
rect 149870 692910 149960 693150
rect 150200 692910 150310 693150
rect 150550 692910 150640 693150
rect 150880 692910 150970 693150
rect 151210 692910 151300 693150
rect 151540 692910 151650 693150
rect 151890 692910 151980 693150
rect 152220 692910 152310 693150
rect 152550 692910 152640 693150
rect 152880 692910 152990 693150
rect 153230 692910 153320 693150
rect 153560 692910 153650 693150
rect 153890 692910 153980 693150
rect 154220 692910 154330 693150
rect 154570 692910 154660 693150
rect 154900 692910 154990 693150
rect 155230 692910 155320 693150
rect 155560 692910 155670 693150
rect 155910 692910 155930 693150
rect 144930 692820 155930 692910
rect 144930 692580 144950 692820
rect 145190 692580 145280 692820
rect 145520 692580 145610 692820
rect 145850 692580 145940 692820
rect 146180 692580 146290 692820
rect 146530 692580 146620 692820
rect 146860 692580 146950 692820
rect 147190 692580 147280 692820
rect 147520 692580 147630 692820
rect 147870 692580 147960 692820
rect 148200 692580 148290 692820
rect 148530 692580 148620 692820
rect 148860 692580 148970 692820
rect 149210 692580 149300 692820
rect 149540 692580 149630 692820
rect 149870 692580 149960 692820
rect 150200 692580 150310 692820
rect 150550 692580 150640 692820
rect 150880 692580 150970 692820
rect 151210 692580 151300 692820
rect 151540 692580 151650 692820
rect 151890 692580 151980 692820
rect 152220 692580 152310 692820
rect 152550 692580 152640 692820
rect 152880 692580 152990 692820
rect 153230 692580 153320 692820
rect 153560 692580 153650 692820
rect 153890 692580 153980 692820
rect 154220 692580 154330 692820
rect 154570 692580 154660 692820
rect 154900 692580 154990 692820
rect 155230 692580 155320 692820
rect 155560 692580 155670 692820
rect 155910 692580 155930 692820
rect 144930 692490 155930 692580
rect 144930 692250 144950 692490
rect 145190 692250 145280 692490
rect 145520 692250 145610 692490
rect 145850 692250 145940 692490
rect 146180 692250 146290 692490
rect 146530 692250 146620 692490
rect 146860 692250 146950 692490
rect 147190 692250 147280 692490
rect 147520 692250 147630 692490
rect 147870 692250 147960 692490
rect 148200 692250 148290 692490
rect 148530 692250 148620 692490
rect 148860 692250 148970 692490
rect 149210 692250 149300 692490
rect 149540 692250 149630 692490
rect 149870 692250 149960 692490
rect 150200 692250 150310 692490
rect 150550 692250 150640 692490
rect 150880 692250 150970 692490
rect 151210 692250 151300 692490
rect 151540 692250 151650 692490
rect 151890 692250 151980 692490
rect 152220 692250 152310 692490
rect 152550 692250 152640 692490
rect 152880 692250 152990 692490
rect 153230 692250 153320 692490
rect 153560 692250 153650 692490
rect 153890 692250 153980 692490
rect 154220 692250 154330 692490
rect 154570 692250 154660 692490
rect 154900 692250 154990 692490
rect 155230 692250 155320 692490
rect 155560 692250 155670 692490
rect 155910 692250 155930 692490
rect 144930 692160 155930 692250
rect 144930 691920 144950 692160
rect 145190 691920 145280 692160
rect 145520 691920 145610 692160
rect 145850 691920 145940 692160
rect 146180 691920 146290 692160
rect 146530 691920 146620 692160
rect 146860 691920 146950 692160
rect 147190 691920 147280 692160
rect 147520 691920 147630 692160
rect 147870 691920 147960 692160
rect 148200 691920 148290 692160
rect 148530 691920 148620 692160
rect 148860 691920 148970 692160
rect 149210 691920 149300 692160
rect 149540 691920 149630 692160
rect 149870 691920 149960 692160
rect 150200 691920 150310 692160
rect 150550 691920 150640 692160
rect 150880 691920 150970 692160
rect 151210 691920 151300 692160
rect 151540 691920 151650 692160
rect 151890 691920 151980 692160
rect 152220 691920 152310 692160
rect 152550 691920 152640 692160
rect 152880 691920 152990 692160
rect 153230 691920 153320 692160
rect 153560 691920 153650 692160
rect 153890 691920 153980 692160
rect 154220 691920 154330 692160
rect 154570 691920 154660 692160
rect 154900 691920 154990 692160
rect 155230 691920 155320 692160
rect 155560 691920 155670 692160
rect 155910 691920 155930 692160
rect 144930 691810 155930 691920
rect 144930 691570 144950 691810
rect 145190 691570 145280 691810
rect 145520 691570 145610 691810
rect 145850 691570 145940 691810
rect 146180 691570 146290 691810
rect 146530 691570 146620 691810
rect 146860 691570 146950 691810
rect 147190 691570 147280 691810
rect 147520 691570 147630 691810
rect 147870 691570 147960 691810
rect 148200 691570 148290 691810
rect 148530 691570 148620 691810
rect 148860 691570 148970 691810
rect 149210 691570 149300 691810
rect 149540 691570 149630 691810
rect 149870 691570 149960 691810
rect 150200 691570 150310 691810
rect 150550 691570 150640 691810
rect 150880 691570 150970 691810
rect 151210 691570 151300 691810
rect 151540 691570 151650 691810
rect 151890 691570 151980 691810
rect 152220 691570 152310 691810
rect 152550 691570 152640 691810
rect 152880 691570 152990 691810
rect 153230 691570 153320 691810
rect 153560 691570 153650 691810
rect 153890 691570 153980 691810
rect 154220 691570 154330 691810
rect 154570 691570 154660 691810
rect 154900 691570 154990 691810
rect 155230 691570 155320 691810
rect 155560 691570 155670 691810
rect 155910 691570 155930 691810
rect 144930 691480 155930 691570
rect 144930 691240 144950 691480
rect 145190 691240 145280 691480
rect 145520 691240 145610 691480
rect 145850 691240 145940 691480
rect 146180 691240 146290 691480
rect 146530 691240 146620 691480
rect 146860 691240 146950 691480
rect 147190 691240 147280 691480
rect 147520 691240 147630 691480
rect 147870 691240 147960 691480
rect 148200 691240 148290 691480
rect 148530 691240 148620 691480
rect 148860 691240 148970 691480
rect 149210 691240 149300 691480
rect 149540 691240 149630 691480
rect 149870 691240 149960 691480
rect 150200 691240 150310 691480
rect 150550 691240 150640 691480
rect 150880 691240 150970 691480
rect 151210 691240 151300 691480
rect 151540 691240 151650 691480
rect 151890 691240 151980 691480
rect 152220 691240 152310 691480
rect 152550 691240 152640 691480
rect 152880 691240 152990 691480
rect 153230 691240 153320 691480
rect 153560 691240 153650 691480
rect 153890 691240 153980 691480
rect 154220 691240 154330 691480
rect 154570 691240 154660 691480
rect 154900 691240 154990 691480
rect 155230 691240 155320 691480
rect 155560 691240 155670 691480
rect 155910 691240 155930 691480
rect 144930 691150 155930 691240
rect 144930 690910 144950 691150
rect 145190 690910 145280 691150
rect 145520 690910 145610 691150
rect 145850 690910 145940 691150
rect 146180 690910 146290 691150
rect 146530 690910 146620 691150
rect 146860 690910 146950 691150
rect 147190 690910 147280 691150
rect 147520 690910 147630 691150
rect 147870 690910 147960 691150
rect 148200 690910 148290 691150
rect 148530 690910 148620 691150
rect 148860 690910 148970 691150
rect 149210 690910 149300 691150
rect 149540 690910 149630 691150
rect 149870 690910 149960 691150
rect 150200 690910 150310 691150
rect 150550 690910 150640 691150
rect 150880 690910 150970 691150
rect 151210 690910 151300 691150
rect 151540 690910 151650 691150
rect 151890 690910 151980 691150
rect 152220 690910 152310 691150
rect 152550 690910 152640 691150
rect 152880 690910 152990 691150
rect 153230 690910 153320 691150
rect 153560 690910 153650 691150
rect 153890 690910 153980 691150
rect 154220 690910 154330 691150
rect 154570 690910 154660 691150
rect 154900 690910 154990 691150
rect 155230 690910 155320 691150
rect 155560 690910 155670 691150
rect 155910 690910 155930 691150
rect 144930 690820 155930 690910
rect 144930 690580 144950 690820
rect 145190 690580 145280 690820
rect 145520 690580 145610 690820
rect 145850 690580 145940 690820
rect 146180 690580 146290 690820
rect 146530 690580 146620 690820
rect 146860 690580 146950 690820
rect 147190 690580 147280 690820
rect 147520 690580 147630 690820
rect 147870 690580 147960 690820
rect 148200 690580 148290 690820
rect 148530 690580 148620 690820
rect 148860 690580 148970 690820
rect 149210 690580 149300 690820
rect 149540 690580 149630 690820
rect 149870 690580 149960 690820
rect 150200 690580 150310 690820
rect 150550 690580 150640 690820
rect 150880 690580 150970 690820
rect 151210 690580 151300 690820
rect 151540 690580 151650 690820
rect 151890 690580 151980 690820
rect 152220 690580 152310 690820
rect 152550 690580 152640 690820
rect 152880 690580 152990 690820
rect 153230 690580 153320 690820
rect 153560 690580 153650 690820
rect 153890 690580 153980 690820
rect 154220 690580 154330 690820
rect 154570 690580 154660 690820
rect 154900 690580 154990 690820
rect 155230 690580 155320 690820
rect 155560 690580 155670 690820
rect 155910 690580 155930 690820
rect 144930 690470 155930 690580
rect 144930 690230 144950 690470
rect 145190 690230 145280 690470
rect 145520 690230 145610 690470
rect 145850 690230 145940 690470
rect 146180 690230 146290 690470
rect 146530 690230 146620 690470
rect 146860 690230 146950 690470
rect 147190 690230 147280 690470
rect 147520 690230 147630 690470
rect 147870 690230 147960 690470
rect 148200 690230 148290 690470
rect 148530 690230 148620 690470
rect 148860 690230 148970 690470
rect 149210 690230 149300 690470
rect 149540 690230 149630 690470
rect 149870 690230 149960 690470
rect 150200 690230 150310 690470
rect 150550 690230 150640 690470
rect 150880 690230 150970 690470
rect 151210 690230 151300 690470
rect 151540 690230 151650 690470
rect 151890 690230 151980 690470
rect 152220 690230 152310 690470
rect 152550 690230 152640 690470
rect 152880 690230 152990 690470
rect 153230 690230 153320 690470
rect 153560 690230 153650 690470
rect 153890 690230 153980 690470
rect 154220 690230 154330 690470
rect 154570 690230 154660 690470
rect 154900 690230 154990 690470
rect 155230 690230 155320 690470
rect 155560 690230 155670 690470
rect 155910 690230 155930 690470
rect 144930 690140 155930 690230
rect 144930 689900 144950 690140
rect 145190 689900 145280 690140
rect 145520 689900 145610 690140
rect 145850 689900 145940 690140
rect 146180 689900 146290 690140
rect 146530 689900 146620 690140
rect 146860 689900 146950 690140
rect 147190 689900 147280 690140
rect 147520 689900 147630 690140
rect 147870 689900 147960 690140
rect 148200 689900 148290 690140
rect 148530 689900 148620 690140
rect 148860 689900 148970 690140
rect 149210 689900 149300 690140
rect 149540 689900 149630 690140
rect 149870 689900 149960 690140
rect 150200 689900 150310 690140
rect 150550 689900 150640 690140
rect 150880 689900 150970 690140
rect 151210 689900 151300 690140
rect 151540 689900 151650 690140
rect 151890 689900 151980 690140
rect 152220 689900 152310 690140
rect 152550 689900 152640 690140
rect 152880 689900 152990 690140
rect 153230 689900 153320 690140
rect 153560 689900 153650 690140
rect 153890 689900 153980 690140
rect 154220 689900 154330 690140
rect 154570 689900 154660 690140
rect 154900 689900 154990 690140
rect 155230 689900 155320 690140
rect 155560 689900 155670 690140
rect 155910 689900 155930 690140
rect 144930 689810 155930 689900
rect 144930 689570 144950 689810
rect 145190 689570 145280 689810
rect 145520 689570 145610 689810
rect 145850 689570 145940 689810
rect 146180 689570 146290 689810
rect 146530 689570 146620 689810
rect 146860 689570 146950 689810
rect 147190 689570 147280 689810
rect 147520 689570 147630 689810
rect 147870 689570 147960 689810
rect 148200 689570 148290 689810
rect 148530 689570 148620 689810
rect 148860 689570 148970 689810
rect 149210 689570 149300 689810
rect 149540 689570 149630 689810
rect 149870 689570 149960 689810
rect 150200 689570 150310 689810
rect 150550 689570 150640 689810
rect 150880 689570 150970 689810
rect 151210 689570 151300 689810
rect 151540 689570 151650 689810
rect 151890 689570 151980 689810
rect 152220 689570 152310 689810
rect 152550 689570 152640 689810
rect 152880 689570 152990 689810
rect 153230 689570 153320 689810
rect 153560 689570 153650 689810
rect 153890 689570 153980 689810
rect 154220 689570 154330 689810
rect 154570 689570 154660 689810
rect 154900 689570 154990 689810
rect 155230 689570 155320 689810
rect 155560 689570 155670 689810
rect 155910 689570 155930 689810
rect 144930 689480 155930 689570
rect 144930 689240 144950 689480
rect 145190 689240 145280 689480
rect 145520 689240 145610 689480
rect 145850 689240 145940 689480
rect 146180 689240 146290 689480
rect 146530 689240 146620 689480
rect 146860 689240 146950 689480
rect 147190 689240 147280 689480
rect 147520 689240 147630 689480
rect 147870 689240 147960 689480
rect 148200 689240 148290 689480
rect 148530 689240 148620 689480
rect 148860 689240 148970 689480
rect 149210 689240 149300 689480
rect 149540 689240 149630 689480
rect 149870 689240 149960 689480
rect 150200 689240 150310 689480
rect 150550 689240 150640 689480
rect 150880 689240 150970 689480
rect 151210 689240 151300 689480
rect 151540 689240 151650 689480
rect 151890 689240 151980 689480
rect 152220 689240 152310 689480
rect 152550 689240 152640 689480
rect 152880 689240 152990 689480
rect 153230 689240 153320 689480
rect 153560 689240 153650 689480
rect 153890 689240 153980 689480
rect 154220 689240 154330 689480
rect 154570 689240 154660 689480
rect 154900 689240 154990 689480
rect 155230 689240 155320 689480
rect 155560 689240 155670 689480
rect 155910 689240 155930 689480
rect 144930 689130 155930 689240
rect 144930 688890 144950 689130
rect 145190 688890 145280 689130
rect 145520 688890 145610 689130
rect 145850 688890 145940 689130
rect 146180 688890 146290 689130
rect 146530 688890 146620 689130
rect 146860 688890 146950 689130
rect 147190 688890 147280 689130
rect 147520 688890 147630 689130
rect 147870 688890 147960 689130
rect 148200 688890 148290 689130
rect 148530 688890 148620 689130
rect 148860 688890 148970 689130
rect 149210 688890 149300 689130
rect 149540 688890 149630 689130
rect 149870 688890 149960 689130
rect 150200 688890 150310 689130
rect 150550 688890 150640 689130
rect 150880 688890 150970 689130
rect 151210 688890 151300 689130
rect 151540 688890 151650 689130
rect 151890 688890 151980 689130
rect 152220 688890 152310 689130
rect 152550 688890 152640 689130
rect 152880 688890 152990 689130
rect 153230 688890 153320 689130
rect 153560 688890 153650 689130
rect 153890 688890 153980 689130
rect 154220 688890 154330 689130
rect 154570 688890 154660 689130
rect 154900 688890 154990 689130
rect 155230 688890 155320 689130
rect 155560 688890 155670 689130
rect 155910 688890 155930 689130
rect 144930 688800 155930 688890
rect 144930 688560 144950 688800
rect 145190 688560 145280 688800
rect 145520 688560 145610 688800
rect 145850 688560 145940 688800
rect 146180 688560 146290 688800
rect 146530 688560 146620 688800
rect 146860 688560 146950 688800
rect 147190 688560 147280 688800
rect 147520 688560 147630 688800
rect 147870 688560 147960 688800
rect 148200 688560 148290 688800
rect 148530 688560 148620 688800
rect 148860 688560 148970 688800
rect 149210 688560 149300 688800
rect 149540 688560 149630 688800
rect 149870 688560 149960 688800
rect 150200 688560 150310 688800
rect 150550 688560 150640 688800
rect 150880 688560 150970 688800
rect 151210 688560 151300 688800
rect 151540 688560 151650 688800
rect 151890 688560 151980 688800
rect 152220 688560 152310 688800
rect 152550 688560 152640 688800
rect 152880 688560 152990 688800
rect 153230 688560 153320 688800
rect 153560 688560 153650 688800
rect 153890 688560 153980 688800
rect 154220 688560 154330 688800
rect 154570 688560 154660 688800
rect 154900 688560 154990 688800
rect 155230 688560 155320 688800
rect 155560 688560 155670 688800
rect 155910 688560 155930 688800
rect 144930 688470 155930 688560
rect 144930 688230 144950 688470
rect 145190 688230 145280 688470
rect 145520 688230 145610 688470
rect 145850 688230 145940 688470
rect 146180 688230 146290 688470
rect 146530 688230 146620 688470
rect 146860 688230 146950 688470
rect 147190 688230 147280 688470
rect 147520 688230 147630 688470
rect 147870 688230 147960 688470
rect 148200 688230 148290 688470
rect 148530 688230 148620 688470
rect 148860 688230 148970 688470
rect 149210 688230 149300 688470
rect 149540 688230 149630 688470
rect 149870 688230 149960 688470
rect 150200 688230 150310 688470
rect 150550 688230 150640 688470
rect 150880 688230 150970 688470
rect 151210 688230 151300 688470
rect 151540 688230 151650 688470
rect 151890 688230 151980 688470
rect 152220 688230 152310 688470
rect 152550 688230 152640 688470
rect 152880 688230 152990 688470
rect 153230 688230 153320 688470
rect 153560 688230 153650 688470
rect 153890 688230 153980 688470
rect 154220 688230 154330 688470
rect 154570 688230 154660 688470
rect 154900 688230 154990 688470
rect 155230 688230 155320 688470
rect 155560 688230 155670 688470
rect 155910 688230 155930 688470
rect 144930 688140 155930 688230
rect 144930 687900 144950 688140
rect 145190 687900 145280 688140
rect 145520 687900 145610 688140
rect 145850 687900 145940 688140
rect 146180 687900 146290 688140
rect 146530 687900 146620 688140
rect 146860 687900 146950 688140
rect 147190 687900 147280 688140
rect 147520 687900 147630 688140
rect 147870 687900 147960 688140
rect 148200 687900 148290 688140
rect 148530 687900 148620 688140
rect 148860 687900 148970 688140
rect 149210 687900 149300 688140
rect 149540 687900 149630 688140
rect 149870 687900 149960 688140
rect 150200 687900 150310 688140
rect 150550 687900 150640 688140
rect 150880 687900 150970 688140
rect 151210 687900 151300 688140
rect 151540 687900 151650 688140
rect 151890 687900 151980 688140
rect 152220 687900 152310 688140
rect 152550 687900 152640 688140
rect 152880 687900 152990 688140
rect 153230 687900 153320 688140
rect 153560 687900 153650 688140
rect 153890 687900 153980 688140
rect 154220 687900 154330 688140
rect 154570 687900 154660 688140
rect 154900 687900 154990 688140
rect 155230 687900 155320 688140
rect 155560 687900 155670 688140
rect 155910 687900 155930 688140
rect 144930 687790 155930 687900
rect 144930 687550 144950 687790
rect 145190 687550 145280 687790
rect 145520 687550 145610 687790
rect 145850 687550 145940 687790
rect 146180 687550 146290 687790
rect 146530 687550 146620 687790
rect 146860 687550 146950 687790
rect 147190 687550 147280 687790
rect 147520 687550 147630 687790
rect 147870 687550 147960 687790
rect 148200 687550 148290 687790
rect 148530 687550 148620 687790
rect 148860 687550 148970 687790
rect 149210 687550 149300 687790
rect 149540 687550 149630 687790
rect 149870 687550 149960 687790
rect 150200 687550 150310 687790
rect 150550 687550 150640 687790
rect 150880 687550 150970 687790
rect 151210 687550 151300 687790
rect 151540 687550 151650 687790
rect 151890 687550 151980 687790
rect 152220 687550 152310 687790
rect 152550 687550 152640 687790
rect 152880 687550 152990 687790
rect 153230 687550 153320 687790
rect 153560 687550 153650 687790
rect 153890 687550 153980 687790
rect 154220 687550 154330 687790
rect 154570 687550 154660 687790
rect 154900 687550 154990 687790
rect 155230 687550 155320 687790
rect 155560 687550 155670 687790
rect 155910 687550 155930 687790
rect 144930 687460 155930 687550
rect 144930 687220 144950 687460
rect 145190 687220 145280 687460
rect 145520 687220 145610 687460
rect 145850 687220 145940 687460
rect 146180 687220 146290 687460
rect 146530 687220 146620 687460
rect 146860 687220 146950 687460
rect 147190 687220 147280 687460
rect 147520 687220 147630 687460
rect 147870 687220 147960 687460
rect 148200 687220 148290 687460
rect 148530 687220 148620 687460
rect 148860 687220 148970 687460
rect 149210 687220 149300 687460
rect 149540 687220 149630 687460
rect 149870 687220 149960 687460
rect 150200 687220 150310 687460
rect 150550 687220 150640 687460
rect 150880 687220 150970 687460
rect 151210 687220 151300 687460
rect 151540 687220 151650 687460
rect 151890 687220 151980 687460
rect 152220 687220 152310 687460
rect 152550 687220 152640 687460
rect 152880 687220 152990 687460
rect 153230 687220 153320 687460
rect 153560 687220 153650 687460
rect 153890 687220 153980 687460
rect 154220 687220 154330 687460
rect 154570 687220 154660 687460
rect 154900 687220 154990 687460
rect 155230 687220 155320 687460
rect 155560 687220 155670 687460
rect 155910 687220 155930 687460
rect 144930 687130 155930 687220
rect 144930 686890 144950 687130
rect 145190 686890 145280 687130
rect 145520 686890 145610 687130
rect 145850 686890 145940 687130
rect 146180 686890 146290 687130
rect 146530 686890 146620 687130
rect 146860 686890 146950 687130
rect 147190 686890 147280 687130
rect 147520 686890 147630 687130
rect 147870 686890 147960 687130
rect 148200 686890 148290 687130
rect 148530 686890 148620 687130
rect 148860 686890 148970 687130
rect 149210 686890 149300 687130
rect 149540 686890 149630 687130
rect 149870 686890 149960 687130
rect 150200 686890 150310 687130
rect 150550 686890 150640 687130
rect 150880 686890 150970 687130
rect 151210 686890 151300 687130
rect 151540 686890 151650 687130
rect 151890 686890 151980 687130
rect 152220 686890 152310 687130
rect 152550 686890 152640 687130
rect 152880 686890 152990 687130
rect 153230 686890 153320 687130
rect 153560 686890 153650 687130
rect 153890 686890 153980 687130
rect 154220 686890 154330 687130
rect 154570 686890 154660 687130
rect 154900 686890 154990 687130
rect 155230 686890 155320 687130
rect 155560 686890 155670 687130
rect 155910 686890 155930 687130
rect 144930 686800 155930 686890
rect 144930 686560 144950 686800
rect 145190 686560 145280 686800
rect 145520 686560 145610 686800
rect 145850 686560 145940 686800
rect 146180 686560 146290 686800
rect 146530 686560 146620 686800
rect 146860 686560 146950 686800
rect 147190 686560 147280 686800
rect 147520 686560 147630 686800
rect 147870 686560 147960 686800
rect 148200 686560 148290 686800
rect 148530 686560 148620 686800
rect 148860 686560 148970 686800
rect 149210 686560 149300 686800
rect 149540 686560 149630 686800
rect 149870 686560 149960 686800
rect 150200 686560 150310 686800
rect 150550 686560 150640 686800
rect 150880 686560 150970 686800
rect 151210 686560 151300 686800
rect 151540 686560 151650 686800
rect 151890 686560 151980 686800
rect 152220 686560 152310 686800
rect 152550 686560 152640 686800
rect 152880 686560 152990 686800
rect 153230 686560 153320 686800
rect 153560 686560 153650 686800
rect 153890 686560 153980 686800
rect 154220 686560 154330 686800
rect 154570 686560 154660 686800
rect 154900 686560 154990 686800
rect 155230 686560 155320 686800
rect 155560 686560 155670 686800
rect 155910 686560 155930 686800
rect 144930 686450 155930 686560
rect 144930 686210 144950 686450
rect 145190 686210 145280 686450
rect 145520 686210 145610 686450
rect 145850 686210 145940 686450
rect 146180 686210 146290 686450
rect 146530 686210 146620 686450
rect 146860 686210 146950 686450
rect 147190 686210 147280 686450
rect 147520 686210 147630 686450
rect 147870 686210 147960 686450
rect 148200 686210 148290 686450
rect 148530 686210 148620 686450
rect 148860 686210 148970 686450
rect 149210 686210 149300 686450
rect 149540 686210 149630 686450
rect 149870 686210 149960 686450
rect 150200 686210 150310 686450
rect 150550 686210 150640 686450
rect 150880 686210 150970 686450
rect 151210 686210 151300 686450
rect 151540 686210 151650 686450
rect 151890 686210 151980 686450
rect 152220 686210 152310 686450
rect 152550 686210 152640 686450
rect 152880 686210 152990 686450
rect 153230 686210 153320 686450
rect 153560 686210 153650 686450
rect 153890 686210 153980 686450
rect 154220 686210 154330 686450
rect 154570 686210 154660 686450
rect 154900 686210 154990 686450
rect 155230 686210 155320 686450
rect 155560 686210 155670 686450
rect 155910 686210 155930 686450
rect 144930 686120 155930 686210
rect 144930 685880 144950 686120
rect 145190 685880 145280 686120
rect 145520 685880 145610 686120
rect 145850 685880 145940 686120
rect 146180 685880 146290 686120
rect 146530 685880 146620 686120
rect 146860 685880 146950 686120
rect 147190 685880 147280 686120
rect 147520 685880 147630 686120
rect 147870 685880 147960 686120
rect 148200 685880 148290 686120
rect 148530 685880 148620 686120
rect 148860 685880 148970 686120
rect 149210 685880 149300 686120
rect 149540 685880 149630 686120
rect 149870 685880 149960 686120
rect 150200 685880 150310 686120
rect 150550 685880 150640 686120
rect 150880 685880 150970 686120
rect 151210 685880 151300 686120
rect 151540 685880 151650 686120
rect 151890 685880 151980 686120
rect 152220 685880 152310 686120
rect 152550 685880 152640 686120
rect 152880 685880 152990 686120
rect 153230 685880 153320 686120
rect 153560 685880 153650 686120
rect 153890 685880 153980 686120
rect 154220 685880 154330 686120
rect 154570 685880 154660 686120
rect 154900 685880 154990 686120
rect 155230 685880 155320 686120
rect 155560 685880 155670 686120
rect 155910 685880 155930 686120
rect 144930 685790 155930 685880
rect 144930 685550 144950 685790
rect 145190 685550 145280 685790
rect 145520 685550 145610 685790
rect 145850 685550 145940 685790
rect 146180 685550 146290 685790
rect 146530 685550 146620 685790
rect 146860 685550 146950 685790
rect 147190 685550 147280 685790
rect 147520 685550 147630 685790
rect 147870 685550 147960 685790
rect 148200 685550 148290 685790
rect 148530 685550 148620 685790
rect 148860 685550 148970 685790
rect 149210 685550 149300 685790
rect 149540 685550 149630 685790
rect 149870 685550 149960 685790
rect 150200 685550 150310 685790
rect 150550 685550 150640 685790
rect 150880 685550 150970 685790
rect 151210 685550 151300 685790
rect 151540 685550 151650 685790
rect 151890 685550 151980 685790
rect 152220 685550 152310 685790
rect 152550 685550 152640 685790
rect 152880 685550 152990 685790
rect 153230 685550 153320 685790
rect 153560 685550 153650 685790
rect 153890 685550 153980 685790
rect 154220 685550 154330 685790
rect 154570 685550 154660 685790
rect 154900 685550 154990 685790
rect 155230 685550 155320 685790
rect 155560 685550 155670 685790
rect 155910 685550 155930 685790
rect 144930 685460 155930 685550
rect 144930 685220 144950 685460
rect 145190 685220 145280 685460
rect 145520 685220 145610 685460
rect 145850 685220 145940 685460
rect 146180 685220 146290 685460
rect 146530 685220 146620 685460
rect 146860 685220 146950 685460
rect 147190 685220 147280 685460
rect 147520 685220 147630 685460
rect 147870 685220 147960 685460
rect 148200 685220 148290 685460
rect 148530 685220 148620 685460
rect 148860 685220 148970 685460
rect 149210 685220 149300 685460
rect 149540 685220 149630 685460
rect 149870 685220 149960 685460
rect 150200 685220 150310 685460
rect 150550 685220 150640 685460
rect 150880 685220 150970 685460
rect 151210 685220 151300 685460
rect 151540 685220 151650 685460
rect 151890 685220 151980 685460
rect 152220 685220 152310 685460
rect 152550 685220 152640 685460
rect 152880 685220 152990 685460
rect 153230 685220 153320 685460
rect 153560 685220 153650 685460
rect 153890 685220 153980 685460
rect 154220 685220 154330 685460
rect 154570 685220 154660 685460
rect 154900 685220 154990 685460
rect 155230 685220 155320 685460
rect 155560 685220 155670 685460
rect 155910 685220 155930 685460
rect 144930 685110 155930 685220
rect 144930 684870 144950 685110
rect 145190 684870 145280 685110
rect 145520 684870 145610 685110
rect 145850 684870 145940 685110
rect 146180 684870 146290 685110
rect 146530 684870 146620 685110
rect 146860 684870 146950 685110
rect 147190 684870 147280 685110
rect 147520 684870 147630 685110
rect 147870 684870 147960 685110
rect 148200 684870 148290 685110
rect 148530 684870 148620 685110
rect 148860 684870 148970 685110
rect 149210 684870 149300 685110
rect 149540 684870 149630 685110
rect 149870 684870 149960 685110
rect 150200 684870 150310 685110
rect 150550 684870 150640 685110
rect 150880 684870 150970 685110
rect 151210 684870 151300 685110
rect 151540 684870 151650 685110
rect 151890 684870 151980 685110
rect 152220 684870 152310 685110
rect 152550 684870 152640 685110
rect 152880 684870 152990 685110
rect 153230 684870 153320 685110
rect 153560 684870 153650 685110
rect 153890 684870 153980 685110
rect 154220 684870 154330 685110
rect 154570 684870 154660 685110
rect 154900 684870 154990 685110
rect 155230 684870 155320 685110
rect 155560 684870 155670 685110
rect 155910 684870 155930 685110
rect 144930 684780 155930 684870
rect 144930 684540 144950 684780
rect 145190 684540 145280 684780
rect 145520 684540 145610 684780
rect 145850 684540 145940 684780
rect 146180 684540 146290 684780
rect 146530 684540 146620 684780
rect 146860 684540 146950 684780
rect 147190 684540 147280 684780
rect 147520 684540 147630 684780
rect 147870 684540 147960 684780
rect 148200 684540 148290 684780
rect 148530 684540 148620 684780
rect 148860 684540 148970 684780
rect 149210 684540 149300 684780
rect 149540 684540 149630 684780
rect 149870 684540 149960 684780
rect 150200 684540 150310 684780
rect 150550 684540 150640 684780
rect 150880 684540 150970 684780
rect 151210 684540 151300 684780
rect 151540 684540 151650 684780
rect 151890 684540 151980 684780
rect 152220 684540 152310 684780
rect 152550 684540 152640 684780
rect 152880 684540 152990 684780
rect 153230 684540 153320 684780
rect 153560 684540 153650 684780
rect 153890 684540 153980 684780
rect 154220 684540 154330 684780
rect 154570 684540 154660 684780
rect 154900 684540 154990 684780
rect 155230 684540 155320 684780
rect 155560 684540 155670 684780
rect 155910 684540 155930 684780
rect 144930 684450 155930 684540
rect 144930 684210 144950 684450
rect 145190 684210 145280 684450
rect 145520 684210 145610 684450
rect 145850 684210 145940 684450
rect 146180 684210 146290 684450
rect 146530 684210 146620 684450
rect 146860 684210 146950 684450
rect 147190 684210 147280 684450
rect 147520 684210 147630 684450
rect 147870 684210 147960 684450
rect 148200 684210 148290 684450
rect 148530 684210 148620 684450
rect 148860 684210 148970 684450
rect 149210 684210 149300 684450
rect 149540 684210 149630 684450
rect 149870 684210 149960 684450
rect 150200 684210 150310 684450
rect 150550 684210 150640 684450
rect 150880 684210 150970 684450
rect 151210 684210 151300 684450
rect 151540 684210 151650 684450
rect 151890 684210 151980 684450
rect 152220 684210 152310 684450
rect 152550 684210 152640 684450
rect 152880 684210 152990 684450
rect 153230 684210 153320 684450
rect 153560 684210 153650 684450
rect 153890 684210 153980 684450
rect 154220 684210 154330 684450
rect 154570 684210 154660 684450
rect 154900 684210 154990 684450
rect 155230 684210 155320 684450
rect 155560 684210 155670 684450
rect 155910 684210 155930 684450
rect 144930 684120 155930 684210
rect 144930 683880 144950 684120
rect 145190 683880 145280 684120
rect 145520 683880 145610 684120
rect 145850 683880 145940 684120
rect 146180 683880 146290 684120
rect 146530 683880 146620 684120
rect 146860 683880 146950 684120
rect 147190 683880 147280 684120
rect 147520 683880 147630 684120
rect 147870 683880 147960 684120
rect 148200 683880 148290 684120
rect 148530 683880 148620 684120
rect 148860 683880 148970 684120
rect 149210 683880 149300 684120
rect 149540 683880 149630 684120
rect 149870 683880 149960 684120
rect 150200 683880 150310 684120
rect 150550 683880 150640 684120
rect 150880 683880 150970 684120
rect 151210 683880 151300 684120
rect 151540 683880 151650 684120
rect 151890 683880 151980 684120
rect 152220 683880 152310 684120
rect 152550 683880 152640 684120
rect 152880 683880 152990 684120
rect 153230 683880 153320 684120
rect 153560 683880 153650 684120
rect 153890 683880 153980 684120
rect 154220 683880 154330 684120
rect 154570 683880 154660 684120
rect 154900 683880 154990 684120
rect 155230 683880 155320 684120
rect 155560 683880 155670 684120
rect 155910 683880 155930 684120
rect 144930 683860 155930 683880
rect 110790 683280 121790 683300
rect 110790 683040 110810 683280
rect 111050 683040 111160 683280
rect 111400 683040 111490 683280
rect 111730 683040 111820 683280
rect 112060 683040 112150 683280
rect 112390 683040 112500 683280
rect 112740 683040 112830 683280
rect 113070 683040 113160 683280
rect 113400 683040 113490 683280
rect 113730 683040 113840 683280
rect 114080 683040 114170 683280
rect 114410 683040 114500 683280
rect 114740 683040 114830 683280
rect 115070 683040 115180 683280
rect 115420 683040 115510 683280
rect 115750 683040 115840 683280
rect 116080 683040 116170 683280
rect 116410 683040 116520 683280
rect 116760 683040 116850 683280
rect 117090 683040 117180 683280
rect 117420 683040 117510 683280
rect 117750 683040 117860 683280
rect 118100 683040 118190 683280
rect 118430 683040 118520 683280
rect 118760 683040 118850 683280
rect 119090 683040 119200 683280
rect 119440 683040 119530 683280
rect 119770 683040 119860 683280
rect 120100 683040 120190 683280
rect 120430 683040 120540 683280
rect 120780 683040 120870 683280
rect 121110 683040 121200 683280
rect 121440 683040 121530 683280
rect 121770 683040 121790 683280
rect 110790 682950 121790 683040
rect 110790 682710 110810 682950
rect 111050 682710 111160 682950
rect 111400 682710 111490 682950
rect 111730 682710 111820 682950
rect 112060 682710 112150 682950
rect 112390 682710 112500 682950
rect 112740 682710 112830 682950
rect 113070 682710 113160 682950
rect 113400 682710 113490 682950
rect 113730 682710 113840 682950
rect 114080 682710 114170 682950
rect 114410 682710 114500 682950
rect 114740 682710 114830 682950
rect 115070 682710 115180 682950
rect 115420 682710 115510 682950
rect 115750 682710 115840 682950
rect 116080 682710 116170 682950
rect 116410 682710 116520 682950
rect 116760 682710 116850 682950
rect 117090 682710 117180 682950
rect 117420 682710 117510 682950
rect 117750 682710 117860 682950
rect 118100 682710 118190 682950
rect 118430 682710 118520 682950
rect 118760 682710 118850 682950
rect 119090 682710 119200 682950
rect 119440 682710 119530 682950
rect 119770 682710 119860 682950
rect 120100 682710 120190 682950
rect 120430 682710 120540 682950
rect 120780 682710 120870 682950
rect 121110 682710 121200 682950
rect 121440 682710 121530 682950
rect 121770 682710 121790 682950
rect 110790 682620 121790 682710
rect 110790 682380 110810 682620
rect 111050 682380 111160 682620
rect 111400 682380 111490 682620
rect 111730 682380 111820 682620
rect 112060 682380 112150 682620
rect 112390 682380 112500 682620
rect 112740 682380 112830 682620
rect 113070 682380 113160 682620
rect 113400 682380 113490 682620
rect 113730 682380 113840 682620
rect 114080 682380 114170 682620
rect 114410 682380 114500 682620
rect 114740 682380 114830 682620
rect 115070 682380 115180 682620
rect 115420 682380 115510 682620
rect 115750 682380 115840 682620
rect 116080 682380 116170 682620
rect 116410 682380 116520 682620
rect 116760 682380 116850 682620
rect 117090 682380 117180 682620
rect 117420 682380 117510 682620
rect 117750 682380 117860 682620
rect 118100 682380 118190 682620
rect 118430 682380 118520 682620
rect 118760 682380 118850 682620
rect 119090 682380 119200 682620
rect 119440 682380 119530 682620
rect 119770 682380 119860 682620
rect 120100 682380 120190 682620
rect 120430 682380 120540 682620
rect 120780 682380 120870 682620
rect 121110 682380 121200 682620
rect 121440 682380 121530 682620
rect 121770 682380 121790 682620
rect 110790 682290 121790 682380
rect 110790 682050 110810 682290
rect 111050 682050 111160 682290
rect 111400 682050 111490 682290
rect 111730 682050 111820 682290
rect 112060 682050 112150 682290
rect 112390 682050 112500 682290
rect 112740 682050 112830 682290
rect 113070 682050 113160 682290
rect 113400 682050 113490 682290
rect 113730 682050 113840 682290
rect 114080 682050 114170 682290
rect 114410 682050 114500 682290
rect 114740 682050 114830 682290
rect 115070 682050 115180 682290
rect 115420 682050 115510 682290
rect 115750 682050 115840 682290
rect 116080 682050 116170 682290
rect 116410 682050 116520 682290
rect 116760 682050 116850 682290
rect 117090 682050 117180 682290
rect 117420 682050 117510 682290
rect 117750 682050 117860 682290
rect 118100 682050 118190 682290
rect 118430 682050 118520 682290
rect 118760 682050 118850 682290
rect 119090 682050 119200 682290
rect 119440 682050 119530 682290
rect 119770 682050 119860 682290
rect 120100 682050 120190 682290
rect 120430 682050 120540 682290
rect 120780 682050 120870 682290
rect 121110 682050 121200 682290
rect 121440 682050 121530 682290
rect 121770 682050 121790 682290
rect 110790 681940 121790 682050
rect 110790 681700 110810 681940
rect 111050 681700 111160 681940
rect 111400 681700 111490 681940
rect 111730 681700 111820 681940
rect 112060 681700 112150 681940
rect 112390 681700 112500 681940
rect 112740 681700 112830 681940
rect 113070 681700 113160 681940
rect 113400 681700 113490 681940
rect 113730 681700 113840 681940
rect 114080 681700 114170 681940
rect 114410 681700 114500 681940
rect 114740 681700 114830 681940
rect 115070 681700 115180 681940
rect 115420 681700 115510 681940
rect 115750 681700 115840 681940
rect 116080 681700 116170 681940
rect 116410 681700 116520 681940
rect 116760 681700 116850 681940
rect 117090 681700 117180 681940
rect 117420 681700 117510 681940
rect 117750 681700 117860 681940
rect 118100 681700 118190 681940
rect 118430 681700 118520 681940
rect 118760 681700 118850 681940
rect 119090 681700 119200 681940
rect 119440 681700 119530 681940
rect 119770 681700 119860 681940
rect 120100 681700 120190 681940
rect 120430 681700 120540 681940
rect 120780 681700 120870 681940
rect 121110 681700 121200 681940
rect 121440 681700 121530 681940
rect 121770 681700 121790 681940
rect 110790 681610 121790 681700
rect 110790 681370 110810 681610
rect 111050 681370 111160 681610
rect 111400 681370 111490 681610
rect 111730 681370 111820 681610
rect 112060 681370 112150 681610
rect 112390 681370 112500 681610
rect 112740 681370 112830 681610
rect 113070 681370 113160 681610
rect 113400 681370 113490 681610
rect 113730 681370 113840 681610
rect 114080 681370 114170 681610
rect 114410 681370 114500 681610
rect 114740 681370 114830 681610
rect 115070 681370 115180 681610
rect 115420 681370 115510 681610
rect 115750 681370 115840 681610
rect 116080 681370 116170 681610
rect 116410 681370 116520 681610
rect 116760 681370 116850 681610
rect 117090 681370 117180 681610
rect 117420 681370 117510 681610
rect 117750 681370 117860 681610
rect 118100 681370 118190 681610
rect 118430 681370 118520 681610
rect 118760 681370 118850 681610
rect 119090 681370 119200 681610
rect 119440 681370 119530 681610
rect 119770 681370 119860 681610
rect 120100 681370 120190 681610
rect 120430 681370 120540 681610
rect 120780 681370 120870 681610
rect 121110 681370 121200 681610
rect 121440 681370 121530 681610
rect 121770 681370 121790 681610
rect 110790 681280 121790 681370
rect 110790 681040 110810 681280
rect 111050 681040 111160 681280
rect 111400 681040 111490 681280
rect 111730 681040 111820 681280
rect 112060 681040 112150 681280
rect 112390 681040 112500 681280
rect 112740 681040 112830 681280
rect 113070 681040 113160 681280
rect 113400 681040 113490 681280
rect 113730 681040 113840 681280
rect 114080 681040 114170 681280
rect 114410 681040 114500 681280
rect 114740 681040 114830 681280
rect 115070 681040 115180 681280
rect 115420 681040 115510 681280
rect 115750 681040 115840 681280
rect 116080 681040 116170 681280
rect 116410 681040 116520 681280
rect 116760 681040 116850 681280
rect 117090 681040 117180 681280
rect 117420 681040 117510 681280
rect 117750 681040 117860 681280
rect 118100 681040 118190 681280
rect 118430 681040 118520 681280
rect 118760 681040 118850 681280
rect 119090 681040 119200 681280
rect 119440 681040 119530 681280
rect 119770 681040 119860 681280
rect 120100 681040 120190 681280
rect 120430 681040 120540 681280
rect 120780 681040 120870 681280
rect 121110 681040 121200 681280
rect 121440 681040 121530 681280
rect 121770 681040 121790 681280
rect 110790 680950 121790 681040
rect 110790 680710 110810 680950
rect 111050 680710 111160 680950
rect 111400 680710 111490 680950
rect 111730 680710 111820 680950
rect 112060 680710 112150 680950
rect 112390 680710 112500 680950
rect 112740 680710 112830 680950
rect 113070 680710 113160 680950
rect 113400 680710 113490 680950
rect 113730 680710 113840 680950
rect 114080 680710 114170 680950
rect 114410 680710 114500 680950
rect 114740 680710 114830 680950
rect 115070 680710 115180 680950
rect 115420 680710 115510 680950
rect 115750 680710 115840 680950
rect 116080 680710 116170 680950
rect 116410 680710 116520 680950
rect 116760 680710 116850 680950
rect 117090 680710 117180 680950
rect 117420 680710 117510 680950
rect 117750 680710 117860 680950
rect 118100 680710 118190 680950
rect 118430 680710 118520 680950
rect 118760 680710 118850 680950
rect 119090 680710 119200 680950
rect 119440 680710 119530 680950
rect 119770 680710 119860 680950
rect 120100 680710 120190 680950
rect 120430 680710 120540 680950
rect 120780 680710 120870 680950
rect 121110 680710 121200 680950
rect 121440 680710 121530 680950
rect 121770 680710 121790 680950
rect 110790 680600 121790 680710
rect 110790 680360 110810 680600
rect 111050 680360 111160 680600
rect 111400 680360 111490 680600
rect 111730 680360 111820 680600
rect 112060 680360 112150 680600
rect 112390 680360 112500 680600
rect 112740 680360 112830 680600
rect 113070 680360 113160 680600
rect 113400 680360 113490 680600
rect 113730 680360 113840 680600
rect 114080 680360 114170 680600
rect 114410 680360 114500 680600
rect 114740 680360 114830 680600
rect 115070 680360 115180 680600
rect 115420 680360 115510 680600
rect 115750 680360 115840 680600
rect 116080 680360 116170 680600
rect 116410 680360 116520 680600
rect 116760 680360 116850 680600
rect 117090 680360 117180 680600
rect 117420 680360 117510 680600
rect 117750 680360 117860 680600
rect 118100 680360 118190 680600
rect 118430 680360 118520 680600
rect 118760 680360 118850 680600
rect 119090 680360 119200 680600
rect 119440 680360 119530 680600
rect 119770 680360 119860 680600
rect 120100 680360 120190 680600
rect 120430 680360 120540 680600
rect 120780 680360 120870 680600
rect 121110 680360 121200 680600
rect 121440 680360 121530 680600
rect 121770 680360 121790 680600
rect 110790 680270 121790 680360
rect 110790 680030 110810 680270
rect 111050 680030 111160 680270
rect 111400 680030 111490 680270
rect 111730 680030 111820 680270
rect 112060 680030 112150 680270
rect 112390 680030 112500 680270
rect 112740 680030 112830 680270
rect 113070 680030 113160 680270
rect 113400 680030 113490 680270
rect 113730 680030 113840 680270
rect 114080 680030 114170 680270
rect 114410 680030 114500 680270
rect 114740 680030 114830 680270
rect 115070 680030 115180 680270
rect 115420 680030 115510 680270
rect 115750 680030 115840 680270
rect 116080 680030 116170 680270
rect 116410 680030 116520 680270
rect 116760 680030 116850 680270
rect 117090 680030 117180 680270
rect 117420 680030 117510 680270
rect 117750 680030 117860 680270
rect 118100 680030 118190 680270
rect 118430 680030 118520 680270
rect 118760 680030 118850 680270
rect 119090 680030 119200 680270
rect 119440 680030 119530 680270
rect 119770 680030 119860 680270
rect 120100 680030 120190 680270
rect 120430 680030 120540 680270
rect 120780 680030 120870 680270
rect 121110 680030 121200 680270
rect 121440 680030 121530 680270
rect 121770 680030 121790 680270
rect 110790 679940 121790 680030
rect 110790 679700 110810 679940
rect 111050 679700 111160 679940
rect 111400 679700 111490 679940
rect 111730 679700 111820 679940
rect 112060 679700 112150 679940
rect 112390 679700 112500 679940
rect 112740 679700 112830 679940
rect 113070 679700 113160 679940
rect 113400 679700 113490 679940
rect 113730 679700 113840 679940
rect 114080 679700 114170 679940
rect 114410 679700 114500 679940
rect 114740 679700 114830 679940
rect 115070 679700 115180 679940
rect 115420 679700 115510 679940
rect 115750 679700 115840 679940
rect 116080 679700 116170 679940
rect 116410 679700 116520 679940
rect 116760 679700 116850 679940
rect 117090 679700 117180 679940
rect 117420 679700 117510 679940
rect 117750 679700 117860 679940
rect 118100 679700 118190 679940
rect 118430 679700 118520 679940
rect 118760 679700 118850 679940
rect 119090 679700 119200 679940
rect 119440 679700 119530 679940
rect 119770 679700 119860 679940
rect 120100 679700 120190 679940
rect 120430 679700 120540 679940
rect 120780 679700 120870 679940
rect 121110 679700 121200 679940
rect 121440 679700 121530 679940
rect 121770 679700 121790 679940
rect 110790 679610 121790 679700
rect 110790 679370 110810 679610
rect 111050 679370 111160 679610
rect 111400 679370 111490 679610
rect 111730 679370 111820 679610
rect 112060 679370 112150 679610
rect 112390 679370 112500 679610
rect 112740 679370 112830 679610
rect 113070 679370 113160 679610
rect 113400 679370 113490 679610
rect 113730 679370 113840 679610
rect 114080 679370 114170 679610
rect 114410 679370 114500 679610
rect 114740 679370 114830 679610
rect 115070 679370 115180 679610
rect 115420 679370 115510 679610
rect 115750 679370 115840 679610
rect 116080 679370 116170 679610
rect 116410 679370 116520 679610
rect 116760 679370 116850 679610
rect 117090 679370 117180 679610
rect 117420 679370 117510 679610
rect 117750 679370 117860 679610
rect 118100 679370 118190 679610
rect 118430 679370 118520 679610
rect 118760 679370 118850 679610
rect 119090 679370 119200 679610
rect 119440 679370 119530 679610
rect 119770 679370 119860 679610
rect 120100 679370 120190 679610
rect 120430 679370 120540 679610
rect 120780 679370 120870 679610
rect 121110 679370 121200 679610
rect 121440 679370 121530 679610
rect 121770 679370 121790 679610
rect 110790 679260 121790 679370
rect 110790 679020 110810 679260
rect 111050 679020 111160 679260
rect 111400 679020 111490 679260
rect 111730 679020 111820 679260
rect 112060 679020 112150 679260
rect 112390 679020 112500 679260
rect 112740 679020 112830 679260
rect 113070 679020 113160 679260
rect 113400 679020 113490 679260
rect 113730 679020 113840 679260
rect 114080 679020 114170 679260
rect 114410 679020 114500 679260
rect 114740 679020 114830 679260
rect 115070 679020 115180 679260
rect 115420 679020 115510 679260
rect 115750 679020 115840 679260
rect 116080 679020 116170 679260
rect 116410 679020 116520 679260
rect 116760 679020 116850 679260
rect 117090 679020 117180 679260
rect 117420 679020 117510 679260
rect 117750 679020 117860 679260
rect 118100 679020 118190 679260
rect 118430 679020 118520 679260
rect 118760 679020 118850 679260
rect 119090 679020 119200 679260
rect 119440 679020 119530 679260
rect 119770 679020 119860 679260
rect 120100 679020 120190 679260
rect 120430 679020 120540 679260
rect 120780 679020 120870 679260
rect 121110 679020 121200 679260
rect 121440 679020 121530 679260
rect 121770 679020 121790 679260
rect 110790 678930 121790 679020
rect 110790 678690 110810 678930
rect 111050 678690 111160 678930
rect 111400 678690 111490 678930
rect 111730 678690 111820 678930
rect 112060 678690 112150 678930
rect 112390 678690 112500 678930
rect 112740 678690 112830 678930
rect 113070 678690 113160 678930
rect 113400 678690 113490 678930
rect 113730 678690 113840 678930
rect 114080 678690 114170 678930
rect 114410 678690 114500 678930
rect 114740 678690 114830 678930
rect 115070 678690 115180 678930
rect 115420 678690 115510 678930
rect 115750 678690 115840 678930
rect 116080 678690 116170 678930
rect 116410 678690 116520 678930
rect 116760 678690 116850 678930
rect 117090 678690 117180 678930
rect 117420 678690 117510 678930
rect 117750 678690 117860 678930
rect 118100 678690 118190 678930
rect 118430 678690 118520 678930
rect 118760 678690 118850 678930
rect 119090 678690 119200 678930
rect 119440 678690 119530 678930
rect 119770 678690 119860 678930
rect 120100 678690 120190 678930
rect 120430 678690 120540 678930
rect 120780 678690 120870 678930
rect 121110 678690 121200 678930
rect 121440 678690 121530 678930
rect 121770 678690 121790 678930
rect 110790 678600 121790 678690
rect 110790 678360 110810 678600
rect 111050 678360 111160 678600
rect 111400 678360 111490 678600
rect 111730 678360 111820 678600
rect 112060 678360 112150 678600
rect 112390 678360 112500 678600
rect 112740 678360 112830 678600
rect 113070 678360 113160 678600
rect 113400 678360 113490 678600
rect 113730 678360 113840 678600
rect 114080 678360 114170 678600
rect 114410 678360 114500 678600
rect 114740 678360 114830 678600
rect 115070 678360 115180 678600
rect 115420 678360 115510 678600
rect 115750 678360 115840 678600
rect 116080 678360 116170 678600
rect 116410 678360 116520 678600
rect 116760 678360 116850 678600
rect 117090 678360 117180 678600
rect 117420 678360 117510 678600
rect 117750 678360 117860 678600
rect 118100 678360 118190 678600
rect 118430 678360 118520 678600
rect 118760 678360 118850 678600
rect 119090 678360 119200 678600
rect 119440 678360 119530 678600
rect 119770 678360 119860 678600
rect 120100 678360 120190 678600
rect 120430 678360 120540 678600
rect 120780 678360 120870 678600
rect 121110 678360 121200 678600
rect 121440 678360 121530 678600
rect 121770 678360 121790 678600
rect 110790 678270 121790 678360
rect 110790 678030 110810 678270
rect 111050 678030 111160 678270
rect 111400 678030 111490 678270
rect 111730 678030 111820 678270
rect 112060 678030 112150 678270
rect 112390 678030 112500 678270
rect 112740 678030 112830 678270
rect 113070 678030 113160 678270
rect 113400 678030 113490 678270
rect 113730 678030 113840 678270
rect 114080 678030 114170 678270
rect 114410 678030 114500 678270
rect 114740 678030 114830 678270
rect 115070 678030 115180 678270
rect 115420 678030 115510 678270
rect 115750 678030 115840 678270
rect 116080 678030 116170 678270
rect 116410 678030 116520 678270
rect 116760 678030 116850 678270
rect 117090 678030 117180 678270
rect 117420 678030 117510 678270
rect 117750 678030 117860 678270
rect 118100 678030 118190 678270
rect 118430 678030 118520 678270
rect 118760 678030 118850 678270
rect 119090 678030 119200 678270
rect 119440 678030 119530 678270
rect 119770 678030 119860 678270
rect 120100 678030 120190 678270
rect 120430 678030 120540 678270
rect 120780 678030 120870 678270
rect 121110 678030 121200 678270
rect 121440 678030 121530 678270
rect 121770 678030 121790 678270
rect 110790 677920 121790 678030
rect 110790 677680 110810 677920
rect 111050 677680 111160 677920
rect 111400 677680 111490 677920
rect 111730 677680 111820 677920
rect 112060 677680 112150 677920
rect 112390 677680 112500 677920
rect 112740 677680 112830 677920
rect 113070 677680 113160 677920
rect 113400 677680 113490 677920
rect 113730 677680 113840 677920
rect 114080 677680 114170 677920
rect 114410 677680 114500 677920
rect 114740 677680 114830 677920
rect 115070 677680 115180 677920
rect 115420 677680 115510 677920
rect 115750 677680 115840 677920
rect 116080 677680 116170 677920
rect 116410 677680 116520 677920
rect 116760 677680 116850 677920
rect 117090 677680 117180 677920
rect 117420 677680 117510 677920
rect 117750 677680 117860 677920
rect 118100 677680 118190 677920
rect 118430 677680 118520 677920
rect 118760 677680 118850 677920
rect 119090 677680 119200 677920
rect 119440 677680 119530 677920
rect 119770 677680 119860 677920
rect 120100 677680 120190 677920
rect 120430 677680 120540 677920
rect 120780 677680 120870 677920
rect 121110 677680 121200 677920
rect 121440 677680 121530 677920
rect 121770 677680 121790 677920
rect 110790 677590 121790 677680
rect 110790 677350 110810 677590
rect 111050 677350 111160 677590
rect 111400 677350 111490 677590
rect 111730 677350 111820 677590
rect 112060 677350 112150 677590
rect 112390 677350 112500 677590
rect 112740 677350 112830 677590
rect 113070 677350 113160 677590
rect 113400 677350 113490 677590
rect 113730 677350 113840 677590
rect 114080 677350 114170 677590
rect 114410 677350 114500 677590
rect 114740 677350 114830 677590
rect 115070 677350 115180 677590
rect 115420 677350 115510 677590
rect 115750 677350 115840 677590
rect 116080 677350 116170 677590
rect 116410 677350 116520 677590
rect 116760 677350 116850 677590
rect 117090 677350 117180 677590
rect 117420 677350 117510 677590
rect 117750 677350 117860 677590
rect 118100 677350 118190 677590
rect 118430 677350 118520 677590
rect 118760 677350 118850 677590
rect 119090 677350 119200 677590
rect 119440 677350 119530 677590
rect 119770 677350 119860 677590
rect 120100 677350 120190 677590
rect 120430 677350 120540 677590
rect 120780 677350 120870 677590
rect 121110 677350 121200 677590
rect 121440 677350 121530 677590
rect 121770 677350 121790 677590
rect 110790 677260 121790 677350
rect 110790 677020 110810 677260
rect 111050 677020 111160 677260
rect 111400 677020 111490 677260
rect 111730 677020 111820 677260
rect 112060 677020 112150 677260
rect 112390 677020 112500 677260
rect 112740 677020 112830 677260
rect 113070 677020 113160 677260
rect 113400 677020 113490 677260
rect 113730 677020 113840 677260
rect 114080 677020 114170 677260
rect 114410 677020 114500 677260
rect 114740 677020 114830 677260
rect 115070 677020 115180 677260
rect 115420 677020 115510 677260
rect 115750 677020 115840 677260
rect 116080 677020 116170 677260
rect 116410 677020 116520 677260
rect 116760 677020 116850 677260
rect 117090 677020 117180 677260
rect 117420 677020 117510 677260
rect 117750 677020 117860 677260
rect 118100 677020 118190 677260
rect 118430 677020 118520 677260
rect 118760 677020 118850 677260
rect 119090 677020 119200 677260
rect 119440 677020 119530 677260
rect 119770 677020 119860 677260
rect 120100 677020 120190 677260
rect 120430 677020 120540 677260
rect 120780 677020 120870 677260
rect 121110 677020 121200 677260
rect 121440 677020 121530 677260
rect 121770 677020 121790 677260
rect 110790 676930 121790 677020
rect 110790 676690 110810 676930
rect 111050 676690 111160 676930
rect 111400 676690 111490 676930
rect 111730 676690 111820 676930
rect 112060 676690 112150 676930
rect 112390 676690 112500 676930
rect 112740 676690 112830 676930
rect 113070 676690 113160 676930
rect 113400 676690 113490 676930
rect 113730 676690 113840 676930
rect 114080 676690 114170 676930
rect 114410 676690 114500 676930
rect 114740 676690 114830 676930
rect 115070 676690 115180 676930
rect 115420 676690 115510 676930
rect 115750 676690 115840 676930
rect 116080 676690 116170 676930
rect 116410 676690 116520 676930
rect 116760 676690 116850 676930
rect 117090 676690 117180 676930
rect 117420 676690 117510 676930
rect 117750 676690 117860 676930
rect 118100 676690 118190 676930
rect 118430 676690 118520 676930
rect 118760 676690 118850 676930
rect 119090 676690 119200 676930
rect 119440 676690 119530 676930
rect 119770 676690 119860 676930
rect 120100 676690 120190 676930
rect 120430 676690 120540 676930
rect 120780 676690 120870 676930
rect 121110 676690 121200 676930
rect 121440 676690 121530 676930
rect 121770 676690 121790 676930
rect 110790 676580 121790 676690
rect 110790 676340 110810 676580
rect 111050 676340 111160 676580
rect 111400 676340 111490 676580
rect 111730 676340 111820 676580
rect 112060 676340 112150 676580
rect 112390 676340 112500 676580
rect 112740 676340 112830 676580
rect 113070 676340 113160 676580
rect 113400 676340 113490 676580
rect 113730 676340 113840 676580
rect 114080 676340 114170 676580
rect 114410 676340 114500 676580
rect 114740 676340 114830 676580
rect 115070 676340 115180 676580
rect 115420 676340 115510 676580
rect 115750 676340 115840 676580
rect 116080 676340 116170 676580
rect 116410 676340 116520 676580
rect 116760 676340 116850 676580
rect 117090 676340 117180 676580
rect 117420 676340 117510 676580
rect 117750 676340 117860 676580
rect 118100 676340 118190 676580
rect 118430 676340 118520 676580
rect 118760 676340 118850 676580
rect 119090 676340 119200 676580
rect 119440 676340 119530 676580
rect 119770 676340 119860 676580
rect 120100 676340 120190 676580
rect 120430 676340 120540 676580
rect 120780 676340 120870 676580
rect 121110 676340 121200 676580
rect 121440 676340 121530 676580
rect 121770 676340 121790 676580
rect 110790 676250 121790 676340
rect 110790 676010 110810 676250
rect 111050 676010 111160 676250
rect 111400 676010 111490 676250
rect 111730 676010 111820 676250
rect 112060 676010 112150 676250
rect 112390 676010 112500 676250
rect 112740 676010 112830 676250
rect 113070 676010 113160 676250
rect 113400 676010 113490 676250
rect 113730 676010 113840 676250
rect 114080 676010 114170 676250
rect 114410 676010 114500 676250
rect 114740 676010 114830 676250
rect 115070 676010 115180 676250
rect 115420 676010 115510 676250
rect 115750 676010 115840 676250
rect 116080 676010 116170 676250
rect 116410 676010 116520 676250
rect 116760 676010 116850 676250
rect 117090 676010 117180 676250
rect 117420 676010 117510 676250
rect 117750 676010 117860 676250
rect 118100 676010 118190 676250
rect 118430 676010 118520 676250
rect 118760 676010 118850 676250
rect 119090 676010 119200 676250
rect 119440 676010 119530 676250
rect 119770 676010 119860 676250
rect 120100 676010 120190 676250
rect 120430 676010 120540 676250
rect 120780 676010 120870 676250
rect 121110 676010 121200 676250
rect 121440 676010 121530 676250
rect 121770 676010 121790 676250
rect 110790 675920 121790 676010
rect 110790 675680 110810 675920
rect 111050 675680 111160 675920
rect 111400 675680 111490 675920
rect 111730 675680 111820 675920
rect 112060 675680 112150 675920
rect 112390 675680 112500 675920
rect 112740 675680 112830 675920
rect 113070 675680 113160 675920
rect 113400 675680 113490 675920
rect 113730 675680 113840 675920
rect 114080 675680 114170 675920
rect 114410 675680 114500 675920
rect 114740 675680 114830 675920
rect 115070 675680 115180 675920
rect 115420 675680 115510 675920
rect 115750 675680 115840 675920
rect 116080 675680 116170 675920
rect 116410 675680 116520 675920
rect 116760 675680 116850 675920
rect 117090 675680 117180 675920
rect 117420 675680 117510 675920
rect 117750 675680 117860 675920
rect 118100 675680 118190 675920
rect 118430 675680 118520 675920
rect 118760 675680 118850 675920
rect 119090 675680 119200 675920
rect 119440 675680 119530 675920
rect 119770 675680 119860 675920
rect 120100 675680 120190 675920
rect 120430 675680 120540 675920
rect 120780 675680 120870 675920
rect 121110 675680 121200 675920
rect 121440 675680 121530 675920
rect 121770 675680 121790 675920
rect 110790 675590 121790 675680
rect 110790 675350 110810 675590
rect 111050 675350 111160 675590
rect 111400 675350 111490 675590
rect 111730 675350 111820 675590
rect 112060 675350 112150 675590
rect 112390 675350 112500 675590
rect 112740 675350 112830 675590
rect 113070 675350 113160 675590
rect 113400 675350 113490 675590
rect 113730 675350 113840 675590
rect 114080 675350 114170 675590
rect 114410 675350 114500 675590
rect 114740 675350 114830 675590
rect 115070 675350 115180 675590
rect 115420 675350 115510 675590
rect 115750 675350 115840 675590
rect 116080 675350 116170 675590
rect 116410 675350 116520 675590
rect 116760 675350 116850 675590
rect 117090 675350 117180 675590
rect 117420 675350 117510 675590
rect 117750 675350 117860 675590
rect 118100 675350 118190 675590
rect 118430 675350 118520 675590
rect 118760 675350 118850 675590
rect 119090 675350 119200 675590
rect 119440 675350 119530 675590
rect 119770 675350 119860 675590
rect 120100 675350 120190 675590
rect 120430 675350 120540 675590
rect 120780 675350 120870 675590
rect 121110 675350 121200 675590
rect 121440 675350 121530 675590
rect 121770 675350 121790 675590
rect 110790 675240 121790 675350
rect 110790 675000 110810 675240
rect 111050 675000 111160 675240
rect 111400 675000 111490 675240
rect 111730 675000 111820 675240
rect 112060 675000 112150 675240
rect 112390 675000 112500 675240
rect 112740 675000 112830 675240
rect 113070 675000 113160 675240
rect 113400 675000 113490 675240
rect 113730 675000 113840 675240
rect 114080 675000 114170 675240
rect 114410 675000 114500 675240
rect 114740 675000 114830 675240
rect 115070 675000 115180 675240
rect 115420 675000 115510 675240
rect 115750 675000 115840 675240
rect 116080 675000 116170 675240
rect 116410 675000 116520 675240
rect 116760 675000 116850 675240
rect 117090 675000 117180 675240
rect 117420 675000 117510 675240
rect 117750 675000 117860 675240
rect 118100 675000 118190 675240
rect 118430 675000 118520 675240
rect 118760 675000 118850 675240
rect 119090 675000 119200 675240
rect 119440 675000 119530 675240
rect 119770 675000 119860 675240
rect 120100 675000 120190 675240
rect 120430 675000 120540 675240
rect 120780 675000 120870 675240
rect 121110 675000 121200 675240
rect 121440 675000 121530 675240
rect 121770 675000 121790 675240
rect 110790 674910 121790 675000
rect 110790 674670 110810 674910
rect 111050 674670 111160 674910
rect 111400 674670 111490 674910
rect 111730 674670 111820 674910
rect 112060 674670 112150 674910
rect 112390 674670 112500 674910
rect 112740 674670 112830 674910
rect 113070 674670 113160 674910
rect 113400 674670 113490 674910
rect 113730 674670 113840 674910
rect 114080 674670 114170 674910
rect 114410 674670 114500 674910
rect 114740 674670 114830 674910
rect 115070 674670 115180 674910
rect 115420 674670 115510 674910
rect 115750 674670 115840 674910
rect 116080 674670 116170 674910
rect 116410 674670 116520 674910
rect 116760 674670 116850 674910
rect 117090 674670 117180 674910
rect 117420 674670 117510 674910
rect 117750 674670 117860 674910
rect 118100 674670 118190 674910
rect 118430 674670 118520 674910
rect 118760 674670 118850 674910
rect 119090 674670 119200 674910
rect 119440 674670 119530 674910
rect 119770 674670 119860 674910
rect 120100 674670 120190 674910
rect 120430 674670 120540 674910
rect 120780 674670 120870 674910
rect 121110 674670 121200 674910
rect 121440 674670 121530 674910
rect 121770 674670 121790 674910
rect 110790 674580 121790 674670
rect 110790 674340 110810 674580
rect 111050 674340 111160 674580
rect 111400 674340 111490 674580
rect 111730 674340 111820 674580
rect 112060 674340 112150 674580
rect 112390 674340 112500 674580
rect 112740 674340 112830 674580
rect 113070 674340 113160 674580
rect 113400 674340 113490 674580
rect 113730 674340 113840 674580
rect 114080 674340 114170 674580
rect 114410 674340 114500 674580
rect 114740 674340 114830 674580
rect 115070 674340 115180 674580
rect 115420 674340 115510 674580
rect 115750 674340 115840 674580
rect 116080 674340 116170 674580
rect 116410 674340 116520 674580
rect 116760 674340 116850 674580
rect 117090 674340 117180 674580
rect 117420 674340 117510 674580
rect 117750 674340 117860 674580
rect 118100 674340 118190 674580
rect 118430 674340 118520 674580
rect 118760 674340 118850 674580
rect 119090 674340 119200 674580
rect 119440 674340 119530 674580
rect 119770 674340 119860 674580
rect 120100 674340 120190 674580
rect 120430 674340 120540 674580
rect 120780 674340 120870 674580
rect 121110 674340 121200 674580
rect 121440 674340 121530 674580
rect 121770 674340 121790 674580
rect 110790 674250 121790 674340
rect 110790 674010 110810 674250
rect 111050 674010 111160 674250
rect 111400 674010 111490 674250
rect 111730 674010 111820 674250
rect 112060 674010 112150 674250
rect 112390 674010 112500 674250
rect 112740 674010 112830 674250
rect 113070 674010 113160 674250
rect 113400 674010 113490 674250
rect 113730 674010 113840 674250
rect 114080 674010 114170 674250
rect 114410 674010 114500 674250
rect 114740 674010 114830 674250
rect 115070 674010 115180 674250
rect 115420 674010 115510 674250
rect 115750 674010 115840 674250
rect 116080 674010 116170 674250
rect 116410 674010 116520 674250
rect 116760 674010 116850 674250
rect 117090 674010 117180 674250
rect 117420 674010 117510 674250
rect 117750 674010 117860 674250
rect 118100 674010 118190 674250
rect 118430 674010 118520 674250
rect 118760 674010 118850 674250
rect 119090 674010 119200 674250
rect 119440 674010 119530 674250
rect 119770 674010 119860 674250
rect 120100 674010 120190 674250
rect 120430 674010 120540 674250
rect 120780 674010 120870 674250
rect 121110 674010 121200 674250
rect 121440 674010 121530 674250
rect 121770 674010 121790 674250
rect 110790 673900 121790 674010
rect 110790 673660 110810 673900
rect 111050 673660 111160 673900
rect 111400 673660 111490 673900
rect 111730 673660 111820 673900
rect 112060 673660 112150 673900
rect 112390 673660 112500 673900
rect 112740 673660 112830 673900
rect 113070 673660 113160 673900
rect 113400 673660 113490 673900
rect 113730 673660 113840 673900
rect 114080 673660 114170 673900
rect 114410 673660 114500 673900
rect 114740 673660 114830 673900
rect 115070 673660 115180 673900
rect 115420 673660 115510 673900
rect 115750 673660 115840 673900
rect 116080 673660 116170 673900
rect 116410 673660 116520 673900
rect 116760 673660 116850 673900
rect 117090 673660 117180 673900
rect 117420 673660 117510 673900
rect 117750 673660 117860 673900
rect 118100 673660 118190 673900
rect 118430 673660 118520 673900
rect 118760 673660 118850 673900
rect 119090 673660 119200 673900
rect 119440 673660 119530 673900
rect 119770 673660 119860 673900
rect 120100 673660 120190 673900
rect 120430 673660 120540 673900
rect 120780 673660 120870 673900
rect 121110 673660 121200 673900
rect 121440 673660 121530 673900
rect 121770 673660 121790 673900
rect 110790 673570 121790 673660
rect 110790 673330 110810 673570
rect 111050 673330 111160 673570
rect 111400 673330 111490 673570
rect 111730 673330 111820 673570
rect 112060 673330 112150 673570
rect 112390 673330 112500 673570
rect 112740 673330 112830 673570
rect 113070 673330 113160 673570
rect 113400 673330 113490 673570
rect 113730 673330 113840 673570
rect 114080 673330 114170 673570
rect 114410 673330 114500 673570
rect 114740 673330 114830 673570
rect 115070 673330 115180 673570
rect 115420 673330 115510 673570
rect 115750 673330 115840 673570
rect 116080 673330 116170 673570
rect 116410 673330 116520 673570
rect 116760 673330 116850 673570
rect 117090 673330 117180 673570
rect 117420 673330 117510 673570
rect 117750 673330 117860 673570
rect 118100 673330 118190 673570
rect 118430 673330 118520 673570
rect 118760 673330 118850 673570
rect 119090 673330 119200 673570
rect 119440 673330 119530 673570
rect 119770 673330 119860 673570
rect 120100 673330 120190 673570
rect 120430 673330 120540 673570
rect 120780 673330 120870 673570
rect 121110 673330 121200 673570
rect 121440 673330 121530 673570
rect 121770 673330 121790 673570
rect 110790 673240 121790 673330
rect 110790 673000 110810 673240
rect 111050 673000 111160 673240
rect 111400 673000 111490 673240
rect 111730 673000 111820 673240
rect 112060 673000 112150 673240
rect 112390 673000 112500 673240
rect 112740 673000 112830 673240
rect 113070 673000 113160 673240
rect 113400 673000 113490 673240
rect 113730 673000 113840 673240
rect 114080 673000 114170 673240
rect 114410 673000 114500 673240
rect 114740 673000 114830 673240
rect 115070 673000 115180 673240
rect 115420 673000 115510 673240
rect 115750 673000 115840 673240
rect 116080 673000 116170 673240
rect 116410 673000 116520 673240
rect 116760 673000 116850 673240
rect 117090 673000 117180 673240
rect 117420 673000 117510 673240
rect 117750 673000 117860 673240
rect 118100 673000 118190 673240
rect 118430 673000 118520 673240
rect 118760 673000 118850 673240
rect 119090 673000 119200 673240
rect 119440 673000 119530 673240
rect 119770 673000 119860 673240
rect 120100 673000 120190 673240
rect 120430 673000 120540 673240
rect 120780 673000 120870 673240
rect 121110 673000 121200 673240
rect 121440 673000 121530 673240
rect 121770 673000 121790 673240
rect 110790 672910 121790 673000
rect 110790 672670 110810 672910
rect 111050 672670 111160 672910
rect 111400 672670 111490 672910
rect 111730 672670 111820 672910
rect 112060 672670 112150 672910
rect 112390 672670 112500 672910
rect 112740 672670 112830 672910
rect 113070 672670 113160 672910
rect 113400 672670 113490 672910
rect 113730 672670 113840 672910
rect 114080 672670 114170 672910
rect 114410 672670 114500 672910
rect 114740 672670 114830 672910
rect 115070 672670 115180 672910
rect 115420 672670 115510 672910
rect 115750 672670 115840 672910
rect 116080 672670 116170 672910
rect 116410 672670 116520 672910
rect 116760 672670 116850 672910
rect 117090 672670 117180 672910
rect 117420 672670 117510 672910
rect 117750 672670 117860 672910
rect 118100 672670 118190 672910
rect 118430 672670 118520 672910
rect 118760 672670 118850 672910
rect 119090 672670 119200 672910
rect 119440 672670 119530 672910
rect 119770 672670 119860 672910
rect 120100 672670 120190 672910
rect 120430 672670 120540 672910
rect 120780 672670 120870 672910
rect 121110 672670 121200 672910
rect 121440 672670 121530 672910
rect 121770 672670 121790 672910
rect 110790 672560 121790 672670
rect 110790 672320 110810 672560
rect 111050 672320 111160 672560
rect 111400 672320 111490 672560
rect 111730 672320 111820 672560
rect 112060 672320 112150 672560
rect 112390 672320 112500 672560
rect 112740 672320 112830 672560
rect 113070 672320 113160 672560
rect 113400 672320 113490 672560
rect 113730 672320 113840 672560
rect 114080 672320 114170 672560
rect 114410 672320 114500 672560
rect 114740 672320 114830 672560
rect 115070 672320 115180 672560
rect 115420 672320 115510 672560
rect 115750 672320 115840 672560
rect 116080 672320 116170 672560
rect 116410 672320 116520 672560
rect 116760 672320 116850 672560
rect 117090 672320 117180 672560
rect 117420 672320 117510 672560
rect 117750 672320 117860 672560
rect 118100 672320 118190 672560
rect 118430 672320 118520 672560
rect 118760 672320 118850 672560
rect 119090 672320 119200 672560
rect 119440 672320 119530 672560
rect 119770 672320 119860 672560
rect 120100 672320 120190 672560
rect 120430 672320 120540 672560
rect 120780 672320 120870 672560
rect 121110 672320 121200 672560
rect 121440 672320 121530 672560
rect 121770 672320 121790 672560
rect 110790 672300 121790 672320
rect 122170 683280 133170 683300
rect 122170 683040 122190 683280
rect 122430 683040 122540 683280
rect 122780 683040 122870 683280
rect 123110 683040 123200 683280
rect 123440 683040 123530 683280
rect 123770 683040 123880 683280
rect 124120 683040 124210 683280
rect 124450 683040 124540 683280
rect 124780 683040 124870 683280
rect 125110 683040 125220 683280
rect 125460 683040 125550 683280
rect 125790 683040 125880 683280
rect 126120 683040 126210 683280
rect 126450 683040 126560 683280
rect 126800 683040 126890 683280
rect 127130 683040 127220 683280
rect 127460 683040 127550 683280
rect 127790 683040 127900 683280
rect 128140 683040 128230 683280
rect 128470 683040 128560 683280
rect 128800 683040 128890 683280
rect 129130 683040 129240 683280
rect 129480 683040 129570 683280
rect 129810 683040 129900 683280
rect 130140 683040 130230 683280
rect 130470 683040 130580 683280
rect 130820 683040 130910 683280
rect 131150 683040 131240 683280
rect 131480 683040 131570 683280
rect 131810 683040 131920 683280
rect 132160 683040 132250 683280
rect 132490 683040 132580 683280
rect 132820 683040 132910 683280
rect 133150 683040 133170 683280
rect 122170 682950 133170 683040
rect 122170 682710 122190 682950
rect 122430 682710 122540 682950
rect 122780 682710 122870 682950
rect 123110 682710 123200 682950
rect 123440 682710 123530 682950
rect 123770 682710 123880 682950
rect 124120 682710 124210 682950
rect 124450 682710 124540 682950
rect 124780 682710 124870 682950
rect 125110 682710 125220 682950
rect 125460 682710 125550 682950
rect 125790 682710 125880 682950
rect 126120 682710 126210 682950
rect 126450 682710 126560 682950
rect 126800 682710 126890 682950
rect 127130 682710 127220 682950
rect 127460 682710 127550 682950
rect 127790 682710 127900 682950
rect 128140 682710 128230 682950
rect 128470 682710 128560 682950
rect 128800 682710 128890 682950
rect 129130 682710 129240 682950
rect 129480 682710 129570 682950
rect 129810 682710 129900 682950
rect 130140 682710 130230 682950
rect 130470 682710 130580 682950
rect 130820 682710 130910 682950
rect 131150 682710 131240 682950
rect 131480 682710 131570 682950
rect 131810 682710 131920 682950
rect 132160 682710 132250 682950
rect 132490 682710 132580 682950
rect 132820 682710 132910 682950
rect 133150 682710 133170 682950
rect 122170 682620 133170 682710
rect 122170 682380 122190 682620
rect 122430 682380 122540 682620
rect 122780 682380 122870 682620
rect 123110 682380 123200 682620
rect 123440 682380 123530 682620
rect 123770 682380 123880 682620
rect 124120 682380 124210 682620
rect 124450 682380 124540 682620
rect 124780 682380 124870 682620
rect 125110 682380 125220 682620
rect 125460 682380 125550 682620
rect 125790 682380 125880 682620
rect 126120 682380 126210 682620
rect 126450 682380 126560 682620
rect 126800 682380 126890 682620
rect 127130 682380 127220 682620
rect 127460 682380 127550 682620
rect 127790 682380 127900 682620
rect 128140 682380 128230 682620
rect 128470 682380 128560 682620
rect 128800 682380 128890 682620
rect 129130 682380 129240 682620
rect 129480 682380 129570 682620
rect 129810 682380 129900 682620
rect 130140 682380 130230 682620
rect 130470 682380 130580 682620
rect 130820 682380 130910 682620
rect 131150 682380 131240 682620
rect 131480 682380 131570 682620
rect 131810 682380 131920 682620
rect 132160 682380 132250 682620
rect 132490 682380 132580 682620
rect 132820 682380 132910 682620
rect 133150 682380 133170 682620
rect 122170 682290 133170 682380
rect 122170 682050 122190 682290
rect 122430 682050 122540 682290
rect 122780 682050 122870 682290
rect 123110 682050 123200 682290
rect 123440 682050 123530 682290
rect 123770 682050 123880 682290
rect 124120 682050 124210 682290
rect 124450 682050 124540 682290
rect 124780 682050 124870 682290
rect 125110 682050 125220 682290
rect 125460 682050 125550 682290
rect 125790 682050 125880 682290
rect 126120 682050 126210 682290
rect 126450 682050 126560 682290
rect 126800 682050 126890 682290
rect 127130 682050 127220 682290
rect 127460 682050 127550 682290
rect 127790 682050 127900 682290
rect 128140 682050 128230 682290
rect 128470 682050 128560 682290
rect 128800 682050 128890 682290
rect 129130 682050 129240 682290
rect 129480 682050 129570 682290
rect 129810 682050 129900 682290
rect 130140 682050 130230 682290
rect 130470 682050 130580 682290
rect 130820 682050 130910 682290
rect 131150 682050 131240 682290
rect 131480 682050 131570 682290
rect 131810 682050 131920 682290
rect 132160 682050 132250 682290
rect 132490 682050 132580 682290
rect 132820 682050 132910 682290
rect 133150 682050 133170 682290
rect 122170 681940 133170 682050
rect 122170 681700 122190 681940
rect 122430 681700 122540 681940
rect 122780 681700 122870 681940
rect 123110 681700 123200 681940
rect 123440 681700 123530 681940
rect 123770 681700 123880 681940
rect 124120 681700 124210 681940
rect 124450 681700 124540 681940
rect 124780 681700 124870 681940
rect 125110 681700 125220 681940
rect 125460 681700 125550 681940
rect 125790 681700 125880 681940
rect 126120 681700 126210 681940
rect 126450 681700 126560 681940
rect 126800 681700 126890 681940
rect 127130 681700 127220 681940
rect 127460 681700 127550 681940
rect 127790 681700 127900 681940
rect 128140 681700 128230 681940
rect 128470 681700 128560 681940
rect 128800 681700 128890 681940
rect 129130 681700 129240 681940
rect 129480 681700 129570 681940
rect 129810 681700 129900 681940
rect 130140 681700 130230 681940
rect 130470 681700 130580 681940
rect 130820 681700 130910 681940
rect 131150 681700 131240 681940
rect 131480 681700 131570 681940
rect 131810 681700 131920 681940
rect 132160 681700 132250 681940
rect 132490 681700 132580 681940
rect 132820 681700 132910 681940
rect 133150 681700 133170 681940
rect 122170 681610 133170 681700
rect 122170 681370 122190 681610
rect 122430 681370 122540 681610
rect 122780 681370 122870 681610
rect 123110 681370 123200 681610
rect 123440 681370 123530 681610
rect 123770 681370 123880 681610
rect 124120 681370 124210 681610
rect 124450 681370 124540 681610
rect 124780 681370 124870 681610
rect 125110 681370 125220 681610
rect 125460 681370 125550 681610
rect 125790 681370 125880 681610
rect 126120 681370 126210 681610
rect 126450 681370 126560 681610
rect 126800 681370 126890 681610
rect 127130 681370 127220 681610
rect 127460 681370 127550 681610
rect 127790 681370 127900 681610
rect 128140 681370 128230 681610
rect 128470 681370 128560 681610
rect 128800 681370 128890 681610
rect 129130 681370 129240 681610
rect 129480 681370 129570 681610
rect 129810 681370 129900 681610
rect 130140 681370 130230 681610
rect 130470 681370 130580 681610
rect 130820 681370 130910 681610
rect 131150 681370 131240 681610
rect 131480 681370 131570 681610
rect 131810 681370 131920 681610
rect 132160 681370 132250 681610
rect 132490 681370 132580 681610
rect 132820 681370 132910 681610
rect 133150 681370 133170 681610
rect 122170 681280 133170 681370
rect 122170 681040 122190 681280
rect 122430 681040 122540 681280
rect 122780 681040 122870 681280
rect 123110 681040 123200 681280
rect 123440 681040 123530 681280
rect 123770 681040 123880 681280
rect 124120 681040 124210 681280
rect 124450 681040 124540 681280
rect 124780 681040 124870 681280
rect 125110 681040 125220 681280
rect 125460 681040 125550 681280
rect 125790 681040 125880 681280
rect 126120 681040 126210 681280
rect 126450 681040 126560 681280
rect 126800 681040 126890 681280
rect 127130 681040 127220 681280
rect 127460 681040 127550 681280
rect 127790 681040 127900 681280
rect 128140 681040 128230 681280
rect 128470 681040 128560 681280
rect 128800 681040 128890 681280
rect 129130 681040 129240 681280
rect 129480 681040 129570 681280
rect 129810 681040 129900 681280
rect 130140 681040 130230 681280
rect 130470 681040 130580 681280
rect 130820 681040 130910 681280
rect 131150 681040 131240 681280
rect 131480 681040 131570 681280
rect 131810 681040 131920 681280
rect 132160 681040 132250 681280
rect 132490 681040 132580 681280
rect 132820 681040 132910 681280
rect 133150 681040 133170 681280
rect 122170 680950 133170 681040
rect 122170 680710 122190 680950
rect 122430 680710 122540 680950
rect 122780 680710 122870 680950
rect 123110 680710 123200 680950
rect 123440 680710 123530 680950
rect 123770 680710 123880 680950
rect 124120 680710 124210 680950
rect 124450 680710 124540 680950
rect 124780 680710 124870 680950
rect 125110 680710 125220 680950
rect 125460 680710 125550 680950
rect 125790 680710 125880 680950
rect 126120 680710 126210 680950
rect 126450 680710 126560 680950
rect 126800 680710 126890 680950
rect 127130 680710 127220 680950
rect 127460 680710 127550 680950
rect 127790 680710 127900 680950
rect 128140 680710 128230 680950
rect 128470 680710 128560 680950
rect 128800 680710 128890 680950
rect 129130 680710 129240 680950
rect 129480 680710 129570 680950
rect 129810 680710 129900 680950
rect 130140 680710 130230 680950
rect 130470 680710 130580 680950
rect 130820 680710 130910 680950
rect 131150 680710 131240 680950
rect 131480 680710 131570 680950
rect 131810 680710 131920 680950
rect 132160 680710 132250 680950
rect 132490 680710 132580 680950
rect 132820 680710 132910 680950
rect 133150 680710 133170 680950
rect 122170 680600 133170 680710
rect 122170 680360 122190 680600
rect 122430 680360 122540 680600
rect 122780 680360 122870 680600
rect 123110 680360 123200 680600
rect 123440 680360 123530 680600
rect 123770 680360 123880 680600
rect 124120 680360 124210 680600
rect 124450 680360 124540 680600
rect 124780 680360 124870 680600
rect 125110 680360 125220 680600
rect 125460 680360 125550 680600
rect 125790 680360 125880 680600
rect 126120 680360 126210 680600
rect 126450 680360 126560 680600
rect 126800 680360 126890 680600
rect 127130 680360 127220 680600
rect 127460 680360 127550 680600
rect 127790 680360 127900 680600
rect 128140 680360 128230 680600
rect 128470 680360 128560 680600
rect 128800 680360 128890 680600
rect 129130 680360 129240 680600
rect 129480 680360 129570 680600
rect 129810 680360 129900 680600
rect 130140 680360 130230 680600
rect 130470 680360 130580 680600
rect 130820 680360 130910 680600
rect 131150 680360 131240 680600
rect 131480 680360 131570 680600
rect 131810 680360 131920 680600
rect 132160 680360 132250 680600
rect 132490 680360 132580 680600
rect 132820 680360 132910 680600
rect 133150 680360 133170 680600
rect 122170 680270 133170 680360
rect 122170 680030 122190 680270
rect 122430 680030 122540 680270
rect 122780 680030 122870 680270
rect 123110 680030 123200 680270
rect 123440 680030 123530 680270
rect 123770 680030 123880 680270
rect 124120 680030 124210 680270
rect 124450 680030 124540 680270
rect 124780 680030 124870 680270
rect 125110 680030 125220 680270
rect 125460 680030 125550 680270
rect 125790 680030 125880 680270
rect 126120 680030 126210 680270
rect 126450 680030 126560 680270
rect 126800 680030 126890 680270
rect 127130 680030 127220 680270
rect 127460 680030 127550 680270
rect 127790 680030 127900 680270
rect 128140 680030 128230 680270
rect 128470 680030 128560 680270
rect 128800 680030 128890 680270
rect 129130 680030 129240 680270
rect 129480 680030 129570 680270
rect 129810 680030 129900 680270
rect 130140 680030 130230 680270
rect 130470 680030 130580 680270
rect 130820 680030 130910 680270
rect 131150 680030 131240 680270
rect 131480 680030 131570 680270
rect 131810 680030 131920 680270
rect 132160 680030 132250 680270
rect 132490 680030 132580 680270
rect 132820 680030 132910 680270
rect 133150 680030 133170 680270
rect 122170 679940 133170 680030
rect 122170 679700 122190 679940
rect 122430 679700 122540 679940
rect 122780 679700 122870 679940
rect 123110 679700 123200 679940
rect 123440 679700 123530 679940
rect 123770 679700 123880 679940
rect 124120 679700 124210 679940
rect 124450 679700 124540 679940
rect 124780 679700 124870 679940
rect 125110 679700 125220 679940
rect 125460 679700 125550 679940
rect 125790 679700 125880 679940
rect 126120 679700 126210 679940
rect 126450 679700 126560 679940
rect 126800 679700 126890 679940
rect 127130 679700 127220 679940
rect 127460 679700 127550 679940
rect 127790 679700 127900 679940
rect 128140 679700 128230 679940
rect 128470 679700 128560 679940
rect 128800 679700 128890 679940
rect 129130 679700 129240 679940
rect 129480 679700 129570 679940
rect 129810 679700 129900 679940
rect 130140 679700 130230 679940
rect 130470 679700 130580 679940
rect 130820 679700 130910 679940
rect 131150 679700 131240 679940
rect 131480 679700 131570 679940
rect 131810 679700 131920 679940
rect 132160 679700 132250 679940
rect 132490 679700 132580 679940
rect 132820 679700 132910 679940
rect 133150 679700 133170 679940
rect 122170 679610 133170 679700
rect 122170 679370 122190 679610
rect 122430 679370 122540 679610
rect 122780 679370 122870 679610
rect 123110 679370 123200 679610
rect 123440 679370 123530 679610
rect 123770 679370 123880 679610
rect 124120 679370 124210 679610
rect 124450 679370 124540 679610
rect 124780 679370 124870 679610
rect 125110 679370 125220 679610
rect 125460 679370 125550 679610
rect 125790 679370 125880 679610
rect 126120 679370 126210 679610
rect 126450 679370 126560 679610
rect 126800 679370 126890 679610
rect 127130 679370 127220 679610
rect 127460 679370 127550 679610
rect 127790 679370 127900 679610
rect 128140 679370 128230 679610
rect 128470 679370 128560 679610
rect 128800 679370 128890 679610
rect 129130 679370 129240 679610
rect 129480 679370 129570 679610
rect 129810 679370 129900 679610
rect 130140 679370 130230 679610
rect 130470 679370 130580 679610
rect 130820 679370 130910 679610
rect 131150 679370 131240 679610
rect 131480 679370 131570 679610
rect 131810 679370 131920 679610
rect 132160 679370 132250 679610
rect 132490 679370 132580 679610
rect 132820 679370 132910 679610
rect 133150 679370 133170 679610
rect 122170 679260 133170 679370
rect 122170 679020 122190 679260
rect 122430 679020 122540 679260
rect 122780 679020 122870 679260
rect 123110 679020 123200 679260
rect 123440 679020 123530 679260
rect 123770 679020 123880 679260
rect 124120 679020 124210 679260
rect 124450 679020 124540 679260
rect 124780 679020 124870 679260
rect 125110 679020 125220 679260
rect 125460 679020 125550 679260
rect 125790 679020 125880 679260
rect 126120 679020 126210 679260
rect 126450 679020 126560 679260
rect 126800 679020 126890 679260
rect 127130 679020 127220 679260
rect 127460 679020 127550 679260
rect 127790 679020 127900 679260
rect 128140 679020 128230 679260
rect 128470 679020 128560 679260
rect 128800 679020 128890 679260
rect 129130 679020 129240 679260
rect 129480 679020 129570 679260
rect 129810 679020 129900 679260
rect 130140 679020 130230 679260
rect 130470 679020 130580 679260
rect 130820 679020 130910 679260
rect 131150 679020 131240 679260
rect 131480 679020 131570 679260
rect 131810 679020 131920 679260
rect 132160 679020 132250 679260
rect 132490 679020 132580 679260
rect 132820 679020 132910 679260
rect 133150 679020 133170 679260
rect 122170 678930 133170 679020
rect 122170 678690 122190 678930
rect 122430 678690 122540 678930
rect 122780 678690 122870 678930
rect 123110 678690 123200 678930
rect 123440 678690 123530 678930
rect 123770 678690 123880 678930
rect 124120 678690 124210 678930
rect 124450 678690 124540 678930
rect 124780 678690 124870 678930
rect 125110 678690 125220 678930
rect 125460 678690 125550 678930
rect 125790 678690 125880 678930
rect 126120 678690 126210 678930
rect 126450 678690 126560 678930
rect 126800 678690 126890 678930
rect 127130 678690 127220 678930
rect 127460 678690 127550 678930
rect 127790 678690 127900 678930
rect 128140 678690 128230 678930
rect 128470 678690 128560 678930
rect 128800 678690 128890 678930
rect 129130 678690 129240 678930
rect 129480 678690 129570 678930
rect 129810 678690 129900 678930
rect 130140 678690 130230 678930
rect 130470 678690 130580 678930
rect 130820 678690 130910 678930
rect 131150 678690 131240 678930
rect 131480 678690 131570 678930
rect 131810 678690 131920 678930
rect 132160 678690 132250 678930
rect 132490 678690 132580 678930
rect 132820 678690 132910 678930
rect 133150 678690 133170 678930
rect 122170 678600 133170 678690
rect 122170 678360 122190 678600
rect 122430 678360 122540 678600
rect 122780 678360 122870 678600
rect 123110 678360 123200 678600
rect 123440 678360 123530 678600
rect 123770 678360 123880 678600
rect 124120 678360 124210 678600
rect 124450 678360 124540 678600
rect 124780 678360 124870 678600
rect 125110 678360 125220 678600
rect 125460 678360 125550 678600
rect 125790 678360 125880 678600
rect 126120 678360 126210 678600
rect 126450 678360 126560 678600
rect 126800 678360 126890 678600
rect 127130 678360 127220 678600
rect 127460 678360 127550 678600
rect 127790 678360 127900 678600
rect 128140 678360 128230 678600
rect 128470 678360 128560 678600
rect 128800 678360 128890 678600
rect 129130 678360 129240 678600
rect 129480 678360 129570 678600
rect 129810 678360 129900 678600
rect 130140 678360 130230 678600
rect 130470 678360 130580 678600
rect 130820 678360 130910 678600
rect 131150 678360 131240 678600
rect 131480 678360 131570 678600
rect 131810 678360 131920 678600
rect 132160 678360 132250 678600
rect 132490 678360 132580 678600
rect 132820 678360 132910 678600
rect 133150 678360 133170 678600
rect 122170 678270 133170 678360
rect 122170 678030 122190 678270
rect 122430 678030 122540 678270
rect 122780 678030 122870 678270
rect 123110 678030 123200 678270
rect 123440 678030 123530 678270
rect 123770 678030 123880 678270
rect 124120 678030 124210 678270
rect 124450 678030 124540 678270
rect 124780 678030 124870 678270
rect 125110 678030 125220 678270
rect 125460 678030 125550 678270
rect 125790 678030 125880 678270
rect 126120 678030 126210 678270
rect 126450 678030 126560 678270
rect 126800 678030 126890 678270
rect 127130 678030 127220 678270
rect 127460 678030 127550 678270
rect 127790 678030 127900 678270
rect 128140 678030 128230 678270
rect 128470 678030 128560 678270
rect 128800 678030 128890 678270
rect 129130 678030 129240 678270
rect 129480 678030 129570 678270
rect 129810 678030 129900 678270
rect 130140 678030 130230 678270
rect 130470 678030 130580 678270
rect 130820 678030 130910 678270
rect 131150 678030 131240 678270
rect 131480 678030 131570 678270
rect 131810 678030 131920 678270
rect 132160 678030 132250 678270
rect 132490 678030 132580 678270
rect 132820 678030 132910 678270
rect 133150 678030 133170 678270
rect 122170 677920 133170 678030
rect 122170 677680 122190 677920
rect 122430 677680 122540 677920
rect 122780 677680 122870 677920
rect 123110 677680 123200 677920
rect 123440 677680 123530 677920
rect 123770 677680 123880 677920
rect 124120 677680 124210 677920
rect 124450 677680 124540 677920
rect 124780 677680 124870 677920
rect 125110 677680 125220 677920
rect 125460 677680 125550 677920
rect 125790 677680 125880 677920
rect 126120 677680 126210 677920
rect 126450 677680 126560 677920
rect 126800 677680 126890 677920
rect 127130 677680 127220 677920
rect 127460 677680 127550 677920
rect 127790 677680 127900 677920
rect 128140 677680 128230 677920
rect 128470 677680 128560 677920
rect 128800 677680 128890 677920
rect 129130 677680 129240 677920
rect 129480 677680 129570 677920
rect 129810 677680 129900 677920
rect 130140 677680 130230 677920
rect 130470 677680 130580 677920
rect 130820 677680 130910 677920
rect 131150 677680 131240 677920
rect 131480 677680 131570 677920
rect 131810 677680 131920 677920
rect 132160 677680 132250 677920
rect 132490 677680 132580 677920
rect 132820 677680 132910 677920
rect 133150 677680 133170 677920
rect 122170 677590 133170 677680
rect 122170 677350 122190 677590
rect 122430 677350 122540 677590
rect 122780 677350 122870 677590
rect 123110 677350 123200 677590
rect 123440 677350 123530 677590
rect 123770 677350 123880 677590
rect 124120 677350 124210 677590
rect 124450 677350 124540 677590
rect 124780 677350 124870 677590
rect 125110 677350 125220 677590
rect 125460 677350 125550 677590
rect 125790 677350 125880 677590
rect 126120 677350 126210 677590
rect 126450 677350 126560 677590
rect 126800 677350 126890 677590
rect 127130 677350 127220 677590
rect 127460 677350 127550 677590
rect 127790 677350 127900 677590
rect 128140 677350 128230 677590
rect 128470 677350 128560 677590
rect 128800 677350 128890 677590
rect 129130 677350 129240 677590
rect 129480 677350 129570 677590
rect 129810 677350 129900 677590
rect 130140 677350 130230 677590
rect 130470 677350 130580 677590
rect 130820 677350 130910 677590
rect 131150 677350 131240 677590
rect 131480 677350 131570 677590
rect 131810 677350 131920 677590
rect 132160 677350 132250 677590
rect 132490 677350 132580 677590
rect 132820 677350 132910 677590
rect 133150 677350 133170 677590
rect 122170 677260 133170 677350
rect 122170 677020 122190 677260
rect 122430 677020 122540 677260
rect 122780 677020 122870 677260
rect 123110 677020 123200 677260
rect 123440 677020 123530 677260
rect 123770 677020 123880 677260
rect 124120 677020 124210 677260
rect 124450 677020 124540 677260
rect 124780 677020 124870 677260
rect 125110 677020 125220 677260
rect 125460 677020 125550 677260
rect 125790 677020 125880 677260
rect 126120 677020 126210 677260
rect 126450 677020 126560 677260
rect 126800 677020 126890 677260
rect 127130 677020 127220 677260
rect 127460 677020 127550 677260
rect 127790 677020 127900 677260
rect 128140 677020 128230 677260
rect 128470 677020 128560 677260
rect 128800 677020 128890 677260
rect 129130 677020 129240 677260
rect 129480 677020 129570 677260
rect 129810 677020 129900 677260
rect 130140 677020 130230 677260
rect 130470 677020 130580 677260
rect 130820 677020 130910 677260
rect 131150 677020 131240 677260
rect 131480 677020 131570 677260
rect 131810 677020 131920 677260
rect 132160 677020 132250 677260
rect 132490 677020 132580 677260
rect 132820 677020 132910 677260
rect 133150 677020 133170 677260
rect 122170 676930 133170 677020
rect 122170 676690 122190 676930
rect 122430 676690 122540 676930
rect 122780 676690 122870 676930
rect 123110 676690 123200 676930
rect 123440 676690 123530 676930
rect 123770 676690 123880 676930
rect 124120 676690 124210 676930
rect 124450 676690 124540 676930
rect 124780 676690 124870 676930
rect 125110 676690 125220 676930
rect 125460 676690 125550 676930
rect 125790 676690 125880 676930
rect 126120 676690 126210 676930
rect 126450 676690 126560 676930
rect 126800 676690 126890 676930
rect 127130 676690 127220 676930
rect 127460 676690 127550 676930
rect 127790 676690 127900 676930
rect 128140 676690 128230 676930
rect 128470 676690 128560 676930
rect 128800 676690 128890 676930
rect 129130 676690 129240 676930
rect 129480 676690 129570 676930
rect 129810 676690 129900 676930
rect 130140 676690 130230 676930
rect 130470 676690 130580 676930
rect 130820 676690 130910 676930
rect 131150 676690 131240 676930
rect 131480 676690 131570 676930
rect 131810 676690 131920 676930
rect 132160 676690 132250 676930
rect 132490 676690 132580 676930
rect 132820 676690 132910 676930
rect 133150 676690 133170 676930
rect 122170 676580 133170 676690
rect 122170 676340 122190 676580
rect 122430 676340 122540 676580
rect 122780 676340 122870 676580
rect 123110 676340 123200 676580
rect 123440 676340 123530 676580
rect 123770 676340 123880 676580
rect 124120 676340 124210 676580
rect 124450 676340 124540 676580
rect 124780 676340 124870 676580
rect 125110 676340 125220 676580
rect 125460 676340 125550 676580
rect 125790 676340 125880 676580
rect 126120 676340 126210 676580
rect 126450 676340 126560 676580
rect 126800 676340 126890 676580
rect 127130 676340 127220 676580
rect 127460 676340 127550 676580
rect 127790 676340 127900 676580
rect 128140 676340 128230 676580
rect 128470 676340 128560 676580
rect 128800 676340 128890 676580
rect 129130 676340 129240 676580
rect 129480 676340 129570 676580
rect 129810 676340 129900 676580
rect 130140 676340 130230 676580
rect 130470 676340 130580 676580
rect 130820 676340 130910 676580
rect 131150 676340 131240 676580
rect 131480 676340 131570 676580
rect 131810 676340 131920 676580
rect 132160 676340 132250 676580
rect 132490 676340 132580 676580
rect 132820 676340 132910 676580
rect 133150 676340 133170 676580
rect 122170 676250 133170 676340
rect 122170 676010 122190 676250
rect 122430 676010 122540 676250
rect 122780 676010 122870 676250
rect 123110 676010 123200 676250
rect 123440 676010 123530 676250
rect 123770 676010 123880 676250
rect 124120 676010 124210 676250
rect 124450 676010 124540 676250
rect 124780 676010 124870 676250
rect 125110 676010 125220 676250
rect 125460 676010 125550 676250
rect 125790 676010 125880 676250
rect 126120 676010 126210 676250
rect 126450 676010 126560 676250
rect 126800 676010 126890 676250
rect 127130 676010 127220 676250
rect 127460 676010 127550 676250
rect 127790 676010 127900 676250
rect 128140 676010 128230 676250
rect 128470 676010 128560 676250
rect 128800 676010 128890 676250
rect 129130 676010 129240 676250
rect 129480 676010 129570 676250
rect 129810 676010 129900 676250
rect 130140 676010 130230 676250
rect 130470 676010 130580 676250
rect 130820 676010 130910 676250
rect 131150 676010 131240 676250
rect 131480 676010 131570 676250
rect 131810 676010 131920 676250
rect 132160 676010 132250 676250
rect 132490 676010 132580 676250
rect 132820 676010 132910 676250
rect 133150 676010 133170 676250
rect 122170 675920 133170 676010
rect 122170 675680 122190 675920
rect 122430 675680 122540 675920
rect 122780 675680 122870 675920
rect 123110 675680 123200 675920
rect 123440 675680 123530 675920
rect 123770 675680 123880 675920
rect 124120 675680 124210 675920
rect 124450 675680 124540 675920
rect 124780 675680 124870 675920
rect 125110 675680 125220 675920
rect 125460 675680 125550 675920
rect 125790 675680 125880 675920
rect 126120 675680 126210 675920
rect 126450 675680 126560 675920
rect 126800 675680 126890 675920
rect 127130 675680 127220 675920
rect 127460 675680 127550 675920
rect 127790 675680 127900 675920
rect 128140 675680 128230 675920
rect 128470 675680 128560 675920
rect 128800 675680 128890 675920
rect 129130 675680 129240 675920
rect 129480 675680 129570 675920
rect 129810 675680 129900 675920
rect 130140 675680 130230 675920
rect 130470 675680 130580 675920
rect 130820 675680 130910 675920
rect 131150 675680 131240 675920
rect 131480 675680 131570 675920
rect 131810 675680 131920 675920
rect 132160 675680 132250 675920
rect 132490 675680 132580 675920
rect 132820 675680 132910 675920
rect 133150 675680 133170 675920
rect 122170 675590 133170 675680
rect 122170 675350 122190 675590
rect 122430 675350 122540 675590
rect 122780 675350 122870 675590
rect 123110 675350 123200 675590
rect 123440 675350 123530 675590
rect 123770 675350 123880 675590
rect 124120 675350 124210 675590
rect 124450 675350 124540 675590
rect 124780 675350 124870 675590
rect 125110 675350 125220 675590
rect 125460 675350 125550 675590
rect 125790 675350 125880 675590
rect 126120 675350 126210 675590
rect 126450 675350 126560 675590
rect 126800 675350 126890 675590
rect 127130 675350 127220 675590
rect 127460 675350 127550 675590
rect 127790 675350 127900 675590
rect 128140 675350 128230 675590
rect 128470 675350 128560 675590
rect 128800 675350 128890 675590
rect 129130 675350 129240 675590
rect 129480 675350 129570 675590
rect 129810 675350 129900 675590
rect 130140 675350 130230 675590
rect 130470 675350 130580 675590
rect 130820 675350 130910 675590
rect 131150 675350 131240 675590
rect 131480 675350 131570 675590
rect 131810 675350 131920 675590
rect 132160 675350 132250 675590
rect 132490 675350 132580 675590
rect 132820 675350 132910 675590
rect 133150 675350 133170 675590
rect 122170 675240 133170 675350
rect 122170 675000 122190 675240
rect 122430 675000 122540 675240
rect 122780 675000 122870 675240
rect 123110 675000 123200 675240
rect 123440 675000 123530 675240
rect 123770 675000 123880 675240
rect 124120 675000 124210 675240
rect 124450 675000 124540 675240
rect 124780 675000 124870 675240
rect 125110 675000 125220 675240
rect 125460 675000 125550 675240
rect 125790 675000 125880 675240
rect 126120 675000 126210 675240
rect 126450 675000 126560 675240
rect 126800 675000 126890 675240
rect 127130 675000 127220 675240
rect 127460 675000 127550 675240
rect 127790 675000 127900 675240
rect 128140 675000 128230 675240
rect 128470 675000 128560 675240
rect 128800 675000 128890 675240
rect 129130 675000 129240 675240
rect 129480 675000 129570 675240
rect 129810 675000 129900 675240
rect 130140 675000 130230 675240
rect 130470 675000 130580 675240
rect 130820 675000 130910 675240
rect 131150 675000 131240 675240
rect 131480 675000 131570 675240
rect 131810 675000 131920 675240
rect 132160 675000 132250 675240
rect 132490 675000 132580 675240
rect 132820 675000 132910 675240
rect 133150 675000 133170 675240
rect 122170 674910 133170 675000
rect 122170 674670 122190 674910
rect 122430 674670 122540 674910
rect 122780 674670 122870 674910
rect 123110 674670 123200 674910
rect 123440 674670 123530 674910
rect 123770 674670 123880 674910
rect 124120 674670 124210 674910
rect 124450 674670 124540 674910
rect 124780 674670 124870 674910
rect 125110 674670 125220 674910
rect 125460 674670 125550 674910
rect 125790 674670 125880 674910
rect 126120 674670 126210 674910
rect 126450 674670 126560 674910
rect 126800 674670 126890 674910
rect 127130 674670 127220 674910
rect 127460 674670 127550 674910
rect 127790 674670 127900 674910
rect 128140 674670 128230 674910
rect 128470 674670 128560 674910
rect 128800 674670 128890 674910
rect 129130 674670 129240 674910
rect 129480 674670 129570 674910
rect 129810 674670 129900 674910
rect 130140 674670 130230 674910
rect 130470 674670 130580 674910
rect 130820 674670 130910 674910
rect 131150 674670 131240 674910
rect 131480 674670 131570 674910
rect 131810 674670 131920 674910
rect 132160 674670 132250 674910
rect 132490 674670 132580 674910
rect 132820 674670 132910 674910
rect 133150 674670 133170 674910
rect 122170 674580 133170 674670
rect 122170 674340 122190 674580
rect 122430 674340 122540 674580
rect 122780 674340 122870 674580
rect 123110 674340 123200 674580
rect 123440 674340 123530 674580
rect 123770 674340 123880 674580
rect 124120 674340 124210 674580
rect 124450 674340 124540 674580
rect 124780 674340 124870 674580
rect 125110 674340 125220 674580
rect 125460 674340 125550 674580
rect 125790 674340 125880 674580
rect 126120 674340 126210 674580
rect 126450 674340 126560 674580
rect 126800 674340 126890 674580
rect 127130 674340 127220 674580
rect 127460 674340 127550 674580
rect 127790 674340 127900 674580
rect 128140 674340 128230 674580
rect 128470 674340 128560 674580
rect 128800 674340 128890 674580
rect 129130 674340 129240 674580
rect 129480 674340 129570 674580
rect 129810 674340 129900 674580
rect 130140 674340 130230 674580
rect 130470 674340 130580 674580
rect 130820 674340 130910 674580
rect 131150 674340 131240 674580
rect 131480 674340 131570 674580
rect 131810 674340 131920 674580
rect 132160 674340 132250 674580
rect 132490 674340 132580 674580
rect 132820 674340 132910 674580
rect 133150 674340 133170 674580
rect 122170 674250 133170 674340
rect 122170 674010 122190 674250
rect 122430 674010 122540 674250
rect 122780 674010 122870 674250
rect 123110 674010 123200 674250
rect 123440 674010 123530 674250
rect 123770 674010 123880 674250
rect 124120 674010 124210 674250
rect 124450 674010 124540 674250
rect 124780 674010 124870 674250
rect 125110 674010 125220 674250
rect 125460 674010 125550 674250
rect 125790 674010 125880 674250
rect 126120 674010 126210 674250
rect 126450 674010 126560 674250
rect 126800 674010 126890 674250
rect 127130 674010 127220 674250
rect 127460 674010 127550 674250
rect 127790 674010 127900 674250
rect 128140 674010 128230 674250
rect 128470 674010 128560 674250
rect 128800 674010 128890 674250
rect 129130 674010 129240 674250
rect 129480 674010 129570 674250
rect 129810 674010 129900 674250
rect 130140 674010 130230 674250
rect 130470 674010 130580 674250
rect 130820 674010 130910 674250
rect 131150 674010 131240 674250
rect 131480 674010 131570 674250
rect 131810 674010 131920 674250
rect 132160 674010 132250 674250
rect 132490 674010 132580 674250
rect 132820 674010 132910 674250
rect 133150 674010 133170 674250
rect 122170 673900 133170 674010
rect 122170 673660 122190 673900
rect 122430 673660 122540 673900
rect 122780 673660 122870 673900
rect 123110 673660 123200 673900
rect 123440 673660 123530 673900
rect 123770 673660 123880 673900
rect 124120 673660 124210 673900
rect 124450 673660 124540 673900
rect 124780 673660 124870 673900
rect 125110 673660 125220 673900
rect 125460 673660 125550 673900
rect 125790 673660 125880 673900
rect 126120 673660 126210 673900
rect 126450 673660 126560 673900
rect 126800 673660 126890 673900
rect 127130 673660 127220 673900
rect 127460 673660 127550 673900
rect 127790 673660 127900 673900
rect 128140 673660 128230 673900
rect 128470 673660 128560 673900
rect 128800 673660 128890 673900
rect 129130 673660 129240 673900
rect 129480 673660 129570 673900
rect 129810 673660 129900 673900
rect 130140 673660 130230 673900
rect 130470 673660 130580 673900
rect 130820 673660 130910 673900
rect 131150 673660 131240 673900
rect 131480 673660 131570 673900
rect 131810 673660 131920 673900
rect 132160 673660 132250 673900
rect 132490 673660 132580 673900
rect 132820 673660 132910 673900
rect 133150 673660 133170 673900
rect 122170 673570 133170 673660
rect 122170 673330 122190 673570
rect 122430 673330 122540 673570
rect 122780 673330 122870 673570
rect 123110 673330 123200 673570
rect 123440 673330 123530 673570
rect 123770 673330 123880 673570
rect 124120 673330 124210 673570
rect 124450 673330 124540 673570
rect 124780 673330 124870 673570
rect 125110 673330 125220 673570
rect 125460 673330 125550 673570
rect 125790 673330 125880 673570
rect 126120 673330 126210 673570
rect 126450 673330 126560 673570
rect 126800 673330 126890 673570
rect 127130 673330 127220 673570
rect 127460 673330 127550 673570
rect 127790 673330 127900 673570
rect 128140 673330 128230 673570
rect 128470 673330 128560 673570
rect 128800 673330 128890 673570
rect 129130 673330 129240 673570
rect 129480 673330 129570 673570
rect 129810 673330 129900 673570
rect 130140 673330 130230 673570
rect 130470 673330 130580 673570
rect 130820 673330 130910 673570
rect 131150 673330 131240 673570
rect 131480 673330 131570 673570
rect 131810 673330 131920 673570
rect 132160 673330 132250 673570
rect 132490 673330 132580 673570
rect 132820 673330 132910 673570
rect 133150 673330 133170 673570
rect 122170 673240 133170 673330
rect 122170 673000 122190 673240
rect 122430 673000 122540 673240
rect 122780 673000 122870 673240
rect 123110 673000 123200 673240
rect 123440 673000 123530 673240
rect 123770 673000 123880 673240
rect 124120 673000 124210 673240
rect 124450 673000 124540 673240
rect 124780 673000 124870 673240
rect 125110 673000 125220 673240
rect 125460 673000 125550 673240
rect 125790 673000 125880 673240
rect 126120 673000 126210 673240
rect 126450 673000 126560 673240
rect 126800 673000 126890 673240
rect 127130 673000 127220 673240
rect 127460 673000 127550 673240
rect 127790 673000 127900 673240
rect 128140 673000 128230 673240
rect 128470 673000 128560 673240
rect 128800 673000 128890 673240
rect 129130 673000 129240 673240
rect 129480 673000 129570 673240
rect 129810 673000 129900 673240
rect 130140 673000 130230 673240
rect 130470 673000 130580 673240
rect 130820 673000 130910 673240
rect 131150 673000 131240 673240
rect 131480 673000 131570 673240
rect 131810 673000 131920 673240
rect 132160 673000 132250 673240
rect 132490 673000 132580 673240
rect 132820 673000 132910 673240
rect 133150 673000 133170 673240
rect 122170 672910 133170 673000
rect 122170 672670 122190 672910
rect 122430 672670 122540 672910
rect 122780 672670 122870 672910
rect 123110 672670 123200 672910
rect 123440 672670 123530 672910
rect 123770 672670 123880 672910
rect 124120 672670 124210 672910
rect 124450 672670 124540 672910
rect 124780 672670 124870 672910
rect 125110 672670 125220 672910
rect 125460 672670 125550 672910
rect 125790 672670 125880 672910
rect 126120 672670 126210 672910
rect 126450 672670 126560 672910
rect 126800 672670 126890 672910
rect 127130 672670 127220 672910
rect 127460 672670 127550 672910
rect 127790 672670 127900 672910
rect 128140 672670 128230 672910
rect 128470 672670 128560 672910
rect 128800 672670 128890 672910
rect 129130 672670 129240 672910
rect 129480 672670 129570 672910
rect 129810 672670 129900 672910
rect 130140 672670 130230 672910
rect 130470 672670 130580 672910
rect 130820 672670 130910 672910
rect 131150 672670 131240 672910
rect 131480 672670 131570 672910
rect 131810 672670 131920 672910
rect 132160 672670 132250 672910
rect 132490 672670 132580 672910
rect 132820 672670 132910 672910
rect 133150 672670 133170 672910
rect 122170 672560 133170 672670
rect 122170 672320 122190 672560
rect 122430 672320 122540 672560
rect 122780 672320 122870 672560
rect 123110 672320 123200 672560
rect 123440 672320 123530 672560
rect 123770 672320 123880 672560
rect 124120 672320 124210 672560
rect 124450 672320 124540 672560
rect 124780 672320 124870 672560
rect 125110 672320 125220 672560
rect 125460 672320 125550 672560
rect 125790 672320 125880 672560
rect 126120 672320 126210 672560
rect 126450 672320 126560 672560
rect 126800 672320 126890 672560
rect 127130 672320 127220 672560
rect 127460 672320 127550 672560
rect 127790 672320 127900 672560
rect 128140 672320 128230 672560
rect 128470 672320 128560 672560
rect 128800 672320 128890 672560
rect 129130 672320 129240 672560
rect 129480 672320 129570 672560
rect 129810 672320 129900 672560
rect 130140 672320 130230 672560
rect 130470 672320 130580 672560
rect 130820 672320 130910 672560
rect 131150 672320 131240 672560
rect 131480 672320 131570 672560
rect 131810 672320 131920 672560
rect 132160 672320 132250 672560
rect 132490 672320 132580 672560
rect 132820 672320 132910 672560
rect 133150 672320 133170 672560
rect 122170 672300 133170 672320
rect 133550 683280 144550 683300
rect 133550 683040 133570 683280
rect 133810 683040 133920 683280
rect 134160 683040 134250 683280
rect 134490 683040 134580 683280
rect 134820 683040 134910 683280
rect 135150 683040 135260 683280
rect 135500 683040 135590 683280
rect 135830 683040 135920 683280
rect 136160 683040 136250 683280
rect 136490 683040 136600 683280
rect 136840 683040 136930 683280
rect 137170 683040 137260 683280
rect 137500 683040 137590 683280
rect 137830 683040 137940 683280
rect 138180 683040 138270 683280
rect 138510 683040 138600 683280
rect 138840 683040 138930 683280
rect 139170 683040 139280 683280
rect 139520 683040 139610 683280
rect 139850 683040 139940 683280
rect 140180 683040 140270 683280
rect 140510 683040 140620 683280
rect 140860 683040 140950 683280
rect 141190 683040 141280 683280
rect 141520 683040 141610 683280
rect 141850 683040 141960 683280
rect 142200 683040 142290 683280
rect 142530 683040 142620 683280
rect 142860 683040 142950 683280
rect 143190 683040 143300 683280
rect 143540 683040 143630 683280
rect 143870 683040 143960 683280
rect 144200 683040 144290 683280
rect 144530 683040 144550 683280
rect 133550 682950 144550 683040
rect 133550 682710 133570 682950
rect 133810 682710 133920 682950
rect 134160 682710 134250 682950
rect 134490 682710 134580 682950
rect 134820 682710 134910 682950
rect 135150 682710 135260 682950
rect 135500 682710 135590 682950
rect 135830 682710 135920 682950
rect 136160 682710 136250 682950
rect 136490 682710 136600 682950
rect 136840 682710 136930 682950
rect 137170 682710 137260 682950
rect 137500 682710 137590 682950
rect 137830 682710 137940 682950
rect 138180 682710 138270 682950
rect 138510 682710 138600 682950
rect 138840 682710 138930 682950
rect 139170 682710 139280 682950
rect 139520 682710 139610 682950
rect 139850 682710 139940 682950
rect 140180 682710 140270 682950
rect 140510 682710 140620 682950
rect 140860 682710 140950 682950
rect 141190 682710 141280 682950
rect 141520 682710 141610 682950
rect 141850 682710 141960 682950
rect 142200 682710 142290 682950
rect 142530 682710 142620 682950
rect 142860 682710 142950 682950
rect 143190 682710 143300 682950
rect 143540 682710 143630 682950
rect 143870 682710 143960 682950
rect 144200 682710 144290 682950
rect 144530 682710 144550 682950
rect 133550 682620 144550 682710
rect 133550 682380 133570 682620
rect 133810 682380 133920 682620
rect 134160 682380 134250 682620
rect 134490 682380 134580 682620
rect 134820 682380 134910 682620
rect 135150 682380 135260 682620
rect 135500 682380 135590 682620
rect 135830 682380 135920 682620
rect 136160 682380 136250 682620
rect 136490 682380 136600 682620
rect 136840 682380 136930 682620
rect 137170 682380 137260 682620
rect 137500 682380 137590 682620
rect 137830 682380 137940 682620
rect 138180 682380 138270 682620
rect 138510 682380 138600 682620
rect 138840 682380 138930 682620
rect 139170 682380 139280 682620
rect 139520 682380 139610 682620
rect 139850 682380 139940 682620
rect 140180 682380 140270 682620
rect 140510 682380 140620 682620
rect 140860 682380 140950 682620
rect 141190 682380 141280 682620
rect 141520 682380 141610 682620
rect 141850 682380 141960 682620
rect 142200 682380 142290 682620
rect 142530 682380 142620 682620
rect 142860 682380 142950 682620
rect 143190 682380 143300 682620
rect 143540 682380 143630 682620
rect 143870 682380 143960 682620
rect 144200 682380 144290 682620
rect 144530 682380 144550 682620
rect 133550 682290 144550 682380
rect 133550 682050 133570 682290
rect 133810 682050 133920 682290
rect 134160 682050 134250 682290
rect 134490 682050 134580 682290
rect 134820 682050 134910 682290
rect 135150 682050 135260 682290
rect 135500 682050 135590 682290
rect 135830 682050 135920 682290
rect 136160 682050 136250 682290
rect 136490 682050 136600 682290
rect 136840 682050 136930 682290
rect 137170 682050 137260 682290
rect 137500 682050 137590 682290
rect 137830 682050 137940 682290
rect 138180 682050 138270 682290
rect 138510 682050 138600 682290
rect 138840 682050 138930 682290
rect 139170 682050 139280 682290
rect 139520 682050 139610 682290
rect 139850 682050 139940 682290
rect 140180 682050 140270 682290
rect 140510 682050 140620 682290
rect 140860 682050 140950 682290
rect 141190 682050 141280 682290
rect 141520 682050 141610 682290
rect 141850 682050 141960 682290
rect 142200 682050 142290 682290
rect 142530 682050 142620 682290
rect 142860 682050 142950 682290
rect 143190 682050 143300 682290
rect 143540 682050 143630 682290
rect 143870 682050 143960 682290
rect 144200 682050 144290 682290
rect 144530 682050 144550 682290
rect 133550 681940 144550 682050
rect 133550 681700 133570 681940
rect 133810 681700 133920 681940
rect 134160 681700 134250 681940
rect 134490 681700 134580 681940
rect 134820 681700 134910 681940
rect 135150 681700 135260 681940
rect 135500 681700 135590 681940
rect 135830 681700 135920 681940
rect 136160 681700 136250 681940
rect 136490 681700 136600 681940
rect 136840 681700 136930 681940
rect 137170 681700 137260 681940
rect 137500 681700 137590 681940
rect 137830 681700 137940 681940
rect 138180 681700 138270 681940
rect 138510 681700 138600 681940
rect 138840 681700 138930 681940
rect 139170 681700 139280 681940
rect 139520 681700 139610 681940
rect 139850 681700 139940 681940
rect 140180 681700 140270 681940
rect 140510 681700 140620 681940
rect 140860 681700 140950 681940
rect 141190 681700 141280 681940
rect 141520 681700 141610 681940
rect 141850 681700 141960 681940
rect 142200 681700 142290 681940
rect 142530 681700 142620 681940
rect 142860 681700 142950 681940
rect 143190 681700 143300 681940
rect 143540 681700 143630 681940
rect 143870 681700 143960 681940
rect 144200 681700 144290 681940
rect 144530 681700 144550 681940
rect 133550 681610 144550 681700
rect 133550 681370 133570 681610
rect 133810 681370 133920 681610
rect 134160 681370 134250 681610
rect 134490 681370 134580 681610
rect 134820 681370 134910 681610
rect 135150 681370 135260 681610
rect 135500 681370 135590 681610
rect 135830 681370 135920 681610
rect 136160 681370 136250 681610
rect 136490 681370 136600 681610
rect 136840 681370 136930 681610
rect 137170 681370 137260 681610
rect 137500 681370 137590 681610
rect 137830 681370 137940 681610
rect 138180 681370 138270 681610
rect 138510 681370 138600 681610
rect 138840 681370 138930 681610
rect 139170 681370 139280 681610
rect 139520 681370 139610 681610
rect 139850 681370 139940 681610
rect 140180 681370 140270 681610
rect 140510 681370 140620 681610
rect 140860 681370 140950 681610
rect 141190 681370 141280 681610
rect 141520 681370 141610 681610
rect 141850 681370 141960 681610
rect 142200 681370 142290 681610
rect 142530 681370 142620 681610
rect 142860 681370 142950 681610
rect 143190 681370 143300 681610
rect 143540 681370 143630 681610
rect 143870 681370 143960 681610
rect 144200 681370 144290 681610
rect 144530 681370 144550 681610
rect 133550 681280 144550 681370
rect 133550 681040 133570 681280
rect 133810 681040 133920 681280
rect 134160 681040 134250 681280
rect 134490 681040 134580 681280
rect 134820 681040 134910 681280
rect 135150 681040 135260 681280
rect 135500 681040 135590 681280
rect 135830 681040 135920 681280
rect 136160 681040 136250 681280
rect 136490 681040 136600 681280
rect 136840 681040 136930 681280
rect 137170 681040 137260 681280
rect 137500 681040 137590 681280
rect 137830 681040 137940 681280
rect 138180 681040 138270 681280
rect 138510 681040 138600 681280
rect 138840 681040 138930 681280
rect 139170 681040 139280 681280
rect 139520 681040 139610 681280
rect 139850 681040 139940 681280
rect 140180 681040 140270 681280
rect 140510 681040 140620 681280
rect 140860 681040 140950 681280
rect 141190 681040 141280 681280
rect 141520 681040 141610 681280
rect 141850 681040 141960 681280
rect 142200 681040 142290 681280
rect 142530 681040 142620 681280
rect 142860 681040 142950 681280
rect 143190 681040 143300 681280
rect 143540 681040 143630 681280
rect 143870 681040 143960 681280
rect 144200 681040 144290 681280
rect 144530 681040 144550 681280
rect 133550 680950 144550 681040
rect 133550 680710 133570 680950
rect 133810 680710 133920 680950
rect 134160 680710 134250 680950
rect 134490 680710 134580 680950
rect 134820 680710 134910 680950
rect 135150 680710 135260 680950
rect 135500 680710 135590 680950
rect 135830 680710 135920 680950
rect 136160 680710 136250 680950
rect 136490 680710 136600 680950
rect 136840 680710 136930 680950
rect 137170 680710 137260 680950
rect 137500 680710 137590 680950
rect 137830 680710 137940 680950
rect 138180 680710 138270 680950
rect 138510 680710 138600 680950
rect 138840 680710 138930 680950
rect 139170 680710 139280 680950
rect 139520 680710 139610 680950
rect 139850 680710 139940 680950
rect 140180 680710 140270 680950
rect 140510 680710 140620 680950
rect 140860 680710 140950 680950
rect 141190 680710 141280 680950
rect 141520 680710 141610 680950
rect 141850 680710 141960 680950
rect 142200 680710 142290 680950
rect 142530 680710 142620 680950
rect 142860 680710 142950 680950
rect 143190 680710 143300 680950
rect 143540 680710 143630 680950
rect 143870 680710 143960 680950
rect 144200 680710 144290 680950
rect 144530 680710 144550 680950
rect 133550 680600 144550 680710
rect 133550 680360 133570 680600
rect 133810 680360 133920 680600
rect 134160 680360 134250 680600
rect 134490 680360 134580 680600
rect 134820 680360 134910 680600
rect 135150 680360 135260 680600
rect 135500 680360 135590 680600
rect 135830 680360 135920 680600
rect 136160 680360 136250 680600
rect 136490 680360 136600 680600
rect 136840 680360 136930 680600
rect 137170 680360 137260 680600
rect 137500 680360 137590 680600
rect 137830 680360 137940 680600
rect 138180 680360 138270 680600
rect 138510 680360 138600 680600
rect 138840 680360 138930 680600
rect 139170 680360 139280 680600
rect 139520 680360 139610 680600
rect 139850 680360 139940 680600
rect 140180 680360 140270 680600
rect 140510 680360 140620 680600
rect 140860 680360 140950 680600
rect 141190 680360 141280 680600
rect 141520 680360 141610 680600
rect 141850 680360 141960 680600
rect 142200 680360 142290 680600
rect 142530 680360 142620 680600
rect 142860 680360 142950 680600
rect 143190 680360 143300 680600
rect 143540 680360 143630 680600
rect 143870 680360 143960 680600
rect 144200 680360 144290 680600
rect 144530 680360 144550 680600
rect 133550 680270 144550 680360
rect 133550 680030 133570 680270
rect 133810 680030 133920 680270
rect 134160 680030 134250 680270
rect 134490 680030 134580 680270
rect 134820 680030 134910 680270
rect 135150 680030 135260 680270
rect 135500 680030 135590 680270
rect 135830 680030 135920 680270
rect 136160 680030 136250 680270
rect 136490 680030 136600 680270
rect 136840 680030 136930 680270
rect 137170 680030 137260 680270
rect 137500 680030 137590 680270
rect 137830 680030 137940 680270
rect 138180 680030 138270 680270
rect 138510 680030 138600 680270
rect 138840 680030 138930 680270
rect 139170 680030 139280 680270
rect 139520 680030 139610 680270
rect 139850 680030 139940 680270
rect 140180 680030 140270 680270
rect 140510 680030 140620 680270
rect 140860 680030 140950 680270
rect 141190 680030 141280 680270
rect 141520 680030 141610 680270
rect 141850 680030 141960 680270
rect 142200 680030 142290 680270
rect 142530 680030 142620 680270
rect 142860 680030 142950 680270
rect 143190 680030 143300 680270
rect 143540 680030 143630 680270
rect 143870 680030 143960 680270
rect 144200 680030 144290 680270
rect 144530 680030 144550 680270
rect 133550 679940 144550 680030
rect 133550 679700 133570 679940
rect 133810 679700 133920 679940
rect 134160 679700 134250 679940
rect 134490 679700 134580 679940
rect 134820 679700 134910 679940
rect 135150 679700 135260 679940
rect 135500 679700 135590 679940
rect 135830 679700 135920 679940
rect 136160 679700 136250 679940
rect 136490 679700 136600 679940
rect 136840 679700 136930 679940
rect 137170 679700 137260 679940
rect 137500 679700 137590 679940
rect 137830 679700 137940 679940
rect 138180 679700 138270 679940
rect 138510 679700 138600 679940
rect 138840 679700 138930 679940
rect 139170 679700 139280 679940
rect 139520 679700 139610 679940
rect 139850 679700 139940 679940
rect 140180 679700 140270 679940
rect 140510 679700 140620 679940
rect 140860 679700 140950 679940
rect 141190 679700 141280 679940
rect 141520 679700 141610 679940
rect 141850 679700 141960 679940
rect 142200 679700 142290 679940
rect 142530 679700 142620 679940
rect 142860 679700 142950 679940
rect 143190 679700 143300 679940
rect 143540 679700 143630 679940
rect 143870 679700 143960 679940
rect 144200 679700 144290 679940
rect 144530 679700 144550 679940
rect 133550 679610 144550 679700
rect 133550 679370 133570 679610
rect 133810 679370 133920 679610
rect 134160 679370 134250 679610
rect 134490 679370 134580 679610
rect 134820 679370 134910 679610
rect 135150 679370 135260 679610
rect 135500 679370 135590 679610
rect 135830 679370 135920 679610
rect 136160 679370 136250 679610
rect 136490 679370 136600 679610
rect 136840 679370 136930 679610
rect 137170 679370 137260 679610
rect 137500 679370 137590 679610
rect 137830 679370 137940 679610
rect 138180 679370 138270 679610
rect 138510 679370 138600 679610
rect 138840 679370 138930 679610
rect 139170 679370 139280 679610
rect 139520 679370 139610 679610
rect 139850 679370 139940 679610
rect 140180 679370 140270 679610
rect 140510 679370 140620 679610
rect 140860 679370 140950 679610
rect 141190 679370 141280 679610
rect 141520 679370 141610 679610
rect 141850 679370 141960 679610
rect 142200 679370 142290 679610
rect 142530 679370 142620 679610
rect 142860 679370 142950 679610
rect 143190 679370 143300 679610
rect 143540 679370 143630 679610
rect 143870 679370 143960 679610
rect 144200 679370 144290 679610
rect 144530 679370 144550 679610
rect 133550 679260 144550 679370
rect 133550 679020 133570 679260
rect 133810 679020 133920 679260
rect 134160 679020 134250 679260
rect 134490 679020 134580 679260
rect 134820 679020 134910 679260
rect 135150 679020 135260 679260
rect 135500 679020 135590 679260
rect 135830 679020 135920 679260
rect 136160 679020 136250 679260
rect 136490 679020 136600 679260
rect 136840 679020 136930 679260
rect 137170 679020 137260 679260
rect 137500 679020 137590 679260
rect 137830 679020 137940 679260
rect 138180 679020 138270 679260
rect 138510 679020 138600 679260
rect 138840 679020 138930 679260
rect 139170 679020 139280 679260
rect 139520 679020 139610 679260
rect 139850 679020 139940 679260
rect 140180 679020 140270 679260
rect 140510 679020 140620 679260
rect 140860 679020 140950 679260
rect 141190 679020 141280 679260
rect 141520 679020 141610 679260
rect 141850 679020 141960 679260
rect 142200 679020 142290 679260
rect 142530 679020 142620 679260
rect 142860 679020 142950 679260
rect 143190 679020 143300 679260
rect 143540 679020 143630 679260
rect 143870 679020 143960 679260
rect 144200 679020 144290 679260
rect 144530 679020 144550 679260
rect 133550 678930 144550 679020
rect 133550 678690 133570 678930
rect 133810 678690 133920 678930
rect 134160 678690 134250 678930
rect 134490 678690 134580 678930
rect 134820 678690 134910 678930
rect 135150 678690 135260 678930
rect 135500 678690 135590 678930
rect 135830 678690 135920 678930
rect 136160 678690 136250 678930
rect 136490 678690 136600 678930
rect 136840 678690 136930 678930
rect 137170 678690 137260 678930
rect 137500 678690 137590 678930
rect 137830 678690 137940 678930
rect 138180 678690 138270 678930
rect 138510 678690 138600 678930
rect 138840 678690 138930 678930
rect 139170 678690 139280 678930
rect 139520 678690 139610 678930
rect 139850 678690 139940 678930
rect 140180 678690 140270 678930
rect 140510 678690 140620 678930
rect 140860 678690 140950 678930
rect 141190 678690 141280 678930
rect 141520 678690 141610 678930
rect 141850 678690 141960 678930
rect 142200 678690 142290 678930
rect 142530 678690 142620 678930
rect 142860 678690 142950 678930
rect 143190 678690 143300 678930
rect 143540 678690 143630 678930
rect 143870 678690 143960 678930
rect 144200 678690 144290 678930
rect 144530 678690 144550 678930
rect 133550 678600 144550 678690
rect 133550 678360 133570 678600
rect 133810 678360 133920 678600
rect 134160 678360 134250 678600
rect 134490 678360 134580 678600
rect 134820 678360 134910 678600
rect 135150 678360 135260 678600
rect 135500 678360 135590 678600
rect 135830 678360 135920 678600
rect 136160 678360 136250 678600
rect 136490 678360 136600 678600
rect 136840 678360 136930 678600
rect 137170 678360 137260 678600
rect 137500 678360 137590 678600
rect 137830 678360 137940 678600
rect 138180 678360 138270 678600
rect 138510 678360 138600 678600
rect 138840 678360 138930 678600
rect 139170 678360 139280 678600
rect 139520 678360 139610 678600
rect 139850 678360 139940 678600
rect 140180 678360 140270 678600
rect 140510 678360 140620 678600
rect 140860 678360 140950 678600
rect 141190 678360 141280 678600
rect 141520 678360 141610 678600
rect 141850 678360 141960 678600
rect 142200 678360 142290 678600
rect 142530 678360 142620 678600
rect 142860 678360 142950 678600
rect 143190 678360 143300 678600
rect 143540 678360 143630 678600
rect 143870 678360 143960 678600
rect 144200 678360 144290 678600
rect 144530 678360 144550 678600
rect 133550 678270 144550 678360
rect 133550 678030 133570 678270
rect 133810 678030 133920 678270
rect 134160 678030 134250 678270
rect 134490 678030 134580 678270
rect 134820 678030 134910 678270
rect 135150 678030 135260 678270
rect 135500 678030 135590 678270
rect 135830 678030 135920 678270
rect 136160 678030 136250 678270
rect 136490 678030 136600 678270
rect 136840 678030 136930 678270
rect 137170 678030 137260 678270
rect 137500 678030 137590 678270
rect 137830 678030 137940 678270
rect 138180 678030 138270 678270
rect 138510 678030 138600 678270
rect 138840 678030 138930 678270
rect 139170 678030 139280 678270
rect 139520 678030 139610 678270
rect 139850 678030 139940 678270
rect 140180 678030 140270 678270
rect 140510 678030 140620 678270
rect 140860 678030 140950 678270
rect 141190 678030 141280 678270
rect 141520 678030 141610 678270
rect 141850 678030 141960 678270
rect 142200 678030 142290 678270
rect 142530 678030 142620 678270
rect 142860 678030 142950 678270
rect 143190 678030 143300 678270
rect 143540 678030 143630 678270
rect 143870 678030 143960 678270
rect 144200 678030 144290 678270
rect 144530 678030 144550 678270
rect 133550 677920 144550 678030
rect 133550 677680 133570 677920
rect 133810 677680 133920 677920
rect 134160 677680 134250 677920
rect 134490 677680 134580 677920
rect 134820 677680 134910 677920
rect 135150 677680 135260 677920
rect 135500 677680 135590 677920
rect 135830 677680 135920 677920
rect 136160 677680 136250 677920
rect 136490 677680 136600 677920
rect 136840 677680 136930 677920
rect 137170 677680 137260 677920
rect 137500 677680 137590 677920
rect 137830 677680 137940 677920
rect 138180 677680 138270 677920
rect 138510 677680 138600 677920
rect 138840 677680 138930 677920
rect 139170 677680 139280 677920
rect 139520 677680 139610 677920
rect 139850 677680 139940 677920
rect 140180 677680 140270 677920
rect 140510 677680 140620 677920
rect 140860 677680 140950 677920
rect 141190 677680 141280 677920
rect 141520 677680 141610 677920
rect 141850 677680 141960 677920
rect 142200 677680 142290 677920
rect 142530 677680 142620 677920
rect 142860 677680 142950 677920
rect 143190 677680 143300 677920
rect 143540 677680 143630 677920
rect 143870 677680 143960 677920
rect 144200 677680 144290 677920
rect 144530 677680 144550 677920
rect 133550 677590 144550 677680
rect 133550 677350 133570 677590
rect 133810 677350 133920 677590
rect 134160 677350 134250 677590
rect 134490 677350 134580 677590
rect 134820 677350 134910 677590
rect 135150 677350 135260 677590
rect 135500 677350 135590 677590
rect 135830 677350 135920 677590
rect 136160 677350 136250 677590
rect 136490 677350 136600 677590
rect 136840 677350 136930 677590
rect 137170 677350 137260 677590
rect 137500 677350 137590 677590
rect 137830 677350 137940 677590
rect 138180 677350 138270 677590
rect 138510 677350 138600 677590
rect 138840 677350 138930 677590
rect 139170 677350 139280 677590
rect 139520 677350 139610 677590
rect 139850 677350 139940 677590
rect 140180 677350 140270 677590
rect 140510 677350 140620 677590
rect 140860 677350 140950 677590
rect 141190 677350 141280 677590
rect 141520 677350 141610 677590
rect 141850 677350 141960 677590
rect 142200 677350 142290 677590
rect 142530 677350 142620 677590
rect 142860 677350 142950 677590
rect 143190 677350 143300 677590
rect 143540 677350 143630 677590
rect 143870 677350 143960 677590
rect 144200 677350 144290 677590
rect 144530 677350 144550 677590
rect 133550 677260 144550 677350
rect 133550 677020 133570 677260
rect 133810 677020 133920 677260
rect 134160 677020 134250 677260
rect 134490 677020 134580 677260
rect 134820 677020 134910 677260
rect 135150 677020 135260 677260
rect 135500 677020 135590 677260
rect 135830 677020 135920 677260
rect 136160 677020 136250 677260
rect 136490 677020 136600 677260
rect 136840 677020 136930 677260
rect 137170 677020 137260 677260
rect 137500 677020 137590 677260
rect 137830 677020 137940 677260
rect 138180 677020 138270 677260
rect 138510 677020 138600 677260
rect 138840 677020 138930 677260
rect 139170 677020 139280 677260
rect 139520 677020 139610 677260
rect 139850 677020 139940 677260
rect 140180 677020 140270 677260
rect 140510 677020 140620 677260
rect 140860 677020 140950 677260
rect 141190 677020 141280 677260
rect 141520 677020 141610 677260
rect 141850 677020 141960 677260
rect 142200 677020 142290 677260
rect 142530 677020 142620 677260
rect 142860 677020 142950 677260
rect 143190 677020 143300 677260
rect 143540 677020 143630 677260
rect 143870 677020 143960 677260
rect 144200 677020 144290 677260
rect 144530 677020 144550 677260
rect 133550 676930 144550 677020
rect 133550 676690 133570 676930
rect 133810 676690 133920 676930
rect 134160 676690 134250 676930
rect 134490 676690 134580 676930
rect 134820 676690 134910 676930
rect 135150 676690 135260 676930
rect 135500 676690 135590 676930
rect 135830 676690 135920 676930
rect 136160 676690 136250 676930
rect 136490 676690 136600 676930
rect 136840 676690 136930 676930
rect 137170 676690 137260 676930
rect 137500 676690 137590 676930
rect 137830 676690 137940 676930
rect 138180 676690 138270 676930
rect 138510 676690 138600 676930
rect 138840 676690 138930 676930
rect 139170 676690 139280 676930
rect 139520 676690 139610 676930
rect 139850 676690 139940 676930
rect 140180 676690 140270 676930
rect 140510 676690 140620 676930
rect 140860 676690 140950 676930
rect 141190 676690 141280 676930
rect 141520 676690 141610 676930
rect 141850 676690 141960 676930
rect 142200 676690 142290 676930
rect 142530 676690 142620 676930
rect 142860 676690 142950 676930
rect 143190 676690 143300 676930
rect 143540 676690 143630 676930
rect 143870 676690 143960 676930
rect 144200 676690 144290 676930
rect 144530 676690 144550 676930
rect 133550 676580 144550 676690
rect 133550 676340 133570 676580
rect 133810 676340 133920 676580
rect 134160 676340 134250 676580
rect 134490 676340 134580 676580
rect 134820 676340 134910 676580
rect 135150 676340 135260 676580
rect 135500 676340 135590 676580
rect 135830 676340 135920 676580
rect 136160 676340 136250 676580
rect 136490 676340 136600 676580
rect 136840 676340 136930 676580
rect 137170 676340 137260 676580
rect 137500 676340 137590 676580
rect 137830 676340 137940 676580
rect 138180 676340 138270 676580
rect 138510 676340 138600 676580
rect 138840 676340 138930 676580
rect 139170 676340 139280 676580
rect 139520 676340 139610 676580
rect 139850 676340 139940 676580
rect 140180 676340 140270 676580
rect 140510 676340 140620 676580
rect 140860 676340 140950 676580
rect 141190 676340 141280 676580
rect 141520 676340 141610 676580
rect 141850 676340 141960 676580
rect 142200 676340 142290 676580
rect 142530 676340 142620 676580
rect 142860 676340 142950 676580
rect 143190 676340 143300 676580
rect 143540 676340 143630 676580
rect 143870 676340 143960 676580
rect 144200 676340 144290 676580
rect 144530 676340 144550 676580
rect 133550 676250 144550 676340
rect 133550 676010 133570 676250
rect 133810 676010 133920 676250
rect 134160 676010 134250 676250
rect 134490 676010 134580 676250
rect 134820 676010 134910 676250
rect 135150 676010 135260 676250
rect 135500 676010 135590 676250
rect 135830 676010 135920 676250
rect 136160 676010 136250 676250
rect 136490 676010 136600 676250
rect 136840 676010 136930 676250
rect 137170 676010 137260 676250
rect 137500 676010 137590 676250
rect 137830 676010 137940 676250
rect 138180 676010 138270 676250
rect 138510 676010 138600 676250
rect 138840 676010 138930 676250
rect 139170 676010 139280 676250
rect 139520 676010 139610 676250
rect 139850 676010 139940 676250
rect 140180 676010 140270 676250
rect 140510 676010 140620 676250
rect 140860 676010 140950 676250
rect 141190 676010 141280 676250
rect 141520 676010 141610 676250
rect 141850 676010 141960 676250
rect 142200 676010 142290 676250
rect 142530 676010 142620 676250
rect 142860 676010 142950 676250
rect 143190 676010 143300 676250
rect 143540 676010 143630 676250
rect 143870 676010 143960 676250
rect 144200 676010 144290 676250
rect 144530 676010 144550 676250
rect 133550 675920 144550 676010
rect 133550 675680 133570 675920
rect 133810 675680 133920 675920
rect 134160 675680 134250 675920
rect 134490 675680 134580 675920
rect 134820 675680 134910 675920
rect 135150 675680 135260 675920
rect 135500 675680 135590 675920
rect 135830 675680 135920 675920
rect 136160 675680 136250 675920
rect 136490 675680 136600 675920
rect 136840 675680 136930 675920
rect 137170 675680 137260 675920
rect 137500 675680 137590 675920
rect 137830 675680 137940 675920
rect 138180 675680 138270 675920
rect 138510 675680 138600 675920
rect 138840 675680 138930 675920
rect 139170 675680 139280 675920
rect 139520 675680 139610 675920
rect 139850 675680 139940 675920
rect 140180 675680 140270 675920
rect 140510 675680 140620 675920
rect 140860 675680 140950 675920
rect 141190 675680 141280 675920
rect 141520 675680 141610 675920
rect 141850 675680 141960 675920
rect 142200 675680 142290 675920
rect 142530 675680 142620 675920
rect 142860 675680 142950 675920
rect 143190 675680 143300 675920
rect 143540 675680 143630 675920
rect 143870 675680 143960 675920
rect 144200 675680 144290 675920
rect 144530 675680 144550 675920
rect 133550 675590 144550 675680
rect 133550 675350 133570 675590
rect 133810 675350 133920 675590
rect 134160 675350 134250 675590
rect 134490 675350 134580 675590
rect 134820 675350 134910 675590
rect 135150 675350 135260 675590
rect 135500 675350 135590 675590
rect 135830 675350 135920 675590
rect 136160 675350 136250 675590
rect 136490 675350 136600 675590
rect 136840 675350 136930 675590
rect 137170 675350 137260 675590
rect 137500 675350 137590 675590
rect 137830 675350 137940 675590
rect 138180 675350 138270 675590
rect 138510 675350 138600 675590
rect 138840 675350 138930 675590
rect 139170 675350 139280 675590
rect 139520 675350 139610 675590
rect 139850 675350 139940 675590
rect 140180 675350 140270 675590
rect 140510 675350 140620 675590
rect 140860 675350 140950 675590
rect 141190 675350 141280 675590
rect 141520 675350 141610 675590
rect 141850 675350 141960 675590
rect 142200 675350 142290 675590
rect 142530 675350 142620 675590
rect 142860 675350 142950 675590
rect 143190 675350 143300 675590
rect 143540 675350 143630 675590
rect 143870 675350 143960 675590
rect 144200 675350 144290 675590
rect 144530 675350 144550 675590
rect 133550 675240 144550 675350
rect 133550 675000 133570 675240
rect 133810 675000 133920 675240
rect 134160 675000 134250 675240
rect 134490 675000 134580 675240
rect 134820 675000 134910 675240
rect 135150 675000 135260 675240
rect 135500 675000 135590 675240
rect 135830 675000 135920 675240
rect 136160 675000 136250 675240
rect 136490 675000 136600 675240
rect 136840 675000 136930 675240
rect 137170 675000 137260 675240
rect 137500 675000 137590 675240
rect 137830 675000 137940 675240
rect 138180 675000 138270 675240
rect 138510 675000 138600 675240
rect 138840 675000 138930 675240
rect 139170 675000 139280 675240
rect 139520 675000 139610 675240
rect 139850 675000 139940 675240
rect 140180 675000 140270 675240
rect 140510 675000 140620 675240
rect 140860 675000 140950 675240
rect 141190 675000 141280 675240
rect 141520 675000 141610 675240
rect 141850 675000 141960 675240
rect 142200 675000 142290 675240
rect 142530 675000 142620 675240
rect 142860 675000 142950 675240
rect 143190 675000 143300 675240
rect 143540 675000 143630 675240
rect 143870 675000 143960 675240
rect 144200 675000 144290 675240
rect 144530 675000 144550 675240
rect 133550 674910 144550 675000
rect 133550 674670 133570 674910
rect 133810 674670 133920 674910
rect 134160 674670 134250 674910
rect 134490 674670 134580 674910
rect 134820 674670 134910 674910
rect 135150 674670 135260 674910
rect 135500 674670 135590 674910
rect 135830 674670 135920 674910
rect 136160 674670 136250 674910
rect 136490 674670 136600 674910
rect 136840 674670 136930 674910
rect 137170 674670 137260 674910
rect 137500 674670 137590 674910
rect 137830 674670 137940 674910
rect 138180 674670 138270 674910
rect 138510 674670 138600 674910
rect 138840 674670 138930 674910
rect 139170 674670 139280 674910
rect 139520 674670 139610 674910
rect 139850 674670 139940 674910
rect 140180 674670 140270 674910
rect 140510 674670 140620 674910
rect 140860 674670 140950 674910
rect 141190 674670 141280 674910
rect 141520 674670 141610 674910
rect 141850 674670 141960 674910
rect 142200 674670 142290 674910
rect 142530 674670 142620 674910
rect 142860 674670 142950 674910
rect 143190 674670 143300 674910
rect 143540 674670 143630 674910
rect 143870 674670 143960 674910
rect 144200 674670 144290 674910
rect 144530 674670 144550 674910
rect 133550 674580 144550 674670
rect 133550 674340 133570 674580
rect 133810 674340 133920 674580
rect 134160 674340 134250 674580
rect 134490 674340 134580 674580
rect 134820 674340 134910 674580
rect 135150 674340 135260 674580
rect 135500 674340 135590 674580
rect 135830 674340 135920 674580
rect 136160 674340 136250 674580
rect 136490 674340 136600 674580
rect 136840 674340 136930 674580
rect 137170 674340 137260 674580
rect 137500 674340 137590 674580
rect 137830 674340 137940 674580
rect 138180 674340 138270 674580
rect 138510 674340 138600 674580
rect 138840 674340 138930 674580
rect 139170 674340 139280 674580
rect 139520 674340 139610 674580
rect 139850 674340 139940 674580
rect 140180 674340 140270 674580
rect 140510 674340 140620 674580
rect 140860 674340 140950 674580
rect 141190 674340 141280 674580
rect 141520 674340 141610 674580
rect 141850 674340 141960 674580
rect 142200 674340 142290 674580
rect 142530 674340 142620 674580
rect 142860 674340 142950 674580
rect 143190 674340 143300 674580
rect 143540 674340 143630 674580
rect 143870 674340 143960 674580
rect 144200 674340 144290 674580
rect 144530 674340 144550 674580
rect 133550 674250 144550 674340
rect 133550 674010 133570 674250
rect 133810 674010 133920 674250
rect 134160 674010 134250 674250
rect 134490 674010 134580 674250
rect 134820 674010 134910 674250
rect 135150 674010 135260 674250
rect 135500 674010 135590 674250
rect 135830 674010 135920 674250
rect 136160 674010 136250 674250
rect 136490 674010 136600 674250
rect 136840 674010 136930 674250
rect 137170 674010 137260 674250
rect 137500 674010 137590 674250
rect 137830 674010 137940 674250
rect 138180 674010 138270 674250
rect 138510 674010 138600 674250
rect 138840 674010 138930 674250
rect 139170 674010 139280 674250
rect 139520 674010 139610 674250
rect 139850 674010 139940 674250
rect 140180 674010 140270 674250
rect 140510 674010 140620 674250
rect 140860 674010 140950 674250
rect 141190 674010 141280 674250
rect 141520 674010 141610 674250
rect 141850 674010 141960 674250
rect 142200 674010 142290 674250
rect 142530 674010 142620 674250
rect 142860 674010 142950 674250
rect 143190 674010 143300 674250
rect 143540 674010 143630 674250
rect 143870 674010 143960 674250
rect 144200 674010 144290 674250
rect 144530 674010 144550 674250
rect 133550 673900 144550 674010
rect 133550 673660 133570 673900
rect 133810 673660 133920 673900
rect 134160 673660 134250 673900
rect 134490 673660 134580 673900
rect 134820 673660 134910 673900
rect 135150 673660 135260 673900
rect 135500 673660 135590 673900
rect 135830 673660 135920 673900
rect 136160 673660 136250 673900
rect 136490 673660 136600 673900
rect 136840 673660 136930 673900
rect 137170 673660 137260 673900
rect 137500 673660 137590 673900
rect 137830 673660 137940 673900
rect 138180 673660 138270 673900
rect 138510 673660 138600 673900
rect 138840 673660 138930 673900
rect 139170 673660 139280 673900
rect 139520 673660 139610 673900
rect 139850 673660 139940 673900
rect 140180 673660 140270 673900
rect 140510 673660 140620 673900
rect 140860 673660 140950 673900
rect 141190 673660 141280 673900
rect 141520 673660 141610 673900
rect 141850 673660 141960 673900
rect 142200 673660 142290 673900
rect 142530 673660 142620 673900
rect 142860 673660 142950 673900
rect 143190 673660 143300 673900
rect 143540 673660 143630 673900
rect 143870 673660 143960 673900
rect 144200 673660 144290 673900
rect 144530 673660 144550 673900
rect 133550 673570 144550 673660
rect 133550 673330 133570 673570
rect 133810 673330 133920 673570
rect 134160 673330 134250 673570
rect 134490 673330 134580 673570
rect 134820 673330 134910 673570
rect 135150 673330 135260 673570
rect 135500 673330 135590 673570
rect 135830 673330 135920 673570
rect 136160 673330 136250 673570
rect 136490 673330 136600 673570
rect 136840 673330 136930 673570
rect 137170 673330 137260 673570
rect 137500 673330 137590 673570
rect 137830 673330 137940 673570
rect 138180 673330 138270 673570
rect 138510 673330 138600 673570
rect 138840 673330 138930 673570
rect 139170 673330 139280 673570
rect 139520 673330 139610 673570
rect 139850 673330 139940 673570
rect 140180 673330 140270 673570
rect 140510 673330 140620 673570
rect 140860 673330 140950 673570
rect 141190 673330 141280 673570
rect 141520 673330 141610 673570
rect 141850 673330 141960 673570
rect 142200 673330 142290 673570
rect 142530 673330 142620 673570
rect 142860 673330 142950 673570
rect 143190 673330 143300 673570
rect 143540 673330 143630 673570
rect 143870 673330 143960 673570
rect 144200 673330 144290 673570
rect 144530 673330 144550 673570
rect 133550 673240 144550 673330
rect 133550 673000 133570 673240
rect 133810 673000 133920 673240
rect 134160 673000 134250 673240
rect 134490 673000 134580 673240
rect 134820 673000 134910 673240
rect 135150 673000 135260 673240
rect 135500 673000 135590 673240
rect 135830 673000 135920 673240
rect 136160 673000 136250 673240
rect 136490 673000 136600 673240
rect 136840 673000 136930 673240
rect 137170 673000 137260 673240
rect 137500 673000 137590 673240
rect 137830 673000 137940 673240
rect 138180 673000 138270 673240
rect 138510 673000 138600 673240
rect 138840 673000 138930 673240
rect 139170 673000 139280 673240
rect 139520 673000 139610 673240
rect 139850 673000 139940 673240
rect 140180 673000 140270 673240
rect 140510 673000 140620 673240
rect 140860 673000 140950 673240
rect 141190 673000 141280 673240
rect 141520 673000 141610 673240
rect 141850 673000 141960 673240
rect 142200 673000 142290 673240
rect 142530 673000 142620 673240
rect 142860 673000 142950 673240
rect 143190 673000 143300 673240
rect 143540 673000 143630 673240
rect 143870 673000 143960 673240
rect 144200 673000 144290 673240
rect 144530 673000 144550 673240
rect 133550 672910 144550 673000
rect 133550 672670 133570 672910
rect 133810 672670 133920 672910
rect 134160 672670 134250 672910
rect 134490 672670 134580 672910
rect 134820 672670 134910 672910
rect 135150 672670 135260 672910
rect 135500 672670 135590 672910
rect 135830 672670 135920 672910
rect 136160 672670 136250 672910
rect 136490 672670 136600 672910
rect 136840 672670 136930 672910
rect 137170 672670 137260 672910
rect 137500 672670 137590 672910
rect 137830 672670 137940 672910
rect 138180 672670 138270 672910
rect 138510 672670 138600 672910
rect 138840 672670 138930 672910
rect 139170 672670 139280 672910
rect 139520 672670 139610 672910
rect 139850 672670 139940 672910
rect 140180 672670 140270 672910
rect 140510 672670 140620 672910
rect 140860 672670 140950 672910
rect 141190 672670 141280 672910
rect 141520 672670 141610 672910
rect 141850 672670 141960 672910
rect 142200 672670 142290 672910
rect 142530 672670 142620 672910
rect 142860 672670 142950 672910
rect 143190 672670 143300 672910
rect 143540 672670 143630 672910
rect 143870 672670 143960 672910
rect 144200 672670 144290 672910
rect 144530 672670 144550 672910
rect 133550 672560 144550 672670
rect 133550 672320 133570 672560
rect 133810 672320 133920 672560
rect 134160 672320 134250 672560
rect 134490 672320 134580 672560
rect 134820 672320 134910 672560
rect 135150 672320 135260 672560
rect 135500 672320 135590 672560
rect 135830 672320 135920 672560
rect 136160 672320 136250 672560
rect 136490 672320 136600 672560
rect 136840 672320 136930 672560
rect 137170 672320 137260 672560
rect 137500 672320 137590 672560
rect 137830 672320 137940 672560
rect 138180 672320 138270 672560
rect 138510 672320 138600 672560
rect 138840 672320 138930 672560
rect 139170 672320 139280 672560
rect 139520 672320 139610 672560
rect 139850 672320 139940 672560
rect 140180 672320 140270 672560
rect 140510 672320 140620 672560
rect 140860 672320 140950 672560
rect 141190 672320 141280 672560
rect 141520 672320 141610 672560
rect 141850 672320 141960 672560
rect 142200 672320 142290 672560
rect 142530 672320 142620 672560
rect 142860 672320 142950 672560
rect 143190 672320 143300 672560
rect 143540 672320 143630 672560
rect 143870 672320 143960 672560
rect 144200 672320 144290 672560
rect 144530 672320 144550 672560
rect 133550 672300 144550 672320
rect 144930 683280 155930 683300
rect 144930 683040 144950 683280
rect 145190 683040 145300 683280
rect 145540 683040 145630 683280
rect 145870 683040 145960 683280
rect 146200 683040 146290 683280
rect 146530 683040 146640 683280
rect 146880 683040 146970 683280
rect 147210 683040 147300 683280
rect 147540 683040 147630 683280
rect 147870 683040 147980 683280
rect 148220 683040 148310 683280
rect 148550 683040 148640 683280
rect 148880 683040 148970 683280
rect 149210 683040 149320 683280
rect 149560 683040 149650 683280
rect 149890 683040 149980 683280
rect 150220 683040 150310 683280
rect 150550 683040 150660 683280
rect 150900 683040 150990 683280
rect 151230 683040 151320 683280
rect 151560 683040 151650 683280
rect 151890 683040 152000 683280
rect 152240 683040 152330 683280
rect 152570 683040 152660 683280
rect 152900 683040 152990 683280
rect 153230 683040 153340 683280
rect 153580 683040 153670 683280
rect 153910 683040 154000 683280
rect 154240 683040 154330 683280
rect 154570 683040 154680 683280
rect 154920 683040 155010 683280
rect 155250 683040 155340 683280
rect 155580 683040 155670 683280
rect 155910 683040 155930 683280
rect 144930 682950 155930 683040
rect 144930 682710 144950 682950
rect 145190 682710 145300 682950
rect 145540 682710 145630 682950
rect 145870 682710 145960 682950
rect 146200 682710 146290 682950
rect 146530 682710 146640 682950
rect 146880 682710 146970 682950
rect 147210 682710 147300 682950
rect 147540 682710 147630 682950
rect 147870 682710 147980 682950
rect 148220 682710 148310 682950
rect 148550 682710 148640 682950
rect 148880 682710 148970 682950
rect 149210 682710 149320 682950
rect 149560 682710 149650 682950
rect 149890 682710 149980 682950
rect 150220 682710 150310 682950
rect 150550 682710 150660 682950
rect 150900 682710 150990 682950
rect 151230 682710 151320 682950
rect 151560 682710 151650 682950
rect 151890 682710 152000 682950
rect 152240 682710 152330 682950
rect 152570 682710 152660 682950
rect 152900 682710 152990 682950
rect 153230 682710 153340 682950
rect 153580 682710 153670 682950
rect 153910 682710 154000 682950
rect 154240 682710 154330 682950
rect 154570 682710 154680 682950
rect 154920 682710 155010 682950
rect 155250 682710 155340 682950
rect 155580 682710 155670 682950
rect 155910 682710 155930 682950
rect 144930 682620 155930 682710
rect 144930 682380 144950 682620
rect 145190 682380 145300 682620
rect 145540 682380 145630 682620
rect 145870 682380 145960 682620
rect 146200 682380 146290 682620
rect 146530 682380 146640 682620
rect 146880 682380 146970 682620
rect 147210 682380 147300 682620
rect 147540 682380 147630 682620
rect 147870 682380 147980 682620
rect 148220 682380 148310 682620
rect 148550 682380 148640 682620
rect 148880 682380 148970 682620
rect 149210 682380 149320 682620
rect 149560 682380 149650 682620
rect 149890 682380 149980 682620
rect 150220 682380 150310 682620
rect 150550 682380 150660 682620
rect 150900 682380 150990 682620
rect 151230 682380 151320 682620
rect 151560 682380 151650 682620
rect 151890 682380 152000 682620
rect 152240 682380 152330 682620
rect 152570 682380 152660 682620
rect 152900 682380 152990 682620
rect 153230 682380 153340 682620
rect 153580 682380 153670 682620
rect 153910 682380 154000 682620
rect 154240 682380 154330 682620
rect 154570 682380 154680 682620
rect 154920 682380 155010 682620
rect 155250 682380 155340 682620
rect 155580 682380 155670 682620
rect 155910 682380 155930 682620
rect 144930 682290 155930 682380
rect 144930 682050 144950 682290
rect 145190 682050 145300 682290
rect 145540 682050 145630 682290
rect 145870 682050 145960 682290
rect 146200 682050 146290 682290
rect 146530 682050 146640 682290
rect 146880 682050 146970 682290
rect 147210 682050 147300 682290
rect 147540 682050 147630 682290
rect 147870 682050 147980 682290
rect 148220 682050 148310 682290
rect 148550 682050 148640 682290
rect 148880 682050 148970 682290
rect 149210 682050 149320 682290
rect 149560 682050 149650 682290
rect 149890 682050 149980 682290
rect 150220 682050 150310 682290
rect 150550 682050 150660 682290
rect 150900 682050 150990 682290
rect 151230 682050 151320 682290
rect 151560 682050 151650 682290
rect 151890 682050 152000 682290
rect 152240 682050 152330 682290
rect 152570 682050 152660 682290
rect 152900 682050 152990 682290
rect 153230 682050 153340 682290
rect 153580 682050 153670 682290
rect 153910 682050 154000 682290
rect 154240 682050 154330 682290
rect 154570 682050 154680 682290
rect 154920 682050 155010 682290
rect 155250 682050 155340 682290
rect 155580 682050 155670 682290
rect 155910 682050 155930 682290
rect 144930 681940 155930 682050
rect 144930 681700 144950 681940
rect 145190 681700 145300 681940
rect 145540 681700 145630 681940
rect 145870 681700 145960 681940
rect 146200 681700 146290 681940
rect 146530 681700 146640 681940
rect 146880 681700 146970 681940
rect 147210 681700 147300 681940
rect 147540 681700 147630 681940
rect 147870 681700 147980 681940
rect 148220 681700 148310 681940
rect 148550 681700 148640 681940
rect 148880 681700 148970 681940
rect 149210 681700 149320 681940
rect 149560 681700 149650 681940
rect 149890 681700 149980 681940
rect 150220 681700 150310 681940
rect 150550 681700 150660 681940
rect 150900 681700 150990 681940
rect 151230 681700 151320 681940
rect 151560 681700 151650 681940
rect 151890 681700 152000 681940
rect 152240 681700 152330 681940
rect 152570 681700 152660 681940
rect 152900 681700 152990 681940
rect 153230 681700 153340 681940
rect 153580 681700 153670 681940
rect 153910 681700 154000 681940
rect 154240 681700 154330 681940
rect 154570 681700 154680 681940
rect 154920 681700 155010 681940
rect 155250 681700 155340 681940
rect 155580 681700 155670 681940
rect 155910 681700 155930 681940
rect 144930 681610 155930 681700
rect 144930 681370 144950 681610
rect 145190 681370 145300 681610
rect 145540 681370 145630 681610
rect 145870 681370 145960 681610
rect 146200 681370 146290 681610
rect 146530 681370 146640 681610
rect 146880 681370 146970 681610
rect 147210 681370 147300 681610
rect 147540 681370 147630 681610
rect 147870 681370 147980 681610
rect 148220 681370 148310 681610
rect 148550 681370 148640 681610
rect 148880 681370 148970 681610
rect 149210 681370 149320 681610
rect 149560 681370 149650 681610
rect 149890 681370 149980 681610
rect 150220 681370 150310 681610
rect 150550 681370 150660 681610
rect 150900 681370 150990 681610
rect 151230 681370 151320 681610
rect 151560 681370 151650 681610
rect 151890 681370 152000 681610
rect 152240 681370 152330 681610
rect 152570 681370 152660 681610
rect 152900 681370 152990 681610
rect 153230 681370 153340 681610
rect 153580 681370 153670 681610
rect 153910 681370 154000 681610
rect 154240 681370 154330 681610
rect 154570 681370 154680 681610
rect 154920 681370 155010 681610
rect 155250 681370 155340 681610
rect 155580 681370 155670 681610
rect 155910 681370 155930 681610
rect 144930 681280 155930 681370
rect 144930 681040 144950 681280
rect 145190 681040 145300 681280
rect 145540 681040 145630 681280
rect 145870 681040 145960 681280
rect 146200 681040 146290 681280
rect 146530 681040 146640 681280
rect 146880 681040 146970 681280
rect 147210 681040 147300 681280
rect 147540 681040 147630 681280
rect 147870 681040 147980 681280
rect 148220 681040 148310 681280
rect 148550 681040 148640 681280
rect 148880 681040 148970 681280
rect 149210 681040 149320 681280
rect 149560 681040 149650 681280
rect 149890 681040 149980 681280
rect 150220 681040 150310 681280
rect 150550 681040 150660 681280
rect 150900 681040 150990 681280
rect 151230 681040 151320 681280
rect 151560 681040 151650 681280
rect 151890 681040 152000 681280
rect 152240 681040 152330 681280
rect 152570 681040 152660 681280
rect 152900 681040 152990 681280
rect 153230 681040 153340 681280
rect 153580 681040 153670 681280
rect 153910 681040 154000 681280
rect 154240 681040 154330 681280
rect 154570 681040 154680 681280
rect 154920 681040 155010 681280
rect 155250 681040 155340 681280
rect 155580 681040 155670 681280
rect 155910 681040 155930 681280
rect 144930 680950 155930 681040
rect 144930 680710 144950 680950
rect 145190 680710 145300 680950
rect 145540 680710 145630 680950
rect 145870 680710 145960 680950
rect 146200 680710 146290 680950
rect 146530 680710 146640 680950
rect 146880 680710 146970 680950
rect 147210 680710 147300 680950
rect 147540 680710 147630 680950
rect 147870 680710 147980 680950
rect 148220 680710 148310 680950
rect 148550 680710 148640 680950
rect 148880 680710 148970 680950
rect 149210 680710 149320 680950
rect 149560 680710 149650 680950
rect 149890 680710 149980 680950
rect 150220 680710 150310 680950
rect 150550 680710 150660 680950
rect 150900 680710 150990 680950
rect 151230 680710 151320 680950
rect 151560 680710 151650 680950
rect 151890 680710 152000 680950
rect 152240 680710 152330 680950
rect 152570 680710 152660 680950
rect 152900 680710 152990 680950
rect 153230 680710 153340 680950
rect 153580 680710 153670 680950
rect 153910 680710 154000 680950
rect 154240 680710 154330 680950
rect 154570 680710 154680 680950
rect 154920 680710 155010 680950
rect 155250 680710 155340 680950
rect 155580 680710 155670 680950
rect 155910 680710 155930 680950
rect 144930 680600 155930 680710
rect 144930 680360 144950 680600
rect 145190 680360 145300 680600
rect 145540 680360 145630 680600
rect 145870 680360 145960 680600
rect 146200 680360 146290 680600
rect 146530 680360 146640 680600
rect 146880 680360 146970 680600
rect 147210 680360 147300 680600
rect 147540 680360 147630 680600
rect 147870 680360 147980 680600
rect 148220 680360 148310 680600
rect 148550 680360 148640 680600
rect 148880 680360 148970 680600
rect 149210 680360 149320 680600
rect 149560 680360 149650 680600
rect 149890 680360 149980 680600
rect 150220 680360 150310 680600
rect 150550 680360 150660 680600
rect 150900 680360 150990 680600
rect 151230 680360 151320 680600
rect 151560 680360 151650 680600
rect 151890 680360 152000 680600
rect 152240 680360 152330 680600
rect 152570 680360 152660 680600
rect 152900 680360 152990 680600
rect 153230 680360 153340 680600
rect 153580 680360 153670 680600
rect 153910 680360 154000 680600
rect 154240 680360 154330 680600
rect 154570 680360 154680 680600
rect 154920 680360 155010 680600
rect 155250 680360 155340 680600
rect 155580 680360 155670 680600
rect 155910 680360 155930 680600
rect 144930 680270 155930 680360
rect 144930 680030 144950 680270
rect 145190 680030 145300 680270
rect 145540 680030 145630 680270
rect 145870 680030 145960 680270
rect 146200 680030 146290 680270
rect 146530 680030 146640 680270
rect 146880 680030 146970 680270
rect 147210 680030 147300 680270
rect 147540 680030 147630 680270
rect 147870 680030 147980 680270
rect 148220 680030 148310 680270
rect 148550 680030 148640 680270
rect 148880 680030 148970 680270
rect 149210 680030 149320 680270
rect 149560 680030 149650 680270
rect 149890 680030 149980 680270
rect 150220 680030 150310 680270
rect 150550 680030 150660 680270
rect 150900 680030 150990 680270
rect 151230 680030 151320 680270
rect 151560 680030 151650 680270
rect 151890 680030 152000 680270
rect 152240 680030 152330 680270
rect 152570 680030 152660 680270
rect 152900 680030 152990 680270
rect 153230 680030 153340 680270
rect 153580 680030 153670 680270
rect 153910 680030 154000 680270
rect 154240 680030 154330 680270
rect 154570 680030 154680 680270
rect 154920 680030 155010 680270
rect 155250 680030 155340 680270
rect 155580 680030 155670 680270
rect 155910 680030 155930 680270
rect 144930 679940 155930 680030
rect 144930 679700 144950 679940
rect 145190 679700 145300 679940
rect 145540 679700 145630 679940
rect 145870 679700 145960 679940
rect 146200 679700 146290 679940
rect 146530 679700 146640 679940
rect 146880 679700 146970 679940
rect 147210 679700 147300 679940
rect 147540 679700 147630 679940
rect 147870 679700 147980 679940
rect 148220 679700 148310 679940
rect 148550 679700 148640 679940
rect 148880 679700 148970 679940
rect 149210 679700 149320 679940
rect 149560 679700 149650 679940
rect 149890 679700 149980 679940
rect 150220 679700 150310 679940
rect 150550 679700 150660 679940
rect 150900 679700 150990 679940
rect 151230 679700 151320 679940
rect 151560 679700 151650 679940
rect 151890 679700 152000 679940
rect 152240 679700 152330 679940
rect 152570 679700 152660 679940
rect 152900 679700 152990 679940
rect 153230 679700 153340 679940
rect 153580 679700 153670 679940
rect 153910 679700 154000 679940
rect 154240 679700 154330 679940
rect 154570 679700 154680 679940
rect 154920 679700 155010 679940
rect 155250 679700 155340 679940
rect 155580 679700 155670 679940
rect 155910 679700 155930 679940
rect 144930 679610 155930 679700
rect 144930 679370 144950 679610
rect 145190 679370 145300 679610
rect 145540 679370 145630 679610
rect 145870 679370 145960 679610
rect 146200 679370 146290 679610
rect 146530 679370 146640 679610
rect 146880 679370 146970 679610
rect 147210 679370 147300 679610
rect 147540 679370 147630 679610
rect 147870 679370 147980 679610
rect 148220 679370 148310 679610
rect 148550 679370 148640 679610
rect 148880 679370 148970 679610
rect 149210 679370 149320 679610
rect 149560 679370 149650 679610
rect 149890 679370 149980 679610
rect 150220 679370 150310 679610
rect 150550 679370 150660 679610
rect 150900 679370 150990 679610
rect 151230 679370 151320 679610
rect 151560 679370 151650 679610
rect 151890 679370 152000 679610
rect 152240 679370 152330 679610
rect 152570 679370 152660 679610
rect 152900 679370 152990 679610
rect 153230 679370 153340 679610
rect 153580 679370 153670 679610
rect 153910 679370 154000 679610
rect 154240 679370 154330 679610
rect 154570 679370 154680 679610
rect 154920 679370 155010 679610
rect 155250 679370 155340 679610
rect 155580 679370 155670 679610
rect 155910 679370 155930 679610
rect 144930 679260 155930 679370
rect 144930 679020 144950 679260
rect 145190 679020 145300 679260
rect 145540 679020 145630 679260
rect 145870 679020 145960 679260
rect 146200 679020 146290 679260
rect 146530 679020 146640 679260
rect 146880 679020 146970 679260
rect 147210 679020 147300 679260
rect 147540 679020 147630 679260
rect 147870 679020 147980 679260
rect 148220 679020 148310 679260
rect 148550 679020 148640 679260
rect 148880 679020 148970 679260
rect 149210 679020 149320 679260
rect 149560 679020 149650 679260
rect 149890 679020 149980 679260
rect 150220 679020 150310 679260
rect 150550 679020 150660 679260
rect 150900 679020 150990 679260
rect 151230 679020 151320 679260
rect 151560 679020 151650 679260
rect 151890 679020 152000 679260
rect 152240 679020 152330 679260
rect 152570 679020 152660 679260
rect 152900 679020 152990 679260
rect 153230 679020 153340 679260
rect 153580 679020 153670 679260
rect 153910 679020 154000 679260
rect 154240 679020 154330 679260
rect 154570 679020 154680 679260
rect 154920 679020 155010 679260
rect 155250 679020 155340 679260
rect 155580 679020 155670 679260
rect 155910 679020 155930 679260
rect 144930 678930 155930 679020
rect 144930 678690 144950 678930
rect 145190 678690 145300 678930
rect 145540 678690 145630 678930
rect 145870 678690 145960 678930
rect 146200 678690 146290 678930
rect 146530 678690 146640 678930
rect 146880 678690 146970 678930
rect 147210 678690 147300 678930
rect 147540 678690 147630 678930
rect 147870 678690 147980 678930
rect 148220 678690 148310 678930
rect 148550 678690 148640 678930
rect 148880 678690 148970 678930
rect 149210 678690 149320 678930
rect 149560 678690 149650 678930
rect 149890 678690 149980 678930
rect 150220 678690 150310 678930
rect 150550 678690 150660 678930
rect 150900 678690 150990 678930
rect 151230 678690 151320 678930
rect 151560 678690 151650 678930
rect 151890 678690 152000 678930
rect 152240 678690 152330 678930
rect 152570 678690 152660 678930
rect 152900 678690 152990 678930
rect 153230 678690 153340 678930
rect 153580 678690 153670 678930
rect 153910 678690 154000 678930
rect 154240 678690 154330 678930
rect 154570 678690 154680 678930
rect 154920 678690 155010 678930
rect 155250 678690 155340 678930
rect 155580 678690 155670 678930
rect 155910 678690 155930 678930
rect 144930 678600 155930 678690
rect 144930 678360 144950 678600
rect 145190 678360 145300 678600
rect 145540 678360 145630 678600
rect 145870 678360 145960 678600
rect 146200 678360 146290 678600
rect 146530 678360 146640 678600
rect 146880 678360 146970 678600
rect 147210 678360 147300 678600
rect 147540 678360 147630 678600
rect 147870 678360 147980 678600
rect 148220 678360 148310 678600
rect 148550 678360 148640 678600
rect 148880 678360 148970 678600
rect 149210 678360 149320 678600
rect 149560 678360 149650 678600
rect 149890 678360 149980 678600
rect 150220 678360 150310 678600
rect 150550 678360 150660 678600
rect 150900 678360 150990 678600
rect 151230 678360 151320 678600
rect 151560 678360 151650 678600
rect 151890 678360 152000 678600
rect 152240 678360 152330 678600
rect 152570 678360 152660 678600
rect 152900 678360 152990 678600
rect 153230 678360 153340 678600
rect 153580 678360 153670 678600
rect 153910 678360 154000 678600
rect 154240 678360 154330 678600
rect 154570 678360 154680 678600
rect 154920 678360 155010 678600
rect 155250 678360 155340 678600
rect 155580 678360 155670 678600
rect 155910 678360 155930 678600
rect 144930 678270 155930 678360
rect 144930 678030 144950 678270
rect 145190 678030 145300 678270
rect 145540 678030 145630 678270
rect 145870 678030 145960 678270
rect 146200 678030 146290 678270
rect 146530 678030 146640 678270
rect 146880 678030 146970 678270
rect 147210 678030 147300 678270
rect 147540 678030 147630 678270
rect 147870 678030 147980 678270
rect 148220 678030 148310 678270
rect 148550 678030 148640 678270
rect 148880 678030 148970 678270
rect 149210 678030 149320 678270
rect 149560 678030 149650 678270
rect 149890 678030 149980 678270
rect 150220 678030 150310 678270
rect 150550 678030 150660 678270
rect 150900 678030 150990 678270
rect 151230 678030 151320 678270
rect 151560 678030 151650 678270
rect 151890 678030 152000 678270
rect 152240 678030 152330 678270
rect 152570 678030 152660 678270
rect 152900 678030 152990 678270
rect 153230 678030 153340 678270
rect 153580 678030 153670 678270
rect 153910 678030 154000 678270
rect 154240 678030 154330 678270
rect 154570 678030 154680 678270
rect 154920 678030 155010 678270
rect 155250 678030 155340 678270
rect 155580 678030 155670 678270
rect 155910 678030 155930 678270
rect 144930 677920 155930 678030
rect 144930 677680 144950 677920
rect 145190 677680 145300 677920
rect 145540 677680 145630 677920
rect 145870 677680 145960 677920
rect 146200 677680 146290 677920
rect 146530 677680 146640 677920
rect 146880 677680 146970 677920
rect 147210 677680 147300 677920
rect 147540 677680 147630 677920
rect 147870 677680 147980 677920
rect 148220 677680 148310 677920
rect 148550 677680 148640 677920
rect 148880 677680 148970 677920
rect 149210 677680 149320 677920
rect 149560 677680 149650 677920
rect 149890 677680 149980 677920
rect 150220 677680 150310 677920
rect 150550 677680 150660 677920
rect 150900 677680 150990 677920
rect 151230 677680 151320 677920
rect 151560 677680 151650 677920
rect 151890 677680 152000 677920
rect 152240 677680 152330 677920
rect 152570 677680 152660 677920
rect 152900 677680 152990 677920
rect 153230 677680 153340 677920
rect 153580 677680 153670 677920
rect 153910 677680 154000 677920
rect 154240 677680 154330 677920
rect 154570 677680 154680 677920
rect 154920 677680 155010 677920
rect 155250 677680 155340 677920
rect 155580 677680 155670 677920
rect 155910 677680 155930 677920
rect 144930 677590 155930 677680
rect 144930 677350 144950 677590
rect 145190 677350 145300 677590
rect 145540 677350 145630 677590
rect 145870 677350 145960 677590
rect 146200 677350 146290 677590
rect 146530 677350 146640 677590
rect 146880 677350 146970 677590
rect 147210 677350 147300 677590
rect 147540 677350 147630 677590
rect 147870 677350 147980 677590
rect 148220 677350 148310 677590
rect 148550 677350 148640 677590
rect 148880 677350 148970 677590
rect 149210 677350 149320 677590
rect 149560 677350 149650 677590
rect 149890 677350 149980 677590
rect 150220 677350 150310 677590
rect 150550 677350 150660 677590
rect 150900 677350 150990 677590
rect 151230 677350 151320 677590
rect 151560 677350 151650 677590
rect 151890 677350 152000 677590
rect 152240 677350 152330 677590
rect 152570 677350 152660 677590
rect 152900 677350 152990 677590
rect 153230 677350 153340 677590
rect 153580 677350 153670 677590
rect 153910 677350 154000 677590
rect 154240 677350 154330 677590
rect 154570 677350 154680 677590
rect 154920 677350 155010 677590
rect 155250 677350 155340 677590
rect 155580 677350 155670 677590
rect 155910 677350 155930 677590
rect 144930 677260 155930 677350
rect 144930 677020 144950 677260
rect 145190 677020 145300 677260
rect 145540 677020 145630 677260
rect 145870 677020 145960 677260
rect 146200 677020 146290 677260
rect 146530 677020 146640 677260
rect 146880 677020 146970 677260
rect 147210 677020 147300 677260
rect 147540 677020 147630 677260
rect 147870 677020 147980 677260
rect 148220 677020 148310 677260
rect 148550 677020 148640 677260
rect 148880 677020 148970 677260
rect 149210 677020 149320 677260
rect 149560 677020 149650 677260
rect 149890 677020 149980 677260
rect 150220 677020 150310 677260
rect 150550 677020 150660 677260
rect 150900 677020 150990 677260
rect 151230 677020 151320 677260
rect 151560 677020 151650 677260
rect 151890 677020 152000 677260
rect 152240 677020 152330 677260
rect 152570 677020 152660 677260
rect 152900 677020 152990 677260
rect 153230 677020 153340 677260
rect 153580 677020 153670 677260
rect 153910 677020 154000 677260
rect 154240 677020 154330 677260
rect 154570 677020 154680 677260
rect 154920 677020 155010 677260
rect 155250 677020 155340 677260
rect 155580 677020 155670 677260
rect 155910 677020 155930 677260
rect 144930 676930 155930 677020
rect 144930 676690 144950 676930
rect 145190 676690 145300 676930
rect 145540 676690 145630 676930
rect 145870 676690 145960 676930
rect 146200 676690 146290 676930
rect 146530 676690 146640 676930
rect 146880 676690 146970 676930
rect 147210 676690 147300 676930
rect 147540 676690 147630 676930
rect 147870 676690 147980 676930
rect 148220 676690 148310 676930
rect 148550 676690 148640 676930
rect 148880 676690 148970 676930
rect 149210 676690 149320 676930
rect 149560 676690 149650 676930
rect 149890 676690 149980 676930
rect 150220 676690 150310 676930
rect 150550 676690 150660 676930
rect 150900 676690 150990 676930
rect 151230 676690 151320 676930
rect 151560 676690 151650 676930
rect 151890 676690 152000 676930
rect 152240 676690 152330 676930
rect 152570 676690 152660 676930
rect 152900 676690 152990 676930
rect 153230 676690 153340 676930
rect 153580 676690 153670 676930
rect 153910 676690 154000 676930
rect 154240 676690 154330 676930
rect 154570 676690 154680 676930
rect 154920 676690 155010 676930
rect 155250 676690 155340 676930
rect 155580 676690 155670 676930
rect 155910 676690 155930 676930
rect 144930 676580 155930 676690
rect 144930 676340 144950 676580
rect 145190 676340 145300 676580
rect 145540 676340 145630 676580
rect 145870 676340 145960 676580
rect 146200 676340 146290 676580
rect 146530 676340 146640 676580
rect 146880 676340 146970 676580
rect 147210 676340 147300 676580
rect 147540 676340 147630 676580
rect 147870 676340 147980 676580
rect 148220 676340 148310 676580
rect 148550 676340 148640 676580
rect 148880 676340 148970 676580
rect 149210 676340 149320 676580
rect 149560 676340 149650 676580
rect 149890 676340 149980 676580
rect 150220 676340 150310 676580
rect 150550 676340 150660 676580
rect 150900 676340 150990 676580
rect 151230 676340 151320 676580
rect 151560 676340 151650 676580
rect 151890 676340 152000 676580
rect 152240 676340 152330 676580
rect 152570 676340 152660 676580
rect 152900 676340 152990 676580
rect 153230 676340 153340 676580
rect 153580 676340 153670 676580
rect 153910 676340 154000 676580
rect 154240 676340 154330 676580
rect 154570 676340 154680 676580
rect 154920 676340 155010 676580
rect 155250 676340 155340 676580
rect 155580 676340 155670 676580
rect 155910 676340 155930 676580
rect 144930 676250 155930 676340
rect 144930 676010 144950 676250
rect 145190 676010 145300 676250
rect 145540 676010 145630 676250
rect 145870 676010 145960 676250
rect 146200 676010 146290 676250
rect 146530 676010 146640 676250
rect 146880 676010 146970 676250
rect 147210 676010 147300 676250
rect 147540 676010 147630 676250
rect 147870 676010 147980 676250
rect 148220 676010 148310 676250
rect 148550 676010 148640 676250
rect 148880 676010 148970 676250
rect 149210 676010 149320 676250
rect 149560 676010 149650 676250
rect 149890 676010 149980 676250
rect 150220 676010 150310 676250
rect 150550 676010 150660 676250
rect 150900 676010 150990 676250
rect 151230 676010 151320 676250
rect 151560 676010 151650 676250
rect 151890 676010 152000 676250
rect 152240 676010 152330 676250
rect 152570 676010 152660 676250
rect 152900 676010 152990 676250
rect 153230 676010 153340 676250
rect 153580 676010 153670 676250
rect 153910 676010 154000 676250
rect 154240 676010 154330 676250
rect 154570 676010 154680 676250
rect 154920 676010 155010 676250
rect 155250 676010 155340 676250
rect 155580 676010 155670 676250
rect 155910 676010 155930 676250
rect 144930 675920 155930 676010
rect 144930 675680 144950 675920
rect 145190 675680 145300 675920
rect 145540 675680 145630 675920
rect 145870 675680 145960 675920
rect 146200 675680 146290 675920
rect 146530 675680 146640 675920
rect 146880 675680 146970 675920
rect 147210 675680 147300 675920
rect 147540 675680 147630 675920
rect 147870 675680 147980 675920
rect 148220 675680 148310 675920
rect 148550 675680 148640 675920
rect 148880 675680 148970 675920
rect 149210 675680 149320 675920
rect 149560 675680 149650 675920
rect 149890 675680 149980 675920
rect 150220 675680 150310 675920
rect 150550 675680 150660 675920
rect 150900 675680 150990 675920
rect 151230 675680 151320 675920
rect 151560 675680 151650 675920
rect 151890 675680 152000 675920
rect 152240 675680 152330 675920
rect 152570 675680 152660 675920
rect 152900 675680 152990 675920
rect 153230 675680 153340 675920
rect 153580 675680 153670 675920
rect 153910 675680 154000 675920
rect 154240 675680 154330 675920
rect 154570 675680 154680 675920
rect 154920 675680 155010 675920
rect 155250 675680 155340 675920
rect 155580 675680 155670 675920
rect 155910 675680 155930 675920
rect 144930 675590 155930 675680
rect 144930 675350 144950 675590
rect 145190 675350 145300 675590
rect 145540 675350 145630 675590
rect 145870 675350 145960 675590
rect 146200 675350 146290 675590
rect 146530 675350 146640 675590
rect 146880 675350 146970 675590
rect 147210 675350 147300 675590
rect 147540 675350 147630 675590
rect 147870 675350 147980 675590
rect 148220 675350 148310 675590
rect 148550 675350 148640 675590
rect 148880 675350 148970 675590
rect 149210 675350 149320 675590
rect 149560 675350 149650 675590
rect 149890 675350 149980 675590
rect 150220 675350 150310 675590
rect 150550 675350 150660 675590
rect 150900 675350 150990 675590
rect 151230 675350 151320 675590
rect 151560 675350 151650 675590
rect 151890 675350 152000 675590
rect 152240 675350 152330 675590
rect 152570 675350 152660 675590
rect 152900 675350 152990 675590
rect 153230 675350 153340 675590
rect 153580 675350 153670 675590
rect 153910 675350 154000 675590
rect 154240 675350 154330 675590
rect 154570 675350 154680 675590
rect 154920 675350 155010 675590
rect 155250 675350 155340 675590
rect 155580 675350 155670 675590
rect 155910 675350 155930 675590
rect 144930 675240 155930 675350
rect 144930 675000 144950 675240
rect 145190 675000 145300 675240
rect 145540 675000 145630 675240
rect 145870 675000 145960 675240
rect 146200 675000 146290 675240
rect 146530 675000 146640 675240
rect 146880 675000 146970 675240
rect 147210 675000 147300 675240
rect 147540 675000 147630 675240
rect 147870 675000 147980 675240
rect 148220 675000 148310 675240
rect 148550 675000 148640 675240
rect 148880 675000 148970 675240
rect 149210 675000 149320 675240
rect 149560 675000 149650 675240
rect 149890 675000 149980 675240
rect 150220 675000 150310 675240
rect 150550 675000 150660 675240
rect 150900 675000 150990 675240
rect 151230 675000 151320 675240
rect 151560 675000 151650 675240
rect 151890 675000 152000 675240
rect 152240 675000 152330 675240
rect 152570 675000 152660 675240
rect 152900 675000 152990 675240
rect 153230 675000 153340 675240
rect 153580 675000 153670 675240
rect 153910 675000 154000 675240
rect 154240 675000 154330 675240
rect 154570 675000 154680 675240
rect 154920 675000 155010 675240
rect 155250 675000 155340 675240
rect 155580 675000 155670 675240
rect 155910 675000 155930 675240
rect 144930 674910 155930 675000
rect 144930 674670 144950 674910
rect 145190 674670 145300 674910
rect 145540 674670 145630 674910
rect 145870 674670 145960 674910
rect 146200 674670 146290 674910
rect 146530 674670 146640 674910
rect 146880 674670 146970 674910
rect 147210 674670 147300 674910
rect 147540 674670 147630 674910
rect 147870 674670 147980 674910
rect 148220 674670 148310 674910
rect 148550 674670 148640 674910
rect 148880 674670 148970 674910
rect 149210 674670 149320 674910
rect 149560 674670 149650 674910
rect 149890 674670 149980 674910
rect 150220 674670 150310 674910
rect 150550 674670 150660 674910
rect 150900 674670 150990 674910
rect 151230 674670 151320 674910
rect 151560 674670 151650 674910
rect 151890 674670 152000 674910
rect 152240 674670 152330 674910
rect 152570 674670 152660 674910
rect 152900 674670 152990 674910
rect 153230 674670 153340 674910
rect 153580 674670 153670 674910
rect 153910 674670 154000 674910
rect 154240 674670 154330 674910
rect 154570 674670 154680 674910
rect 154920 674670 155010 674910
rect 155250 674670 155340 674910
rect 155580 674670 155670 674910
rect 155910 674670 155930 674910
rect 144930 674580 155930 674670
rect 144930 674340 144950 674580
rect 145190 674340 145300 674580
rect 145540 674340 145630 674580
rect 145870 674340 145960 674580
rect 146200 674340 146290 674580
rect 146530 674340 146640 674580
rect 146880 674340 146970 674580
rect 147210 674340 147300 674580
rect 147540 674340 147630 674580
rect 147870 674340 147980 674580
rect 148220 674340 148310 674580
rect 148550 674340 148640 674580
rect 148880 674340 148970 674580
rect 149210 674340 149320 674580
rect 149560 674340 149650 674580
rect 149890 674340 149980 674580
rect 150220 674340 150310 674580
rect 150550 674340 150660 674580
rect 150900 674340 150990 674580
rect 151230 674340 151320 674580
rect 151560 674340 151650 674580
rect 151890 674340 152000 674580
rect 152240 674340 152330 674580
rect 152570 674340 152660 674580
rect 152900 674340 152990 674580
rect 153230 674340 153340 674580
rect 153580 674340 153670 674580
rect 153910 674340 154000 674580
rect 154240 674340 154330 674580
rect 154570 674340 154680 674580
rect 154920 674340 155010 674580
rect 155250 674340 155340 674580
rect 155580 674340 155670 674580
rect 155910 674340 155930 674580
rect 144930 674250 155930 674340
rect 144930 674010 144950 674250
rect 145190 674010 145300 674250
rect 145540 674010 145630 674250
rect 145870 674010 145960 674250
rect 146200 674010 146290 674250
rect 146530 674010 146640 674250
rect 146880 674010 146970 674250
rect 147210 674010 147300 674250
rect 147540 674010 147630 674250
rect 147870 674010 147980 674250
rect 148220 674010 148310 674250
rect 148550 674010 148640 674250
rect 148880 674010 148970 674250
rect 149210 674010 149320 674250
rect 149560 674010 149650 674250
rect 149890 674010 149980 674250
rect 150220 674010 150310 674250
rect 150550 674010 150660 674250
rect 150900 674010 150990 674250
rect 151230 674010 151320 674250
rect 151560 674010 151650 674250
rect 151890 674010 152000 674250
rect 152240 674010 152330 674250
rect 152570 674010 152660 674250
rect 152900 674010 152990 674250
rect 153230 674010 153340 674250
rect 153580 674010 153670 674250
rect 153910 674010 154000 674250
rect 154240 674010 154330 674250
rect 154570 674010 154680 674250
rect 154920 674010 155010 674250
rect 155250 674010 155340 674250
rect 155580 674010 155670 674250
rect 155910 674010 155930 674250
rect 144930 673900 155930 674010
rect 144930 673660 144950 673900
rect 145190 673660 145300 673900
rect 145540 673660 145630 673900
rect 145870 673660 145960 673900
rect 146200 673660 146290 673900
rect 146530 673660 146640 673900
rect 146880 673660 146970 673900
rect 147210 673660 147300 673900
rect 147540 673660 147630 673900
rect 147870 673660 147980 673900
rect 148220 673660 148310 673900
rect 148550 673660 148640 673900
rect 148880 673660 148970 673900
rect 149210 673660 149320 673900
rect 149560 673660 149650 673900
rect 149890 673660 149980 673900
rect 150220 673660 150310 673900
rect 150550 673660 150660 673900
rect 150900 673660 150990 673900
rect 151230 673660 151320 673900
rect 151560 673660 151650 673900
rect 151890 673660 152000 673900
rect 152240 673660 152330 673900
rect 152570 673660 152660 673900
rect 152900 673660 152990 673900
rect 153230 673660 153340 673900
rect 153580 673660 153670 673900
rect 153910 673660 154000 673900
rect 154240 673660 154330 673900
rect 154570 673660 154680 673900
rect 154920 673660 155010 673900
rect 155250 673660 155340 673900
rect 155580 673660 155670 673900
rect 155910 673660 155930 673900
rect 144930 673570 155930 673660
rect 144930 673330 144950 673570
rect 145190 673330 145300 673570
rect 145540 673330 145630 673570
rect 145870 673330 145960 673570
rect 146200 673330 146290 673570
rect 146530 673330 146640 673570
rect 146880 673330 146970 673570
rect 147210 673330 147300 673570
rect 147540 673330 147630 673570
rect 147870 673330 147980 673570
rect 148220 673330 148310 673570
rect 148550 673330 148640 673570
rect 148880 673330 148970 673570
rect 149210 673330 149320 673570
rect 149560 673330 149650 673570
rect 149890 673330 149980 673570
rect 150220 673330 150310 673570
rect 150550 673330 150660 673570
rect 150900 673330 150990 673570
rect 151230 673330 151320 673570
rect 151560 673330 151650 673570
rect 151890 673330 152000 673570
rect 152240 673330 152330 673570
rect 152570 673330 152660 673570
rect 152900 673330 152990 673570
rect 153230 673330 153340 673570
rect 153580 673330 153670 673570
rect 153910 673330 154000 673570
rect 154240 673330 154330 673570
rect 154570 673330 154680 673570
rect 154920 673330 155010 673570
rect 155250 673330 155340 673570
rect 155580 673330 155670 673570
rect 155910 673330 155930 673570
rect 144930 673240 155930 673330
rect 144930 673000 144950 673240
rect 145190 673000 145300 673240
rect 145540 673000 145630 673240
rect 145870 673000 145960 673240
rect 146200 673000 146290 673240
rect 146530 673000 146640 673240
rect 146880 673000 146970 673240
rect 147210 673000 147300 673240
rect 147540 673000 147630 673240
rect 147870 673000 147980 673240
rect 148220 673000 148310 673240
rect 148550 673000 148640 673240
rect 148880 673000 148970 673240
rect 149210 673000 149320 673240
rect 149560 673000 149650 673240
rect 149890 673000 149980 673240
rect 150220 673000 150310 673240
rect 150550 673000 150660 673240
rect 150900 673000 150990 673240
rect 151230 673000 151320 673240
rect 151560 673000 151650 673240
rect 151890 673000 152000 673240
rect 152240 673000 152330 673240
rect 152570 673000 152660 673240
rect 152900 673000 152990 673240
rect 153230 673000 153340 673240
rect 153580 673000 153670 673240
rect 153910 673000 154000 673240
rect 154240 673000 154330 673240
rect 154570 673000 154680 673240
rect 154920 673000 155010 673240
rect 155250 673000 155340 673240
rect 155580 673000 155670 673240
rect 155910 673000 155930 673240
rect 144930 672910 155930 673000
rect 144930 672670 144950 672910
rect 145190 672670 145300 672910
rect 145540 672670 145630 672910
rect 145870 672670 145960 672910
rect 146200 672670 146290 672910
rect 146530 672670 146640 672910
rect 146880 672670 146970 672910
rect 147210 672670 147300 672910
rect 147540 672670 147630 672910
rect 147870 672670 147980 672910
rect 148220 672670 148310 672910
rect 148550 672670 148640 672910
rect 148880 672670 148970 672910
rect 149210 672670 149320 672910
rect 149560 672670 149650 672910
rect 149890 672670 149980 672910
rect 150220 672670 150310 672910
rect 150550 672670 150660 672910
rect 150900 672670 150990 672910
rect 151230 672670 151320 672910
rect 151560 672670 151650 672910
rect 151890 672670 152000 672910
rect 152240 672670 152330 672910
rect 152570 672670 152660 672910
rect 152900 672670 152990 672910
rect 153230 672670 153340 672910
rect 153580 672670 153670 672910
rect 153910 672670 154000 672910
rect 154240 672670 154330 672910
rect 154570 672670 154680 672910
rect 154920 672670 155010 672910
rect 155250 672670 155340 672910
rect 155580 672670 155670 672910
rect 155910 672670 155930 672910
rect 144930 672560 155930 672670
rect 144930 672320 144950 672560
rect 145190 672320 145300 672560
rect 145540 672320 145630 672560
rect 145870 672320 145960 672560
rect 146200 672320 146290 672560
rect 146530 672320 146640 672560
rect 146880 672320 146970 672560
rect 147210 672320 147300 672560
rect 147540 672320 147630 672560
rect 147870 672320 147980 672560
rect 148220 672320 148310 672560
rect 148550 672320 148640 672560
rect 148880 672320 148970 672560
rect 149210 672320 149320 672560
rect 149560 672320 149650 672560
rect 149890 672320 149980 672560
rect 150220 672320 150310 672560
rect 150550 672320 150660 672560
rect 150900 672320 150990 672560
rect 151230 672320 151320 672560
rect 151560 672320 151650 672560
rect 151890 672320 152000 672560
rect 152240 672320 152330 672560
rect 152570 672320 152660 672560
rect 152900 672320 152990 672560
rect 153230 672320 153340 672560
rect 153580 672320 153670 672560
rect 153910 672320 154000 672560
rect 154240 672320 154330 672560
rect 154570 672320 154680 672560
rect 154920 672320 155010 672560
rect 155250 672320 155340 672560
rect 155580 672320 155670 672560
rect 155910 672320 155930 672560
rect 144930 672300 155930 672320
rect 110790 671900 121790 671920
rect 110790 671660 110810 671900
rect 111050 671660 111140 671900
rect 111380 671660 111470 671900
rect 111710 671660 111800 671900
rect 112040 671660 112150 671900
rect 112390 671660 112480 671900
rect 112720 671660 112810 671900
rect 113050 671660 113140 671900
rect 113380 671660 113490 671900
rect 113730 671660 113820 671900
rect 114060 671660 114150 671900
rect 114390 671660 114480 671900
rect 114720 671660 114830 671900
rect 115070 671660 115160 671900
rect 115400 671660 115490 671900
rect 115730 671660 115820 671900
rect 116060 671660 116170 671900
rect 116410 671660 116500 671900
rect 116740 671660 116830 671900
rect 117070 671660 117160 671900
rect 117400 671660 117510 671900
rect 117750 671660 117840 671900
rect 118080 671660 118170 671900
rect 118410 671660 118500 671900
rect 118740 671660 118850 671900
rect 119090 671660 119180 671900
rect 119420 671660 119510 671900
rect 119750 671660 119840 671900
rect 120080 671660 120190 671900
rect 120430 671660 120520 671900
rect 120760 671660 120850 671900
rect 121090 671660 121180 671900
rect 121420 671660 121530 671900
rect 121770 671660 121790 671900
rect 110790 671550 121790 671660
rect 110790 671310 110810 671550
rect 111050 671310 111140 671550
rect 111380 671310 111470 671550
rect 111710 671310 111800 671550
rect 112040 671310 112150 671550
rect 112390 671310 112480 671550
rect 112720 671310 112810 671550
rect 113050 671310 113140 671550
rect 113380 671310 113490 671550
rect 113730 671310 113820 671550
rect 114060 671310 114150 671550
rect 114390 671310 114480 671550
rect 114720 671310 114830 671550
rect 115070 671310 115160 671550
rect 115400 671310 115490 671550
rect 115730 671310 115820 671550
rect 116060 671310 116170 671550
rect 116410 671310 116500 671550
rect 116740 671310 116830 671550
rect 117070 671310 117160 671550
rect 117400 671310 117510 671550
rect 117750 671310 117840 671550
rect 118080 671310 118170 671550
rect 118410 671310 118500 671550
rect 118740 671310 118850 671550
rect 119090 671310 119180 671550
rect 119420 671310 119510 671550
rect 119750 671310 119840 671550
rect 120080 671310 120190 671550
rect 120430 671310 120520 671550
rect 120760 671310 120850 671550
rect 121090 671310 121180 671550
rect 121420 671310 121530 671550
rect 121770 671310 121790 671550
rect 110790 671220 121790 671310
rect 110790 670980 110810 671220
rect 111050 670980 111140 671220
rect 111380 670980 111470 671220
rect 111710 670980 111800 671220
rect 112040 670980 112150 671220
rect 112390 670980 112480 671220
rect 112720 670980 112810 671220
rect 113050 670980 113140 671220
rect 113380 670980 113490 671220
rect 113730 670980 113820 671220
rect 114060 670980 114150 671220
rect 114390 670980 114480 671220
rect 114720 670980 114830 671220
rect 115070 670980 115160 671220
rect 115400 670980 115490 671220
rect 115730 670980 115820 671220
rect 116060 670980 116170 671220
rect 116410 670980 116500 671220
rect 116740 670980 116830 671220
rect 117070 670980 117160 671220
rect 117400 670980 117510 671220
rect 117750 670980 117840 671220
rect 118080 670980 118170 671220
rect 118410 670980 118500 671220
rect 118740 670980 118850 671220
rect 119090 670980 119180 671220
rect 119420 670980 119510 671220
rect 119750 670980 119840 671220
rect 120080 670980 120190 671220
rect 120430 670980 120520 671220
rect 120760 670980 120850 671220
rect 121090 670980 121180 671220
rect 121420 670980 121530 671220
rect 121770 670980 121790 671220
rect 110790 670890 121790 670980
rect 110790 670650 110810 670890
rect 111050 670650 111140 670890
rect 111380 670650 111470 670890
rect 111710 670650 111800 670890
rect 112040 670650 112150 670890
rect 112390 670650 112480 670890
rect 112720 670650 112810 670890
rect 113050 670650 113140 670890
rect 113380 670650 113490 670890
rect 113730 670650 113820 670890
rect 114060 670650 114150 670890
rect 114390 670650 114480 670890
rect 114720 670650 114830 670890
rect 115070 670650 115160 670890
rect 115400 670650 115490 670890
rect 115730 670650 115820 670890
rect 116060 670650 116170 670890
rect 116410 670650 116500 670890
rect 116740 670650 116830 670890
rect 117070 670650 117160 670890
rect 117400 670650 117510 670890
rect 117750 670650 117840 670890
rect 118080 670650 118170 670890
rect 118410 670650 118500 670890
rect 118740 670650 118850 670890
rect 119090 670650 119180 670890
rect 119420 670650 119510 670890
rect 119750 670650 119840 670890
rect 120080 670650 120190 670890
rect 120430 670650 120520 670890
rect 120760 670650 120850 670890
rect 121090 670650 121180 670890
rect 121420 670650 121530 670890
rect 121770 670650 121790 670890
rect 110790 670560 121790 670650
rect 110790 670320 110810 670560
rect 111050 670320 111140 670560
rect 111380 670320 111470 670560
rect 111710 670320 111800 670560
rect 112040 670320 112150 670560
rect 112390 670320 112480 670560
rect 112720 670320 112810 670560
rect 113050 670320 113140 670560
rect 113380 670320 113490 670560
rect 113730 670320 113820 670560
rect 114060 670320 114150 670560
rect 114390 670320 114480 670560
rect 114720 670320 114830 670560
rect 115070 670320 115160 670560
rect 115400 670320 115490 670560
rect 115730 670320 115820 670560
rect 116060 670320 116170 670560
rect 116410 670320 116500 670560
rect 116740 670320 116830 670560
rect 117070 670320 117160 670560
rect 117400 670320 117510 670560
rect 117750 670320 117840 670560
rect 118080 670320 118170 670560
rect 118410 670320 118500 670560
rect 118740 670320 118850 670560
rect 119090 670320 119180 670560
rect 119420 670320 119510 670560
rect 119750 670320 119840 670560
rect 120080 670320 120190 670560
rect 120430 670320 120520 670560
rect 120760 670320 120850 670560
rect 121090 670320 121180 670560
rect 121420 670320 121530 670560
rect 121770 670320 121790 670560
rect 110790 670210 121790 670320
rect 110790 669970 110810 670210
rect 111050 669970 111140 670210
rect 111380 669970 111470 670210
rect 111710 669970 111800 670210
rect 112040 669970 112150 670210
rect 112390 669970 112480 670210
rect 112720 669970 112810 670210
rect 113050 669970 113140 670210
rect 113380 669970 113490 670210
rect 113730 669970 113820 670210
rect 114060 669970 114150 670210
rect 114390 669970 114480 670210
rect 114720 669970 114830 670210
rect 115070 669970 115160 670210
rect 115400 669970 115490 670210
rect 115730 669970 115820 670210
rect 116060 669970 116170 670210
rect 116410 669970 116500 670210
rect 116740 669970 116830 670210
rect 117070 669970 117160 670210
rect 117400 669970 117510 670210
rect 117750 669970 117840 670210
rect 118080 669970 118170 670210
rect 118410 669970 118500 670210
rect 118740 669970 118850 670210
rect 119090 669970 119180 670210
rect 119420 669970 119510 670210
rect 119750 669970 119840 670210
rect 120080 669970 120190 670210
rect 120430 669970 120520 670210
rect 120760 669970 120850 670210
rect 121090 669970 121180 670210
rect 121420 669970 121530 670210
rect 121770 669970 121790 670210
rect 110790 669880 121790 669970
rect 110790 669640 110810 669880
rect 111050 669640 111140 669880
rect 111380 669640 111470 669880
rect 111710 669640 111800 669880
rect 112040 669640 112150 669880
rect 112390 669640 112480 669880
rect 112720 669640 112810 669880
rect 113050 669640 113140 669880
rect 113380 669640 113490 669880
rect 113730 669640 113820 669880
rect 114060 669640 114150 669880
rect 114390 669640 114480 669880
rect 114720 669640 114830 669880
rect 115070 669640 115160 669880
rect 115400 669640 115490 669880
rect 115730 669640 115820 669880
rect 116060 669640 116170 669880
rect 116410 669640 116500 669880
rect 116740 669640 116830 669880
rect 117070 669640 117160 669880
rect 117400 669640 117510 669880
rect 117750 669640 117840 669880
rect 118080 669640 118170 669880
rect 118410 669640 118500 669880
rect 118740 669640 118850 669880
rect 119090 669640 119180 669880
rect 119420 669640 119510 669880
rect 119750 669640 119840 669880
rect 120080 669640 120190 669880
rect 120430 669640 120520 669880
rect 120760 669640 120850 669880
rect 121090 669640 121180 669880
rect 121420 669640 121530 669880
rect 121770 669640 121790 669880
rect 110790 669550 121790 669640
rect 110790 669310 110810 669550
rect 111050 669310 111140 669550
rect 111380 669310 111470 669550
rect 111710 669310 111800 669550
rect 112040 669310 112150 669550
rect 112390 669310 112480 669550
rect 112720 669310 112810 669550
rect 113050 669310 113140 669550
rect 113380 669310 113490 669550
rect 113730 669310 113820 669550
rect 114060 669310 114150 669550
rect 114390 669310 114480 669550
rect 114720 669310 114830 669550
rect 115070 669310 115160 669550
rect 115400 669310 115490 669550
rect 115730 669310 115820 669550
rect 116060 669310 116170 669550
rect 116410 669310 116500 669550
rect 116740 669310 116830 669550
rect 117070 669310 117160 669550
rect 117400 669310 117510 669550
rect 117750 669310 117840 669550
rect 118080 669310 118170 669550
rect 118410 669310 118500 669550
rect 118740 669310 118850 669550
rect 119090 669310 119180 669550
rect 119420 669310 119510 669550
rect 119750 669310 119840 669550
rect 120080 669310 120190 669550
rect 120430 669310 120520 669550
rect 120760 669310 120850 669550
rect 121090 669310 121180 669550
rect 121420 669310 121530 669550
rect 121770 669310 121790 669550
rect 110790 669220 121790 669310
rect 110790 668980 110810 669220
rect 111050 668980 111140 669220
rect 111380 668980 111470 669220
rect 111710 668980 111800 669220
rect 112040 668980 112150 669220
rect 112390 668980 112480 669220
rect 112720 668980 112810 669220
rect 113050 668980 113140 669220
rect 113380 668980 113490 669220
rect 113730 668980 113820 669220
rect 114060 668980 114150 669220
rect 114390 668980 114480 669220
rect 114720 668980 114830 669220
rect 115070 668980 115160 669220
rect 115400 668980 115490 669220
rect 115730 668980 115820 669220
rect 116060 668980 116170 669220
rect 116410 668980 116500 669220
rect 116740 668980 116830 669220
rect 117070 668980 117160 669220
rect 117400 668980 117510 669220
rect 117750 668980 117840 669220
rect 118080 668980 118170 669220
rect 118410 668980 118500 669220
rect 118740 668980 118850 669220
rect 119090 668980 119180 669220
rect 119420 668980 119510 669220
rect 119750 668980 119840 669220
rect 120080 668980 120190 669220
rect 120430 668980 120520 669220
rect 120760 668980 120850 669220
rect 121090 668980 121180 669220
rect 121420 668980 121530 669220
rect 121770 668980 121790 669220
rect 110790 668870 121790 668980
rect 110790 668630 110810 668870
rect 111050 668630 111140 668870
rect 111380 668630 111470 668870
rect 111710 668630 111800 668870
rect 112040 668630 112150 668870
rect 112390 668630 112480 668870
rect 112720 668630 112810 668870
rect 113050 668630 113140 668870
rect 113380 668630 113490 668870
rect 113730 668630 113820 668870
rect 114060 668630 114150 668870
rect 114390 668630 114480 668870
rect 114720 668630 114830 668870
rect 115070 668630 115160 668870
rect 115400 668630 115490 668870
rect 115730 668630 115820 668870
rect 116060 668630 116170 668870
rect 116410 668630 116500 668870
rect 116740 668630 116830 668870
rect 117070 668630 117160 668870
rect 117400 668630 117510 668870
rect 117750 668630 117840 668870
rect 118080 668630 118170 668870
rect 118410 668630 118500 668870
rect 118740 668630 118850 668870
rect 119090 668630 119180 668870
rect 119420 668630 119510 668870
rect 119750 668630 119840 668870
rect 120080 668630 120190 668870
rect 120430 668630 120520 668870
rect 120760 668630 120850 668870
rect 121090 668630 121180 668870
rect 121420 668630 121530 668870
rect 121770 668630 121790 668870
rect 110790 668540 121790 668630
rect 110790 668300 110810 668540
rect 111050 668300 111140 668540
rect 111380 668300 111470 668540
rect 111710 668300 111800 668540
rect 112040 668300 112150 668540
rect 112390 668300 112480 668540
rect 112720 668300 112810 668540
rect 113050 668300 113140 668540
rect 113380 668300 113490 668540
rect 113730 668300 113820 668540
rect 114060 668300 114150 668540
rect 114390 668300 114480 668540
rect 114720 668300 114830 668540
rect 115070 668300 115160 668540
rect 115400 668300 115490 668540
rect 115730 668300 115820 668540
rect 116060 668300 116170 668540
rect 116410 668300 116500 668540
rect 116740 668300 116830 668540
rect 117070 668300 117160 668540
rect 117400 668300 117510 668540
rect 117750 668300 117840 668540
rect 118080 668300 118170 668540
rect 118410 668300 118500 668540
rect 118740 668300 118850 668540
rect 119090 668300 119180 668540
rect 119420 668300 119510 668540
rect 119750 668300 119840 668540
rect 120080 668300 120190 668540
rect 120430 668300 120520 668540
rect 120760 668300 120850 668540
rect 121090 668300 121180 668540
rect 121420 668300 121530 668540
rect 121770 668300 121790 668540
rect 110790 668210 121790 668300
rect 110790 667970 110810 668210
rect 111050 667970 111140 668210
rect 111380 667970 111470 668210
rect 111710 667970 111800 668210
rect 112040 667970 112150 668210
rect 112390 667970 112480 668210
rect 112720 667970 112810 668210
rect 113050 667970 113140 668210
rect 113380 667970 113490 668210
rect 113730 667970 113820 668210
rect 114060 667970 114150 668210
rect 114390 667970 114480 668210
rect 114720 667970 114830 668210
rect 115070 667970 115160 668210
rect 115400 667970 115490 668210
rect 115730 667970 115820 668210
rect 116060 667970 116170 668210
rect 116410 667970 116500 668210
rect 116740 667970 116830 668210
rect 117070 667970 117160 668210
rect 117400 667970 117510 668210
rect 117750 667970 117840 668210
rect 118080 667970 118170 668210
rect 118410 667970 118500 668210
rect 118740 667970 118850 668210
rect 119090 667970 119180 668210
rect 119420 667970 119510 668210
rect 119750 667970 119840 668210
rect 120080 667970 120190 668210
rect 120430 667970 120520 668210
rect 120760 667970 120850 668210
rect 121090 667970 121180 668210
rect 121420 667970 121530 668210
rect 121770 667970 121790 668210
rect 110790 667880 121790 667970
rect 110790 667640 110810 667880
rect 111050 667640 111140 667880
rect 111380 667640 111470 667880
rect 111710 667640 111800 667880
rect 112040 667640 112150 667880
rect 112390 667640 112480 667880
rect 112720 667640 112810 667880
rect 113050 667640 113140 667880
rect 113380 667640 113490 667880
rect 113730 667640 113820 667880
rect 114060 667640 114150 667880
rect 114390 667640 114480 667880
rect 114720 667640 114830 667880
rect 115070 667640 115160 667880
rect 115400 667640 115490 667880
rect 115730 667640 115820 667880
rect 116060 667640 116170 667880
rect 116410 667640 116500 667880
rect 116740 667640 116830 667880
rect 117070 667640 117160 667880
rect 117400 667640 117510 667880
rect 117750 667640 117840 667880
rect 118080 667640 118170 667880
rect 118410 667640 118500 667880
rect 118740 667640 118850 667880
rect 119090 667640 119180 667880
rect 119420 667640 119510 667880
rect 119750 667640 119840 667880
rect 120080 667640 120190 667880
rect 120430 667640 120520 667880
rect 120760 667640 120850 667880
rect 121090 667640 121180 667880
rect 121420 667640 121530 667880
rect 121770 667640 121790 667880
rect 110790 667530 121790 667640
rect 110790 667290 110810 667530
rect 111050 667290 111140 667530
rect 111380 667290 111470 667530
rect 111710 667290 111800 667530
rect 112040 667290 112150 667530
rect 112390 667290 112480 667530
rect 112720 667290 112810 667530
rect 113050 667290 113140 667530
rect 113380 667290 113490 667530
rect 113730 667290 113820 667530
rect 114060 667290 114150 667530
rect 114390 667290 114480 667530
rect 114720 667290 114830 667530
rect 115070 667290 115160 667530
rect 115400 667290 115490 667530
rect 115730 667290 115820 667530
rect 116060 667290 116170 667530
rect 116410 667290 116500 667530
rect 116740 667290 116830 667530
rect 117070 667290 117160 667530
rect 117400 667290 117510 667530
rect 117750 667290 117840 667530
rect 118080 667290 118170 667530
rect 118410 667290 118500 667530
rect 118740 667290 118850 667530
rect 119090 667290 119180 667530
rect 119420 667290 119510 667530
rect 119750 667290 119840 667530
rect 120080 667290 120190 667530
rect 120430 667290 120520 667530
rect 120760 667290 120850 667530
rect 121090 667290 121180 667530
rect 121420 667290 121530 667530
rect 121770 667290 121790 667530
rect 110790 667200 121790 667290
rect 110790 666960 110810 667200
rect 111050 666960 111140 667200
rect 111380 666960 111470 667200
rect 111710 666960 111800 667200
rect 112040 666960 112150 667200
rect 112390 666960 112480 667200
rect 112720 666960 112810 667200
rect 113050 666960 113140 667200
rect 113380 666960 113490 667200
rect 113730 666960 113820 667200
rect 114060 666960 114150 667200
rect 114390 666960 114480 667200
rect 114720 666960 114830 667200
rect 115070 666960 115160 667200
rect 115400 666960 115490 667200
rect 115730 666960 115820 667200
rect 116060 666960 116170 667200
rect 116410 666960 116500 667200
rect 116740 666960 116830 667200
rect 117070 666960 117160 667200
rect 117400 666960 117510 667200
rect 117750 666960 117840 667200
rect 118080 666960 118170 667200
rect 118410 666960 118500 667200
rect 118740 666960 118850 667200
rect 119090 666960 119180 667200
rect 119420 666960 119510 667200
rect 119750 666960 119840 667200
rect 120080 666960 120190 667200
rect 120430 666960 120520 667200
rect 120760 666960 120850 667200
rect 121090 666960 121180 667200
rect 121420 666960 121530 667200
rect 121770 666960 121790 667200
rect 110790 666870 121790 666960
rect 110790 666630 110810 666870
rect 111050 666630 111140 666870
rect 111380 666630 111470 666870
rect 111710 666630 111800 666870
rect 112040 666630 112150 666870
rect 112390 666630 112480 666870
rect 112720 666630 112810 666870
rect 113050 666630 113140 666870
rect 113380 666630 113490 666870
rect 113730 666630 113820 666870
rect 114060 666630 114150 666870
rect 114390 666630 114480 666870
rect 114720 666630 114830 666870
rect 115070 666630 115160 666870
rect 115400 666630 115490 666870
rect 115730 666630 115820 666870
rect 116060 666630 116170 666870
rect 116410 666630 116500 666870
rect 116740 666630 116830 666870
rect 117070 666630 117160 666870
rect 117400 666630 117510 666870
rect 117750 666630 117840 666870
rect 118080 666630 118170 666870
rect 118410 666630 118500 666870
rect 118740 666630 118850 666870
rect 119090 666630 119180 666870
rect 119420 666630 119510 666870
rect 119750 666630 119840 666870
rect 120080 666630 120190 666870
rect 120430 666630 120520 666870
rect 120760 666630 120850 666870
rect 121090 666630 121180 666870
rect 121420 666630 121530 666870
rect 121770 666630 121790 666870
rect 110790 666540 121790 666630
rect 110790 666300 110810 666540
rect 111050 666300 111140 666540
rect 111380 666300 111470 666540
rect 111710 666300 111800 666540
rect 112040 666300 112150 666540
rect 112390 666300 112480 666540
rect 112720 666300 112810 666540
rect 113050 666300 113140 666540
rect 113380 666300 113490 666540
rect 113730 666300 113820 666540
rect 114060 666300 114150 666540
rect 114390 666300 114480 666540
rect 114720 666300 114830 666540
rect 115070 666300 115160 666540
rect 115400 666300 115490 666540
rect 115730 666300 115820 666540
rect 116060 666300 116170 666540
rect 116410 666300 116500 666540
rect 116740 666300 116830 666540
rect 117070 666300 117160 666540
rect 117400 666300 117510 666540
rect 117750 666300 117840 666540
rect 118080 666300 118170 666540
rect 118410 666300 118500 666540
rect 118740 666300 118850 666540
rect 119090 666300 119180 666540
rect 119420 666300 119510 666540
rect 119750 666300 119840 666540
rect 120080 666300 120190 666540
rect 120430 666300 120520 666540
rect 120760 666300 120850 666540
rect 121090 666300 121180 666540
rect 121420 666300 121530 666540
rect 121770 666300 121790 666540
rect 110790 666190 121790 666300
rect 110790 665950 110810 666190
rect 111050 665950 111140 666190
rect 111380 665950 111470 666190
rect 111710 665950 111800 666190
rect 112040 665950 112150 666190
rect 112390 665950 112480 666190
rect 112720 665950 112810 666190
rect 113050 665950 113140 666190
rect 113380 665950 113490 666190
rect 113730 665950 113820 666190
rect 114060 665950 114150 666190
rect 114390 665950 114480 666190
rect 114720 665950 114830 666190
rect 115070 665950 115160 666190
rect 115400 665950 115490 666190
rect 115730 665950 115820 666190
rect 116060 665950 116170 666190
rect 116410 665950 116500 666190
rect 116740 665950 116830 666190
rect 117070 665950 117160 666190
rect 117400 665950 117510 666190
rect 117750 665950 117840 666190
rect 118080 665950 118170 666190
rect 118410 665950 118500 666190
rect 118740 665950 118850 666190
rect 119090 665950 119180 666190
rect 119420 665950 119510 666190
rect 119750 665950 119840 666190
rect 120080 665950 120190 666190
rect 120430 665950 120520 666190
rect 120760 665950 120850 666190
rect 121090 665950 121180 666190
rect 121420 665950 121530 666190
rect 121770 665950 121790 666190
rect 110790 665860 121790 665950
rect 110790 665620 110810 665860
rect 111050 665620 111140 665860
rect 111380 665620 111470 665860
rect 111710 665620 111800 665860
rect 112040 665620 112150 665860
rect 112390 665620 112480 665860
rect 112720 665620 112810 665860
rect 113050 665620 113140 665860
rect 113380 665620 113490 665860
rect 113730 665620 113820 665860
rect 114060 665620 114150 665860
rect 114390 665620 114480 665860
rect 114720 665620 114830 665860
rect 115070 665620 115160 665860
rect 115400 665620 115490 665860
rect 115730 665620 115820 665860
rect 116060 665620 116170 665860
rect 116410 665620 116500 665860
rect 116740 665620 116830 665860
rect 117070 665620 117160 665860
rect 117400 665620 117510 665860
rect 117750 665620 117840 665860
rect 118080 665620 118170 665860
rect 118410 665620 118500 665860
rect 118740 665620 118850 665860
rect 119090 665620 119180 665860
rect 119420 665620 119510 665860
rect 119750 665620 119840 665860
rect 120080 665620 120190 665860
rect 120430 665620 120520 665860
rect 120760 665620 120850 665860
rect 121090 665620 121180 665860
rect 121420 665620 121530 665860
rect 121770 665620 121790 665860
rect 110790 665530 121790 665620
rect 110790 665290 110810 665530
rect 111050 665290 111140 665530
rect 111380 665290 111470 665530
rect 111710 665290 111800 665530
rect 112040 665290 112150 665530
rect 112390 665290 112480 665530
rect 112720 665290 112810 665530
rect 113050 665290 113140 665530
rect 113380 665290 113490 665530
rect 113730 665290 113820 665530
rect 114060 665290 114150 665530
rect 114390 665290 114480 665530
rect 114720 665290 114830 665530
rect 115070 665290 115160 665530
rect 115400 665290 115490 665530
rect 115730 665290 115820 665530
rect 116060 665290 116170 665530
rect 116410 665290 116500 665530
rect 116740 665290 116830 665530
rect 117070 665290 117160 665530
rect 117400 665290 117510 665530
rect 117750 665290 117840 665530
rect 118080 665290 118170 665530
rect 118410 665290 118500 665530
rect 118740 665290 118850 665530
rect 119090 665290 119180 665530
rect 119420 665290 119510 665530
rect 119750 665290 119840 665530
rect 120080 665290 120190 665530
rect 120430 665290 120520 665530
rect 120760 665290 120850 665530
rect 121090 665290 121180 665530
rect 121420 665290 121530 665530
rect 121770 665290 121790 665530
rect 110790 665200 121790 665290
rect 110790 664960 110810 665200
rect 111050 664960 111140 665200
rect 111380 664960 111470 665200
rect 111710 664960 111800 665200
rect 112040 664960 112150 665200
rect 112390 664960 112480 665200
rect 112720 664960 112810 665200
rect 113050 664960 113140 665200
rect 113380 664960 113490 665200
rect 113730 664960 113820 665200
rect 114060 664960 114150 665200
rect 114390 664960 114480 665200
rect 114720 664960 114830 665200
rect 115070 664960 115160 665200
rect 115400 664960 115490 665200
rect 115730 664960 115820 665200
rect 116060 664960 116170 665200
rect 116410 664960 116500 665200
rect 116740 664960 116830 665200
rect 117070 664960 117160 665200
rect 117400 664960 117510 665200
rect 117750 664960 117840 665200
rect 118080 664960 118170 665200
rect 118410 664960 118500 665200
rect 118740 664960 118850 665200
rect 119090 664960 119180 665200
rect 119420 664960 119510 665200
rect 119750 664960 119840 665200
rect 120080 664960 120190 665200
rect 120430 664960 120520 665200
rect 120760 664960 120850 665200
rect 121090 664960 121180 665200
rect 121420 664960 121530 665200
rect 121770 664960 121790 665200
rect 110790 664850 121790 664960
rect 110790 664610 110810 664850
rect 111050 664610 111140 664850
rect 111380 664610 111470 664850
rect 111710 664610 111800 664850
rect 112040 664610 112150 664850
rect 112390 664610 112480 664850
rect 112720 664610 112810 664850
rect 113050 664610 113140 664850
rect 113380 664610 113490 664850
rect 113730 664610 113820 664850
rect 114060 664610 114150 664850
rect 114390 664610 114480 664850
rect 114720 664610 114830 664850
rect 115070 664610 115160 664850
rect 115400 664610 115490 664850
rect 115730 664610 115820 664850
rect 116060 664610 116170 664850
rect 116410 664610 116500 664850
rect 116740 664610 116830 664850
rect 117070 664610 117160 664850
rect 117400 664610 117510 664850
rect 117750 664610 117840 664850
rect 118080 664610 118170 664850
rect 118410 664610 118500 664850
rect 118740 664610 118850 664850
rect 119090 664610 119180 664850
rect 119420 664610 119510 664850
rect 119750 664610 119840 664850
rect 120080 664610 120190 664850
rect 120430 664610 120520 664850
rect 120760 664610 120850 664850
rect 121090 664610 121180 664850
rect 121420 664610 121530 664850
rect 121770 664610 121790 664850
rect 110790 664520 121790 664610
rect 110790 664280 110810 664520
rect 111050 664280 111140 664520
rect 111380 664280 111470 664520
rect 111710 664280 111800 664520
rect 112040 664280 112150 664520
rect 112390 664280 112480 664520
rect 112720 664280 112810 664520
rect 113050 664280 113140 664520
rect 113380 664280 113490 664520
rect 113730 664280 113820 664520
rect 114060 664280 114150 664520
rect 114390 664280 114480 664520
rect 114720 664280 114830 664520
rect 115070 664280 115160 664520
rect 115400 664280 115490 664520
rect 115730 664280 115820 664520
rect 116060 664280 116170 664520
rect 116410 664280 116500 664520
rect 116740 664280 116830 664520
rect 117070 664280 117160 664520
rect 117400 664280 117510 664520
rect 117750 664280 117840 664520
rect 118080 664280 118170 664520
rect 118410 664280 118500 664520
rect 118740 664280 118850 664520
rect 119090 664280 119180 664520
rect 119420 664280 119510 664520
rect 119750 664280 119840 664520
rect 120080 664280 120190 664520
rect 120430 664280 120520 664520
rect 120760 664280 120850 664520
rect 121090 664280 121180 664520
rect 121420 664280 121530 664520
rect 121770 664280 121790 664520
rect 110790 664190 121790 664280
rect 110790 663950 110810 664190
rect 111050 663950 111140 664190
rect 111380 663950 111470 664190
rect 111710 663950 111800 664190
rect 112040 663950 112150 664190
rect 112390 663950 112480 664190
rect 112720 663950 112810 664190
rect 113050 663950 113140 664190
rect 113380 663950 113490 664190
rect 113730 663950 113820 664190
rect 114060 663950 114150 664190
rect 114390 663950 114480 664190
rect 114720 663950 114830 664190
rect 115070 663950 115160 664190
rect 115400 663950 115490 664190
rect 115730 663950 115820 664190
rect 116060 663950 116170 664190
rect 116410 663950 116500 664190
rect 116740 663950 116830 664190
rect 117070 663950 117160 664190
rect 117400 663950 117510 664190
rect 117750 663950 117840 664190
rect 118080 663950 118170 664190
rect 118410 663950 118500 664190
rect 118740 663950 118850 664190
rect 119090 663950 119180 664190
rect 119420 663950 119510 664190
rect 119750 663950 119840 664190
rect 120080 663950 120190 664190
rect 120430 663950 120520 664190
rect 120760 663950 120850 664190
rect 121090 663950 121180 664190
rect 121420 663950 121530 664190
rect 121770 663950 121790 664190
rect 110790 663860 121790 663950
rect 110790 663620 110810 663860
rect 111050 663620 111140 663860
rect 111380 663620 111470 663860
rect 111710 663620 111800 663860
rect 112040 663620 112150 663860
rect 112390 663620 112480 663860
rect 112720 663620 112810 663860
rect 113050 663620 113140 663860
rect 113380 663620 113490 663860
rect 113730 663620 113820 663860
rect 114060 663620 114150 663860
rect 114390 663620 114480 663860
rect 114720 663620 114830 663860
rect 115070 663620 115160 663860
rect 115400 663620 115490 663860
rect 115730 663620 115820 663860
rect 116060 663620 116170 663860
rect 116410 663620 116500 663860
rect 116740 663620 116830 663860
rect 117070 663620 117160 663860
rect 117400 663620 117510 663860
rect 117750 663620 117840 663860
rect 118080 663620 118170 663860
rect 118410 663620 118500 663860
rect 118740 663620 118850 663860
rect 119090 663620 119180 663860
rect 119420 663620 119510 663860
rect 119750 663620 119840 663860
rect 120080 663620 120190 663860
rect 120430 663620 120520 663860
rect 120760 663620 120850 663860
rect 121090 663620 121180 663860
rect 121420 663620 121530 663860
rect 121770 663620 121790 663860
rect 110790 663510 121790 663620
rect 110790 663270 110810 663510
rect 111050 663270 111140 663510
rect 111380 663270 111470 663510
rect 111710 663270 111800 663510
rect 112040 663270 112150 663510
rect 112390 663270 112480 663510
rect 112720 663270 112810 663510
rect 113050 663270 113140 663510
rect 113380 663270 113490 663510
rect 113730 663270 113820 663510
rect 114060 663270 114150 663510
rect 114390 663270 114480 663510
rect 114720 663270 114830 663510
rect 115070 663270 115160 663510
rect 115400 663270 115490 663510
rect 115730 663270 115820 663510
rect 116060 663270 116170 663510
rect 116410 663270 116500 663510
rect 116740 663270 116830 663510
rect 117070 663270 117160 663510
rect 117400 663270 117510 663510
rect 117750 663270 117840 663510
rect 118080 663270 118170 663510
rect 118410 663270 118500 663510
rect 118740 663270 118850 663510
rect 119090 663270 119180 663510
rect 119420 663270 119510 663510
rect 119750 663270 119840 663510
rect 120080 663270 120190 663510
rect 120430 663270 120520 663510
rect 120760 663270 120850 663510
rect 121090 663270 121180 663510
rect 121420 663270 121530 663510
rect 121770 663270 121790 663510
rect 110790 663180 121790 663270
rect 110790 662940 110810 663180
rect 111050 662940 111140 663180
rect 111380 662940 111470 663180
rect 111710 662940 111800 663180
rect 112040 662940 112150 663180
rect 112390 662940 112480 663180
rect 112720 662940 112810 663180
rect 113050 662940 113140 663180
rect 113380 662940 113490 663180
rect 113730 662940 113820 663180
rect 114060 662940 114150 663180
rect 114390 662940 114480 663180
rect 114720 662940 114830 663180
rect 115070 662940 115160 663180
rect 115400 662940 115490 663180
rect 115730 662940 115820 663180
rect 116060 662940 116170 663180
rect 116410 662940 116500 663180
rect 116740 662940 116830 663180
rect 117070 662940 117160 663180
rect 117400 662940 117510 663180
rect 117750 662940 117840 663180
rect 118080 662940 118170 663180
rect 118410 662940 118500 663180
rect 118740 662940 118850 663180
rect 119090 662940 119180 663180
rect 119420 662940 119510 663180
rect 119750 662940 119840 663180
rect 120080 662940 120190 663180
rect 120430 662940 120520 663180
rect 120760 662940 120850 663180
rect 121090 662940 121180 663180
rect 121420 662940 121530 663180
rect 121770 662940 121790 663180
rect 110790 662850 121790 662940
rect 110790 662610 110810 662850
rect 111050 662610 111140 662850
rect 111380 662610 111470 662850
rect 111710 662610 111800 662850
rect 112040 662610 112150 662850
rect 112390 662610 112480 662850
rect 112720 662610 112810 662850
rect 113050 662610 113140 662850
rect 113380 662610 113490 662850
rect 113730 662610 113820 662850
rect 114060 662610 114150 662850
rect 114390 662610 114480 662850
rect 114720 662610 114830 662850
rect 115070 662610 115160 662850
rect 115400 662610 115490 662850
rect 115730 662610 115820 662850
rect 116060 662610 116170 662850
rect 116410 662610 116500 662850
rect 116740 662610 116830 662850
rect 117070 662610 117160 662850
rect 117400 662610 117510 662850
rect 117750 662610 117840 662850
rect 118080 662610 118170 662850
rect 118410 662610 118500 662850
rect 118740 662610 118850 662850
rect 119090 662610 119180 662850
rect 119420 662610 119510 662850
rect 119750 662610 119840 662850
rect 120080 662610 120190 662850
rect 120430 662610 120520 662850
rect 120760 662610 120850 662850
rect 121090 662610 121180 662850
rect 121420 662610 121530 662850
rect 121770 662610 121790 662850
rect 110790 662520 121790 662610
rect 110790 662280 110810 662520
rect 111050 662280 111140 662520
rect 111380 662280 111470 662520
rect 111710 662280 111800 662520
rect 112040 662280 112150 662520
rect 112390 662280 112480 662520
rect 112720 662280 112810 662520
rect 113050 662280 113140 662520
rect 113380 662280 113490 662520
rect 113730 662280 113820 662520
rect 114060 662280 114150 662520
rect 114390 662280 114480 662520
rect 114720 662280 114830 662520
rect 115070 662280 115160 662520
rect 115400 662280 115490 662520
rect 115730 662280 115820 662520
rect 116060 662280 116170 662520
rect 116410 662280 116500 662520
rect 116740 662280 116830 662520
rect 117070 662280 117160 662520
rect 117400 662280 117510 662520
rect 117750 662280 117840 662520
rect 118080 662280 118170 662520
rect 118410 662280 118500 662520
rect 118740 662280 118850 662520
rect 119090 662280 119180 662520
rect 119420 662280 119510 662520
rect 119750 662280 119840 662520
rect 120080 662280 120190 662520
rect 120430 662280 120520 662520
rect 120760 662280 120850 662520
rect 121090 662280 121180 662520
rect 121420 662280 121530 662520
rect 121770 662280 121790 662520
rect 110790 662170 121790 662280
rect 110790 661930 110810 662170
rect 111050 661930 111140 662170
rect 111380 661930 111470 662170
rect 111710 661930 111800 662170
rect 112040 661930 112150 662170
rect 112390 661930 112480 662170
rect 112720 661930 112810 662170
rect 113050 661930 113140 662170
rect 113380 661930 113490 662170
rect 113730 661930 113820 662170
rect 114060 661930 114150 662170
rect 114390 661930 114480 662170
rect 114720 661930 114830 662170
rect 115070 661930 115160 662170
rect 115400 661930 115490 662170
rect 115730 661930 115820 662170
rect 116060 661930 116170 662170
rect 116410 661930 116500 662170
rect 116740 661930 116830 662170
rect 117070 661930 117160 662170
rect 117400 661930 117510 662170
rect 117750 661930 117840 662170
rect 118080 661930 118170 662170
rect 118410 661930 118500 662170
rect 118740 661930 118850 662170
rect 119090 661930 119180 662170
rect 119420 661930 119510 662170
rect 119750 661930 119840 662170
rect 120080 661930 120190 662170
rect 120430 661930 120520 662170
rect 120760 661930 120850 662170
rect 121090 661930 121180 662170
rect 121420 661930 121530 662170
rect 121770 661930 121790 662170
rect 110790 661840 121790 661930
rect 110790 661600 110810 661840
rect 111050 661600 111140 661840
rect 111380 661600 111470 661840
rect 111710 661600 111800 661840
rect 112040 661600 112150 661840
rect 112390 661600 112480 661840
rect 112720 661600 112810 661840
rect 113050 661600 113140 661840
rect 113380 661600 113490 661840
rect 113730 661600 113820 661840
rect 114060 661600 114150 661840
rect 114390 661600 114480 661840
rect 114720 661600 114830 661840
rect 115070 661600 115160 661840
rect 115400 661600 115490 661840
rect 115730 661600 115820 661840
rect 116060 661600 116170 661840
rect 116410 661600 116500 661840
rect 116740 661600 116830 661840
rect 117070 661600 117160 661840
rect 117400 661600 117510 661840
rect 117750 661600 117840 661840
rect 118080 661600 118170 661840
rect 118410 661600 118500 661840
rect 118740 661600 118850 661840
rect 119090 661600 119180 661840
rect 119420 661600 119510 661840
rect 119750 661600 119840 661840
rect 120080 661600 120190 661840
rect 120430 661600 120520 661840
rect 120760 661600 120850 661840
rect 121090 661600 121180 661840
rect 121420 661600 121530 661840
rect 121770 661600 121790 661840
rect 110790 661510 121790 661600
rect 110790 661270 110810 661510
rect 111050 661270 111140 661510
rect 111380 661270 111470 661510
rect 111710 661270 111800 661510
rect 112040 661270 112150 661510
rect 112390 661270 112480 661510
rect 112720 661270 112810 661510
rect 113050 661270 113140 661510
rect 113380 661270 113490 661510
rect 113730 661270 113820 661510
rect 114060 661270 114150 661510
rect 114390 661270 114480 661510
rect 114720 661270 114830 661510
rect 115070 661270 115160 661510
rect 115400 661270 115490 661510
rect 115730 661270 115820 661510
rect 116060 661270 116170 661510
rect 116410 661270 116500 661510
rect 116740 661270 116830 661510
rect 117070 661270 117160 661510
rect 117400 661270 117510 661510
rect 117750 661270 117840 661510
rect 118080 661270 118170 661510
rect 118410 661270 118500 661510
rect 118740 661270 118850 661510
rect 119090 661270 119180 661510
rect 119420 661270 119510 661510
rect 119750 661270 119840 661510
rect 120080 661270 120190 661510
rect 120430 661270 120520 661510
rect 120760 661270 120850 661510
rect 121090 661270 121180 661510
rect 121420 661270 121530 661510
rect 121770 661270 121790 661510
rect 110790 661180 121790 661270
rect 110790 660940 110810 661180
rect 111050 660940 111140 661180
rect 111380 660940 111470 661180
rect 111710 660940 111800 661180
rect 112040 660940 112150 661180
rect 112390 660940 112480 661180
rect 112720 660940 112810 661180
rect 113050 660940 113140 661180
rect 113380 660940 113490 661180
rect 113730 660940 113820 661180
rect 114060 660940 114150 661180
rect 114390 660940 114480 661180
rect 114720 660940 114830 661180
rect 115070 660940 115160 661180
rect 115400 660940 115490 661180
rect 115730 660940 115820 661180
rect 116060 660940 116170 661180
rect 116410 660940 116500 661180
rect 116740 660940 116830 661180
rect 117070 660940 117160 661180
rect 117400 660940 117510 661180
rect 117750 660940 117840 661180
rect 118080 660940 118170 661180
rect 118410 660940 118500 661180
rect 118740 660940 118850 661180
rect 119090 660940 119180 661180
rect 119420 660940 119510 661180
rect 119750 660940 119840 661180
rect 120080 660940 120190 661180
rect 120430 660940 120520 661180
rect 120760 660940 120850 661180
rect 121090 660940 121180 661180
rect 121420 660940 121530 661180
rect 121770 660940 121790 661180
rect 110790 660920 121790 660940
rect 122170 671900 133170 671920
rect 122170 671660 122190 671900
rect 122430 671660 122520 671900
rect 122760 671660 122850 671900
rect 123090 671660 123180 671900
rect 123420 671660 123530 671900
rect 123770 671660 123860 671900
rect 124100 671660 124190 671900
rect 124430 671660 124520 671900
rect 124760 671660 124870 671900
rect 125110 671660 125200 671900
rect 125440 671660 125530 671900
rect 125770 671660 125860 671900
rect 126100 671660 126210 671900
rect 126450 671660 126540 671900
rect 126780 671660 126870 671900
rect 127110 671660 127200 671900
rect 127440 671660 127550 671900
rect 127790 671660 127880 671900
rect 128120 671660 128210 671900
rect 128450 671660 128540 671900
rect 128780 671660 128890 671900
rect 129130 671660 129220 671900
rect 129460 671660 129550 671900
rect 129790 671660 129880 671900
rect 130120 671660 130230 671900
rect 130470 671660 130560 671900
rect 130800 671660 130890 671900
rect 131130 671660 131220 671900
rect 131460 671660 131570 671900
rect 131810 671660 131900 671900
rect 132140 671660 132230 671900
rect 132470 671660 132560 671900
rect 132800 671660 132910 671900
rect 133150 671660 133170 671900
rect 122170 671550 133170 671660
rect 122170 671310 122190 671550
rect 122430 671310 122520 671550
rect 122760 671310 122850 671550
rect 123090 671310 123180 671550
rect 123420 671310 123530 671550
rect 123770 671310 123860 671550
rect 124100 671310 124190 671550
rect 124430 671310 124520 671550
rect 124760 671310 124870 671550
rect 125110 671310 125200 671550
rect 125440 671310 125530 671550
rect 125770 671310 125860 671550
rect 126100 671310 126210 671550
rect 126450 671310 126540 671550
rect 126780 671310 126870 671550
rect 127110 671310 127200 671550
rect 127440 671310 127550 671550
rect 127790 671310 127880 671550
rect 128120 671310 128210 671550
rect 128450 671310 128540 671550
rect 128780 671310 128890 671550
rect 129130 671310 129220 671550
rect 129460 671310 129550 671550
rect 129790 671310 129880 671550
rect 130120 671310 130230 671550
rect 130470 671310 130560 671550
rect 130800 671310 130890 671550
rect 131130 671310 131220 671550
rect 131460 671310 131570 671550
rect 131810 671310 131900 671550
rect 132140 671310 132230 671550
rect 132470 671310 132560 671550
rect 132800 671310 132910 671550
rect 133150 671310 133170 671550
rect 122170 671220 133170 671310
rect 122170 670980 122190 671220
rect 122430 670980 122520 671220
rect 122760 670980 122850 671220
rect 123090 670980 123180 671220
rect 123420 670980 123530 671220
rect 123770 670980 123860 671220
rect 124100 670980 124190 671220
rect 124430 670980 124520 671220
rect 124760 670980 124870 671220
rect 125110 670980 125200 671220
rect 125440 670980 125530 671220
rect 125770 670980 125860 671220
rect 126100 670980 126210 671220
rect 126450 670980 126540 671220
rect 126780 670980 126870 671220
rect 127110 670980 127200 671220
rect 127440 670980 127550 671220
rect 127790 670980 127880 671220
rect 128120 670980 128210 671220
rect 128450 670980 128540 671220
rect 128780 670980 128890 671220
rect 129130 670980 129220 671220
rect 129460 670980 129550 671220
rect 129790 670980 129880 671220
rect 130120 670980 130230 671220
rect 130470 670980 130560 671220
rect 130800 670980 130890 671220
rect 131130 670980 131220 671220
rect 131460 670980 131570 671220
rect 131810 670980 131900 671220
rect 132140 670980 132230 671220
rect 132470 670980 132560 671220
rect 132800 670980 132910 671220
rect 133150 670980 133170 671220
rect 122170 670890 133170 670980
rect 122170 670650 122190 670890
rect 122430 670650 122520 670890
rect 122760 670650 122850 670890
rect 123090 670650 123180 670890
rect 123420 670650 123530 670890
rect 123770 670650 123860 670890
rect 124100 670650 124190 670890
rect 124430 670650 124520 670890
rect 124760 670650 124870 670890
rect 125110 670650 125200 670890
rect 125440 670650 125530 670890
rect 125770 670650 125860 670890
rect 126100 670650 126210 670890
rect 126450 670650 126540 670890
rect 126780 670650 126870 670890
rect 127110 670650 127200 670890
rect 127440 670650 127550 670890
rect 127790 670650 127880 670890
rect 128120 670650 128210 670890
rect 128450 670650 128540 670890
rect 128780 670650 128890 670890
rect 129130 670650 129220 670890
rect 129460 670650 129550 670890
rect 129790 670650 129880 670890
rect 130120 670650 130230 670890
rect 130470 670650 130560 670890
rect 130800 670650 130890 670890
rect 131130 670650 131220 670890
rect 131460 670650 131570 670890
rect 131810 670650 131900 670890
rect 132140 670650 132230 670890
rect 132470 670650 132560 670890
rect 132800 670650 132910 670890
rect 133150 670650 133170 670890
rect 122170 670560 133170 670650
rect 122170 670320 122190 670560
rect 122430 670320 122520 670560
rect 122760 670320 122850 670560
rect 123090 670320 123180 670560
rect 123420 670320 123530 670560
rect 123770 670320 123860 670560
rect 124100 670320 124190 670560
rect 124430 670320 124520 670560
rect 124760 670320 124870 670560
rect 125110 670320 125200 670560
rect 125440 670320 125530 670560
rect 125770 670320 125860 670560
rect 126100 670320 126210 670560
rect 126450 670320 126540 670560
rect 126780 670320 126870 670560
rect 127110 670320 127200 670560
rect 127440 670320 127550 670560
rect 127790 670320 127880 670560
rect 128120 670320 128210 670560
rect 128450 670320 128540 670560
rect 128780 670320 128890 670560
rect 129130 670320 129220 670560
rect 129460 670320 129550 670560
rect 129790 670320 129880 670560
rect 130120 670320 130230 670560
rect 130470 670320 130560 670560
rect 130800 670320 130890 670560
rect 131130 670320 131220 670560
rect 131460 670320 131570 670560
rect 131810 670320 131900 670560
rect 132140 670320 132230 670560
rect 132470 670320 132560 670560
rect 132800 670320 132910 670560
rect 133150 670320 133170 670560
rect 122170 670210 133170 670320
rect 122170 669970 122190 670210
rect 122430 669970 122520 670210
rect 122760 669970 122850 670210
rect 123090 669970 123180 670210
rect 123420 669970 123530 670210
rect 123770 669970 123860 670210
rect 124100 669970 124190 670210
rect 124430 669970 124520 670210
rect 124760 669970 124870 670210
rect 125110 669970 125200 670210
rect 125440 669970 125530 670210
rect 125770 669970 125860 670210
rect 126100 669970 126210 670210
rect 126450 669970 126540 670210
rect 126780 669970 126870 670210
rect 127110 669970 127200 670210
rect 127440 669970 127550 670210
rect 127790 669970 127880 670210
rect 128120 669970 128210 670210
rect 128450 669970 128540 670210
rect 128780 669970 128890 670210
rect 129130 669970 129220 670210
rect 129460 669970 129550 670210
rect 129790 669970 129880 670210
rect 130120 669970 130230 670210
rect 130470 669970 130560 670210
rect 130800 669970 130890 670210
rect 131130 669970 131220 670210
rect 131460 669970 131570 670210
rect 131810 669970 131900 670210
rect 132140 669970 132230 670210
rect 132470 669970 132560 670210
rect 132800 669970 132910 670210
rect 133150 669970 133170 670210
rect 122170 669880 133170 669970
rect 122170 669640 122190 669880
rect 122430 669640 122520 669880
rect 122760 669640 122850 669880
rect 123090 669640 123180 669880
rect 123420 669640 123530 669880
rect 123770 669640 123860 669880
rect 124100 669640 124190 669880
rect 124430 669640 124520 669880
rect 124760 669640 124870 669880
rect 125110 669640 125200 669880
rect 125440 669640 125530 669880
rect 125770 669640 125860 669880
rect 126100 669640 126210 669880
rect 126450 669640 126540 669880
rect 126780 669640 126870 669880
rect 127110 669640 127200 669880
rect 127440 669640 127550 669880
rect 127790 669640 127880 669880
rect 128120 669640 128210 669880
rect 128450 669640 128540 669880
rect 128780 669640 128890 669880
rect 129130 669640 129220 669880
rect 129460 669640 129550 669880
rect 129790 669640 129880 669880
rect 130120 669640 130230 669880
rect 130470 669640 130560 669880
rect 130800 669640 130890 669880
rect 131130 669640 131220 669880
rect 131460 669640 131570 669880
rect 131810 669640 131900 669880
rect 132140 669640 132230 669880
rect 132470 669640 132560 669880
rect 132800 669640 132910 669880
rect 133150 669640 133170 669880
rect 122170 669550 133170 669640
rect 122170 669310 122190 669550
rect 122430 669310 122520 669550
rect 122760 669310 122850 669550
rect 123090 669310 123180 669550
rect 123420 669310 123530 669550
rect 123770 669310 123860 669550
rect 124100 669310 124190 669550
rect 124430 669310 124520 669550
rect 124760 669310 124870 669550
rect 125110 669310 125200 669550
rect 125440 669310 125530 669550
rect 125770 669310 125860 669550
rect 126100 669310 126210 669550
rect 126450 669310 126540 669550
rect 126780 669310 126870 669550
rect 127110 669310 127200 669550
rect 127440 669310 127550 669550
rect 127790 669310 127880 669550
rect 128120 669310 128210 669550
rect 128450 669310 128540 669550
rect 128780 669310 128890 669550
rect 129130 669310 129220 669550
rect 129460 669310 129550 669550
rect 129790 669310 129880 669550
rect 130120 669310 130230 669550
rect 130470 669310 130560 669550
rect 130800 669310 130890 669550
rect 131130 669310 131220 669550
rect 131460 669310 131570 669550
rect 131810 669310 131900 669550
rect 132140 669310 132230 669550
rect 132470 669310 132560 669550
rect 132800 669310 132910 669550
rect 133150 669310 133170 669550
rect 122170 669220 133170 669310
rect 122170 668980 122190 669220
rect 122430 668980 122520 669220
rect 122760 668980 122850 669220
rect 123090 668980 123180 669220
rect 123420 668980 123530 669220
rect 123770 668980 123860 669220
rect 124100 668980 124190 669220
rect 124430 668980 124520 669220
rect 124760 668980 124870 669220
rect 125110 668980 125200 669220
rect 125440 668980 125530 669220
rect 125770 668980 125860 669220
rect 126100 668980 126210 669220
rect 126450 668980 126540 669220
rect 126780 668980 126870 669220
rect 127110 668980 127200 669220
rect 127440 668980 127550 669220
rect 127790 668980 127880 669220
rect 128120 668980 128210 669220
rect 128450 668980 128540 669220
rect 128780 668980 128890 669220
rect 129130 668980 129220 669220
rect 129460 668980 129550 669220
rect 129790 668980 129880 669220
rect 130120 668980 130230 669220
rect 130470 668980 130560 669220
rect 130800 668980 130890 669220
rect 131130 668980 131220 669220
rect 131460 668980 131570 669220
rect 131810 668980 131900 669220
rect 132140 668980 132230 669220
rect 132470 668980 132560 669220
rect 132800 668980 132910 669220
rect 133150 668980 133170 669220
rect 122170 668870 133170 668980
rect 122170 668630 122190 668870
rect 122430 668630 122520 668870
rect 122760 668630 122850 668870
rect 123090 668630 123180 668870
rect 123420 668630 123530 668870
rect 123770 668630 123860 668870
rect 124100 668630 124190 668870
rect 124430 668630 124520 668870
rect 124760 668630 124870 668870
rect 125110 668630 125200 668870
rect 125440 668630 125530 668870
rect 125770 668630 125860 668870
rect 126100 668630 126210 668870
rect 126450 668630 126540 668870
rect 126780 668630 126870 668870
rect 127110 668630 127200 668870
rect 127440 668630 127550 668870
rect 127790 668630 127880 668870
rect 128120 668630 128210 668870
rect 128450 668630 128540 668870
rect 128780 668630 128890 668870
rect 129130 668630 129220 668870
rect 129460 668630 129550 668870
rect 129790 668630 129880 668870
rect 130120 668630 130230 668870
rect 130470 668630 130560 668870
rect 130800 668630 130890 668870
rect 131130 668630 131220 668870
rect 131460 668630 131570 668870
rect 131810 668630 131900 668870
rect 132140 668630 132230 668870
rect 132470 668630 132560 668870
rect 132800 668630 132910 668870
rect 133150 668630 133170 668870
rect 122170 668540 133170 668630
rect 122170 668300 122190 668540
rect 122430 668300 122520 668540
rect 122760 668300 122850 668540
rect 123090 668300 123180 668540
rect 123420 668300 123530 668540
rect 123770 668300 123860 668540
rect 124100 668300 124190 668540
rect 124430 668300 124520 668540
rect 124760 668300 124870 668540
rect 125110 668300 125200 668540
rect 125440 668300 125530 668540
rect 125770 668300 125860 668540
rect 126100 668300 126210 668540
rect 126450 668300 126540 668540
rect 126780 668300 126870 668540
rect 127110 668300 127200 668540
rect 127440 668300 127550 668540
rect 127790 668300 127880 668540
rect 128120 668300 128210 668540
rect 128450 668300 128540 668540
rect 128780 668300 128890 668540
rect 129130 668300 129220 668540
rect 129460 668300 129550 668540
rect 129790 668300 129880 668540
rect 130120 668300 130230 668540
rect 130470 668300 130560 668540
rect 130800 668300 130890 668540
rect 131130 668300 131220 668540
rect 131460 668300 131570 668540
rect 131810 668300 131900 668540
rect 132140 668300 132230 668540
rect 132470 668300 132560 668540
rect 132800 668300 132910 668540
rect 133150 668300 133170 668540
rect 122170 668210 133170 668300
rect 122170 667970 122190 668210
rect 122430 667970 122520 668210
rect 122760 667970 122850 668210
rect 123090 667970 123180 668210
rect 123420 667970 123530 668210
rect 123770 667970 123860 668210
rect 124100 667970 124190 668210
rect 124430 667970 124520 668210
rect 124760 667970 124870 668210
rect 125110 667970 125200 668210
rect 125440 667970 125530 668210
rect 125770 667970 125860 668210
rect 126100 667970 126210 668210
rect 126450 667970 126540 668210
rect 126780 667970 126870 668210
rect 127110 667970 127200 668210
rect 127440 667970 127550 668210
rect 127790 667970 127880 668210
rect 128120 667970 128210 668210
rect 128450 667970 128540 668210
rect 128780 667970 128890 668210
rect 129130 667970 129220 668210
rect 129460 667970 129550 668210
rect 129790 667970 129880 668210
rect 130120 667970 130230 668210
rect 130470 667970 130560 668210
rect 130800 667970 130890 668210
rect 131130 667970 131220 668210
rect 131460 667970 131570 668210
rect 131810 667970 131900 668210
rect 132140 667970 132230 668210
rect 132470 667970 132560 668210
rect 132800 667970 132910 668210
rect 133150 667970 133170 668210
rect 122170 667880 133170 667970
rect 122170 667640 122190 667880
rect 122430 667640 122520 667880
rect 122760 667640 122850 667880
rect 123090 667640 123180 667880
rect 123420 667640 123530 667880
rect 123770 667640 123860 667880
rect 124100 667640 124190 667880
rect 124430 667640 124520 667880
rect 124760 667640 124870 667880
rect 125110 667640 125200 667880
rect 125440 667640 125530 667880
rect 125770 667640 125860 667880
rect 126100 667640 126210 667880
rect 126450 667640 126540 667880
rect 126780 667640 126870 667880
rect 127110 667640 127200 667880
rect 127440 667640 127550 667880
rect 127790 667640 127880 667880
rect 128120 667640 128210 667880
rect 128450 667640 128540 667880
rect 128780 667640 128890 667880
rect 129130 667640 129220 667880
rect 129460 667640 129550 667880
rect 129790 667640 129880 667880
rect 130120 667640 130230 667880
rect 130470 667640 130560 667880
rect 130800 667640 130890 667880
rect 131130 667640 131220 667880
rect 131460 667640 131570 667880
rect 131810 667640 131900 667880
rect 132140 667640 132230 667880
rect 132470 667640 132560 667880
rect 132800 667640 132910 667880
rect 133150 667640 133170 667880
rect 122170 667530 133170 667640
rect 122170 667290 122190 667530
rect 122430 667290 122520 667530
rect 122760 667290 122850 667530
rect 123090 667290 123180 667530
rect 123420 667290 123530 667530
rect 123770 667290 123860 667530
rect 124100 667290 124190 667530
rect 124430 667290 124520 667530
rect 124760 667290 124870 667530
rect 125110 667290 125200 667530
rect 125440 667290 125530 667530
rect 125770 667290 125860 667530
rect 126100 667290 126210 667530
rect 126450 667290 126540 667530
rect 126780 667290 126870 667530
rect 127110 667290 127200 667530
rect 127440 667290 127550 667530
rect 127790 667290 127880 667530
rect 128120 667290 128210 667530
rect 128450 667290 128540 667530
rect 128780 667290 128890 667530
rect 129130 667290 129220 667530
rect 129460 667290 129550 667530
rect 129790 667290 129880 667530
rect 130120 667290 130230 667530
rect 130470 667290 130560 667530
rect 130800 667290 130890 667530
rect 131130 667290 131220 667530
rect 131460 667290 131570 667530
rect 131810 667290 131900 667530
rect 132140 667290 132230 667530
rect 132470 667290 132560 667530
rect 132800 667290 132910 667530
rect 133150 667290 133170 667530
rect 122170 667200 133170 667290
rect 122170 666960 122190 667200
rect 122430 666960 122520 667200
rect 122760 666960 122850 667200
rect 123090 666960 123180 667200
rect 123420 666960 123530 667200
rect 123770 666960 123860 667200
rect 124100 666960 124190 667200
rect 124430 666960 124520 667200
rect 124760 666960 124870 667200
rect 125110 666960 125200 667200
rect 125440 666960 125530 667200
rect 125770 666960 125860 667200
rect 126100 666960 126210 667200
rect 126450 666960 126540 667200
rect 126780 666960 126870 667200
rect 127110 666960 127200 667200
rect 127440 666960 127550 667200
rect 127790 666960 127880 667200
rect 128120 666960 128210 667200
rect 128450 666960 128540 667200
rect 128780 666960 128890 667200
rect 129130 666960 129220 667200
rect 129460 666960 129550 667200
rect 129790 666960 129880 667200
rect 130120 666960 130230 667200
rect 130470 666960 130560 667200
rect 130800 666960 130890 667200
rect 131130 666960 131220 667200
rect 131460 666960 131570 667200
rect 131810 666960 131900 667200
rect 132140 666960 132230 667200
rect 132470 666960 132560 667200
rect 132800 666960 132910 667200
rect 133150 666960 133170 667200
rect 122170 666870 133170 666960
rect 122170 666630 122190 666870
rect 122430 666630 122520 666870
rect 122760 666630 122850 666870
rect 123090 666630 123180 666870
rect 123420 666630 123530 666870
rect 123770 666630 123860 666870
rect 124100 666630 124190 666870
rect 124430 666630 124520 666870
rect 124760 666630 124870 666870
rect 125110 666630 125200 666870
rect 125440 666630 125530 666870
rect 125770 666630 125860 666870
rect 126100 666630 126210 666870
rect 126450 666630 126540 666870
rect 126780 666630 126870 666870
rect 127110 666630 127200 666870
rect 127440 666630 127550 666870
rect 127790 666630 127880 666870
rect 128120 666630 128210 666870
rect 128450 666630 128540 666870
rect 128780 666630 128890 666870
rect 129130 666630 129220 666870
rect 129460 666630 129550 666870
rect 129790 666630 129880 666870
rect 130120 666630 130230 666870
rect 130470 666630 130560 666870
rect 130800 666630 130890 666870
rect 131130 666630 131220 666870
rect 131460 666630 131570 666870
rect 131810 666630 131900 666870
rect 132140 666630 132230 666870
rect 132470 666630 132560 666870
rect 132800 666630 132910 666870
rect 133150 666630 133170 666870
rect 122170 666540 133170 666630
rect 122170 666300 122190 666540
rect 122430 666300 122520 666540
rect 122760 666300 122850 666540
rect 123090 666300 123180 666540
rect 123420 666300 123530 666540
rect 123770 666300 123860 666540
rect 124100 666300 124190 666540
rect 124430 666300 124520 666540
rect 124760 666300 124870 666540
rect 125110 666300 125200 666540
rect 125440 666300 125530 666540
rect 125770 666300 125860 666540
rect 126100 666300 126210 666540
rect 126450 666300 126540 666540
rect 126780 666300 126870 666540
rect 127110 666300 127200 666540
rect 127440 666300 127550 666540
rect 127790 666300 127880 666540
rect 128120 666300 128210 666540
rect 128450 666300 128540 666540
rect 128780 666300 128890 666540
rect 129130 666300 129220 666540
rect 129460 666300 129550 666540
rect 129790 666300 129880 666540
rect 130120 666300 130230 666540
rect 130470 666300 130560 666540
rect 130800 666300 130890 666540
rect 131130 666300 131220 666540
rect 131460 666300 131570 666540
rect 131810 666300 131900 666540
rect 132140 666300 132230 666540
rect 132470 666300 132560 666540
rect 132800 666300 132910 666540
rect 133150 666300 133170 666540
rect 122170 666190 133170 666300
rect 122170 665950 122190 666190
rect 122430 665950 122520 666190
rect 122760 665950 122850 666190
rect 123090 665950 123180 666190
rect 123420 665950 123530 666190
rect 123770 665950 123860 666190
rect 124100 665950 124190 666190
rect 124430 665950 124520 666190
rect 124760 665950 124870 666190
rect 125110 665950 125200 666190
rect 125440 665950 125530 666190
rect 125770 665950 125860 666190
rect 126100 665950 126210 666190
rect 126450 665950 126540 666190
rect 126780 665950 126870 666190
rect 127110 665950 127200 666190
rect 127440 665950 127550 666190
rect 127790 665950 127880 666190
rect 128120 665950 128210 666190
rect 128450 665950 128540 666190
rect 128780 665950 128890 666190
rect 129130 665950 129220 666190
rect 129460 665950 129550 666190
rect 129790 665950 129880 666190
rect 130120 665950 130230 666190
rect 130470 665950 130560 666190
rect 130800 665950 130890 666190
rect 131130 665950 131220 666190
rect 131460 665950 131570 666190
rect 131810 665950 131900 666190
rect 132140 665950 132230 666190
rect 132470 665950 132560 666190
rect 132800 665950 132910 666190
rect 133150 665950 133170 666190
rect 122170 665860 133170 665950
rect 122170 665620 122190 665860
rect 122430 665620 122520 665860
rect 122760 665620 122850 665860
rect 123090 665620 123180 665860
rect 123420 665620 123530 665860
rect 123770 665620 123860 665860
rect 124100 665620 124190 665860
rect 124430 665620 124520 665860
rect 124760 665620 124870 665860
rect 125110 665620 125200 665860
rect 125440 665620 125530 665860
rect 125770 665620 125860 665860
rect 126100 665620 126210 665860
rect 126450 665620 126540 665860
rect 126780 665620 126870 665860
rect 127110 665620 127200 665860
rect 127440 665620 127550 665860
rect 127790 665620 127880 665860
rect 128120 665620 128210 665860
rect 128450 665620 128540 665860
rect 128780 665620 128890 665860
rect 129130 665620 129220 665860
rect 129460 665620 129550 665860
rect 129790 665620 129880 665860
rect 130120 665620 130230 665860
rect 130470 665620 130560 665860
rect 130800 665620 130890 665860
rect 131130 665620 131220 665860
rect 131460 665620 131570 665860
rect 131810 665620 131900 665860
rect 132140 665620 132230 665860
rect 132470 665620 132560 665860
rect 132800 665620 132910 665860
rect 133150 665620 133170 665860
rect 122170 665530 133170 665620
rect 122170 665290 122190 665530
rect 122430 665290 122520 665530
rect 122760 665290 122850 665530
rect 123090 665290 123180 665530
rect 123420 665290 123530 665530
rect 123770 665290 123860 665530
rect 124100 665290 124190 665530
rect 124430 665290 124520 665530
rect 124760 665290 124870 665530
rect 125110 665290 125200 665530
rect 125440 665290 125530 665530
rect 125770 665290 125860 665530
rect 126100 665290 126210 665530
rect 126450 665290 126540 665530
rect 126780 665290 126870 665530
rect 127110 665290 127200 665530
rect 127440 665290 127550 665530
rect 127790 665290 127880 665530
rect 128120 665290 128210 665530
rect 128450 665290 128540 665530
rect 128780 665290 128890 665530
rect 129130 665290 129220 665530
rect 129460 665290 129550 665530
rect 129790 665290 129880 665530
rect 130120 665290 130230 665530
rect 130470 665290 130560 665530
rect 130800 665290 130890 665530
rect 131130 665290 131220 665530
rect 131460 665290 131570 665530
rect 131810 665290 131900 665530
rect 132140 665290 132230 665530
rect 132470 665290 132560 665530
rect 132800 665290 132910 665530
rect 133150 665290 133170 665530
rect 122170 665200 133170 665290
rect 122170 664960 122190 665200
rect 122430 664960 122520 665200
rect 122760 664960 122850 665200
rect 123090 664960 123180 665200
rect 123420 664960 123530 665200
rect 123770 664960 123860 665200
rect 124100 664960 124190 665200
rect 124430 664960 124520 665200
rect 124760 664960 124870 665200
rect 125110 664960 125200 665200
rect 125440 664960 125530 665200
rect 125770 664960 125860 665200
rect 126100 664960 126210 665200
rect 126450 664960 126540 665200
rect 126780 664960 126870 665200
rect 127110 664960 127200 665200
rect 127440 664960 127550 665200
rect 127790 664960 127880 665200
rect 128120 664960 128210 665200
rect 128450 664960 128540 665200
rect 128780 664960 128890 665200
rect 129130 664960 129220 665200
rect 129460 664960 129550 665200
rect 129790 664960 129880 665200
rect 130120 664960 130230 665200
rect 130470 664960 130560 665200
rect 130800 664960 130890 665200
rect 131130 664960 131220 665200
rect 131460 664960 131570 665200
rect 131810 664960 131900 665200
rect 132140 664960 132230 665200
rect 132470 664960 132560 665200
rect 132800 664960 132910 665200
rect 133150 664960 133170 665200
rect 122170 664850 133170 664960
rect 122170 664610 122190 664850
rect 122430 664610 122520 664850
rect 122760 664610 122850 664850
rect 123090 664610 123180 664850
rect 123420 664610 123530 664850
rect 123770 664610 123860 664850
rect 124100 664610 124190 664850
rect 124430 664610 124520 664850
rect 124760 664610 124870 664850
rect 125110 664610 125200 664850
rect 125440 664610 125530 664850
rect 125770 664610 125860 664850
rect 126100 664610 126210 664850
rect 126450 664610 126540 664850
rect 126780 664610 126870 664850
rect 127110 664610 127200 664850
rect 127440 664610 127550 664850
rect 127790 664610 127880 664850
rect 128120 664610 128210 664850
rect 128450 664610 128540 664850
rect 128780 664610 128890 664850
rect 129130 664610 129220 664850
rect 129460 664610 129550 664850
rect 129790 664610 129880 664850
rect 130120 664610 130230 664850
rect 130470 664610 130560 664850
rect 130800 664610 130890 664850
rect 131130 664610 131220 664850
rect 131460 664610 131570 664850
rect 131810 664610 131900 664850
rect 132140 664610 132230 664850
rect 132470 664610 132560 664850
rect 132800 664610 132910 664850
rect 133150 664610 133170 664850
rect 122170 664520 133170 664610
rect 122170 664280 122190 664520
rect 122430 664280 122520 664520
rect 122760 664280 122850 664520
rect 123090 664280 123180 664520
rect 123420 664280 123530 664520
rect 123770 664280 123860 664520
rect 124100 664280 124190 664520
rect 124430 664280 124520 664520
rect 124760 664280 124870 664520
rect 125110 664280 125200 664520
rect 125440 664280 125530 664520
rect 125770 664280 125860 664520
rect 126100 664280 126210 664520
rect 126450 664280 126540 664520
rect 126780 664280 126870 664520
rect 127110 664280 127200 664520
rect 127440 664280 127550 664520
rect 127790 664280 127880 664520
rect 128120 664280 128210 664520
rect 128450 664280 128540 664520
rect 128780 664280 128890 664520
rect 129130 664280 129220 664520
rect 129460 664280 129550 664520
rect 129790 664280 129880 664520
rect 130120 664280 130230 664520
rect 130470 664280 130560 664520
rect 130800 664280 130890 664520
rect 131130 664280 131220 664520
rect 131460 664280 131570 664520
rect 131810 664280 131900 664520
rect 132140 664280 132230 664520
rect 132470 664280 132560 664520
rect 132800 664280 132910 664520
rect 133150 664280 133170 664520
rect 122170 664190 133170 664280
rect 122170 663950 122190 664190
rect 122430 663950 122520 664190
rect 122760 663950 122850 664190
rect 123090 663950 123180 664190
rect 123420 663950 123530 664190
rect 123770 663950 123860 664190
rect 124100 663950 124190 664190
rect 124430 663950 124520 664190
rect 124760 663950 124870 664190
rect 125110 663950 125200 664190
rect 125440 663950 125530 664190
rect 125770 663950 125860 664190
rect 126100 663950 126210 664190
rect 126450 663950 126540 664190
rect 126780 663950 126870 664190
rect 127110 663950 127200 664190
rect 127440 663950 127550 664190
rect 127790 663950 127880 664190
rect 128120 663950 128210 664190
rect 128450 663950 128540 664190
rect 128780 663950 128890 664190
rect 129130 663950 129220 664190
rect 129460 663950 129550 664190
rect 129790 663950 129880 664190
rect 130120 663950 130230 664190
rect 130470 663950 130560 664190
rect 130800 663950 130890 664190
rect 131130 663950 131220 664190
rect 131460 663950 131570 664190
rect 131810 663950 131900 664190
rect 132140 663950 132230 664190
rect 132470 663950 132560 664190
rect 132800 663950 132910 664190
rect 133150 663950 133170 664190
rect 122170 663860 133170 663950
rect 122170 663620 122190 663860
rect 122430 663620 122520 663860
rect 122760 663620 122850 663860
rect 123090 663620 123180 663860
rect 123420 663620 123530 663860
rect 123770 663620 123860 663860
rect 124100 663620 124190 663860
rect 124430 663620 124520 663860
rect 124760 663620 124870 663860
rect 125110 663620 125200 663860
rect 125440 663620 125530 663860
rect 125770 663620 125860 663860
rect 126100 663620 126210 663860
rect 126450 663620 126540 663860
rect 126780 663620 126870 663860
rect 127110 663620 127200 663860
rect 127440 663620 127550 663860
rect 127790 663620 127880 663860
rect 128120 663620 128210 663860
rect 128450 663620 128540 663860
rect 128780 663620 128890 663860
rect 129130 663620 129220 663860
rect 129460 663620 129550 663860
rect 129790 663620 129880 663860
rect 130120 663620 130230 663860
rect 130470 663620 130560 663860
rect 130800 663620 130890 663860
rect 131130 663620 131220 663860
rect 131460 663620 131570 663860
rect 131810 663620 131900 663860
rect 132140 663620 132230 663860
rect 132470 663620 132560 663860
rect 132800 663620 132910 663860
rect 133150 663620 133170 663860
rect 122170 663510 133170 663620
rect 122170 663270 122190 663510
rect 122430 663270 122520 663510
rect 122760 663270 122850 663510
rect 123090 663270 123180 663510
rect 123420 663270 123530 663510
rect 123770 663270 123860 663510
rect 124100 663270 124190 663510
rect 124430 663270 124520 663510
rect 124760 663270 124870 663510
rect 125110 663270 125200 663510
rect 125440 663270 125530 663510
rect 125770 663270 125860 663510
rect 126100 663270 126210 663510
rect 126450 663270 126540 663510
rect 126780 663270 126870 663510
rect 127110 663270 127200 663510
rect 127440 663270 127550 663510
rect 127790 663270 127880 663510
rect 128120 663270 128210 663510
rect 128450 663270 128540 663510
rect 128780 663270 128890 663510
rect 129130 663270 129220 663510
rect 129460 663270 129550 663510
rect 129790 663270 129880 663510
rect 130120 663270 130230 663510
rect 130470 663270 130560 663510
rect 130800 663270 130890 663510
rect 131130 663270 131220 663510
rect 131460 663270 131570 663510
rect 131810 663270 131900 663510
rect 132140 663270 132230 663510
rect 132470 663270 132560 663510
rect 132800 663270 132910 663510
rect 133150 663270 133170 663510
rect 122170 663180 133170 663270
rect 122170 662940 122190 663180
rect 122430 662940 122520 663180
rect 122760 662940 122850 663180
rect 123090 662940 123180 663180
rect 123420 662940 123530 663180
rect 123770 662940 123860 663180
rect 124100 662940 124190 663180
rect 124430 662940 124520 663180
rect 124760 662940 124870 663180
rect 125110 662940 125200 663180
rect 125440 662940 125530 663180
rect 125770 662940 125860 663180
rect 126100 662940 126210 663180
rect 126450 662940 126540 663180
rect 126780 662940 126870 663180
rect 127110 662940 127200 663180
rect 127440 662940 127550 663180
rect 127790 662940 127880 663180
rect 128120 662940 128210 663180
rect 128450 662940 128540 663180
rect 128780 662940 128890 663180
rect 129130 662940 129220 663180
rect 129460 662940 129550 663180
rect 129790 662940 129880 663180
rect 130120 662940 130230 663180
rect 130470 662940 130560 663180
rect 130800 662940 130890 663180
rect 131130 662940 131220 663180
rect 131460 662940 131570 663180
rect 131810 662940 131900 663180
rect 132140 662940 132230 663180
rect 132470 662940 132560 663180
rect 132800 662940 132910 663180
rect 133150 662940 133170 663180
rect 122170 662850 133170 662940
rect 122170 662610 122190 662850
rect 122430 662610 122520 662850
rect 122760 662610 122850 662850
rect 123090 662610 123180 662850
rect 123420 662610 123530 662850
rect 123770 662610 123860 662850
rect 124100 662610 124190 662850
rect 124430 662610 124520 662850
rect 124760 662610 124870 662850
rect 125110 662610 125200 662850
rect 125440 662610 125530 662850
rect 125770 662610 125860 662850
rect 126100 662610 126210 662850
rect 126450 662610 126540 662850
rect 126780 662610 126870 662850
rect 127110 662610 127200 662850
rect 127440 662610 127550 662850
rect 127790 662610 127880 662850
rect 128120 662610 128210 662850
rect 128450 662610 128540 662850
rect 128780 662610 128890 662850
rect 129130 662610 129220 662850
rect 129460 662610 129550 662850
rect 129790 662610 129880 662850
rect 130120 662610 130230 662850
rect 130470 662610 130560 662850
rect 130800 662610 130890 662850
rect 131130 662610 131220 662850
rect 131460 662610 131570 662850
rect 131810 662610 131900 662850
rect 132140 662610 132230 662850
rect 132470 662610 132560 662850
rect 132800 662610 132910 662850
rect 133150 662610 133170 662850
rect 122170 662520 133170 662610
rect 122170 662280 122190 662520
rect 122430 662280 122520 662520
rect 122760 662280 122850 662520
rect 123090 662280 123180 662520
rect 123420 662280 123530 662520
rect 123770 662280 123860 662520
rect 124100 662280 124190 662520
rect 124430 662280 124520 662520
rect 124760 662280 124870 662520
rect 125110 662280 125200 662520
rect 125440 662280 125530 662520
rect 125770 662280 125860 662520
rect 126100 662280 126210 662520
rect 126450 662280 126540 662520
rect 126780 662280 126870 662520
rect 127110 662280 127200 662520
rect 127440 662280 127550 662520
rect 127790 662280 127880 662520
rect 128120 662280 128210 662520
rect 128450 662280 128540 662520
rect 128780 662280 128890 662520
rect 129130 662280 129220 662520
rect 129460 662280 129550 662520
rect 129790 662280 129880 662520
rect 130120 662280 130230 662520
rect 130470 662280 130560 662520
rect 130800 662280 130890 662520
rect 131130 662280 131220 662520
rect 131460 662280 131570 662520
rect 131810 662280 131900 662520
rect 132140 662280 132230 662520
rect 132470 662280 132560 662520
rect 132800 662280 132910 662520
rect 133150 662280 133170 662520
rect 122170 662170 133170 662280
rect 122170 661930 122190 662170
rect 122430 661930 122520 662170
rect 122760 661930 122850 662170
rect 123090 661930 123180 662170
rect 123420 661930 123530 662170
rect 123770 661930 123860 662170
rect 124100 661930 124190 662170
rect 124430 661930 124520 662170
rect 124760 661930 124870 662170
rect 125110 661930 125200 662170
rect 125440 661930 125530 662170
rect 125770 661930 125860 662170
rect 126100 661930 126210 662170
rect 126450 661930 126540 662170
rect 126780 661930 126870 662170
rect 127110 661930 127200 662170
rect 127440 661930 127550 662170
rect 127790 661930 127880 662170
rect 128120 661930 128210 662170
rect 128450 661930 128540 662170
rect 128780 661930 128890 662170
rect 129130 661930 129220 662170
rect 129460 661930 129550 662170
rect 129790 661930 129880 662170
rect 130120 661930 130230 662170
rect 130470 661930 130560 662170
rect 130800 661930 130890 662170
rect 131130 661930 131220 662170
rect 131460 661930 131570 662170
rect 131810 661930 131900 662170
rect 132140 661930 132230 662170
rect 132470 661930 132560 662170
rect 132800 661930 132910 662170
rect 133150 661930 133170 662170
rect 122170 661840 133170 661930
rect 122170 661600 122190 661840
rect 122430 661600 122520 661840
rect 122760 661600 122850 661840
rect 123090 661600 123180 661840
rect 123420 661600 123530 661840
rect 123770 661600 123860 661840
rect 124100 661600 124190 661840
rect 124430 661600 124520 661840
rect 124760 661600 124870 661840
rect 125110 661600 125200 661840
rect 125440 661600 125530 661840
rect 125770 661600 125860 661840
rect 126100 661600 126210 661840
rect 126450 661600 126540 661840
rect 126780 661600 126870 661840
rect 127110 661600 127200 661840
rect 127440 661600 127550 661840
rect 127790 661600 127880 661840
rect 128120 661600 128210 661840
rect 128450 661600 128540 661840
rect 128780 661600 128890 661840
rect 129130 661600 129220 661840
rect 129460 661600 129550 661840
rect 129790 661600 129880 661840
rect 130120 661600 130230 661840
rect 130470 661600 130560 661840
rect 130800 661600 130890 661840
rect 131130 661600 131220 661840
rect 131460 661600 131570 661840
rect 131810 661600 131900 661840
rect 132140 661600 132230 661840
rect 132470 661600 132560 661840
rect 132800 661600 132910 661840
rect 133150 661600 133170 661840
rect 122170 661510 133170 661600
rect 122170 661270 122190 661510
rect 122430 661270 122520 661510
rect 122760 661270 122850 661510
rect 123090 661270 123180 661510
rect 123420 661270 123530 661510
rect 123770 661270 123860 661510
rect 124100 661270 124190 661510
rect 124430 661270 124520 661510
rect 124760 661270 124870 661510
rect 125110 661270 125200 661510
rect 125440 661270 125530 661510
rect 125770 661270 125860 661510
rect 126100 661270 126210 661510
rect 126450 661270 126540 661510
rect 126780 661270 126870 661510
rect 127110 661270 127200 661510
rect 127440 661270 127550 661510
rect 127790 661270 127880 661510
rect 128120 661270 128210 661510
rect 128450 661270 128540 661510
rect 128780 661270 128890 661510
rect 129130 661270 129220 661510
rect 129460 661270 129550 661510
rect 129790 661270 129880 661510
rect 130120 661270 130230 661510
rect 130470 661270 130560 661510
rect 130800 661270 130890 661510
rect 131130 661270 131220 661510
rect 131460 661270 131570 661510
rect 131810 661270 131900 661510
rect 132140 661270 132230 661510
rect 132470 661270 132560 661510
rect 132800 661270 132910 661510
rect 133150 661270 133170 661510
rect 122170 661180 133170 661270
rect 122170 660940 122190 661180
rect 122430 660940 122520 661180
rect 122760 660940 122850 661180
rect 123090 660940 123180 661180
rect 123420 660940 123530 661180
rect 123770 660940 123860 661180
rect 124100 660940 124190 661180
rect 124430 660940 124520 661180
rect 124760 660940 124870 661180
rect 125110 660940 125200 661180
rect 125440 660940 125530 661180
rect 125770 660940 125860 661180
rect 126100 660940 126210 661180
rect 126450 660940 126540 661180
rect 126780 660940 126870 661180
rect 127110 660940 127200 661180
rect 127440 660940 127550 661180
rect 127790 660940 127880 661180
rect 128120 660940 128210 661180
rect 128450 660940 128540 661180
rect 128780 660940 128890 661180
rect 129130 660940 129220 661180
rect 129460 660940 129550 661180
rect 129790 660940 129880 661180
rect 130120 660940 130230 661180
rect 130470 660940 130560 661180
rect 130800 660940 130890 661180
rect 131130 660940 131220 661180
rect 131460 660940 131570 661180
rect 131810 660940 131900 661180
rect 132140 660940 132230 661180
rect 132470 660940 132560 661180
rect 132800 660940 132910 661180
rect 133150 660940 133170 661180
rect 122170 660920 133170 660940
rect 133550 671900 144550 671920
rect 133550 671660 133570 671900
rect 133810 671660 133900 671900
rect 134140 671660 134230 671900
rect 134470 671660 134560 671900
rect 134800 671660 134910 671900
rect 135150 671660 135240 671900
rect 135480 671660 135570 671900
rect 135810 671660 135900 671900
rect 136140 671660 136250 671900
rect 136490 671660 136580 671900
rect 136820 671660 136910 671900
rect 137150 671660 137240 671900
rect 137480 671660 137590 671900
rect 137830 671660 137920 671900
rect 138160 671660 138250 671900
rect 138490 671660 138580 671900
rect 138820 671660 138930 671900
rect 139170 671660 139260 671900
rect 139500 671660 139590 671900
rect 139830 671660 139920 671900
rect 140160 671660 140270 671900
rect 140510 671660 140600 671900
rect 140840 671660 140930 671900
rect 141170 671660 141260 671900
rect 141500 671660 141610 671900
rect 141850 671660 141940 671900
rect 142180 671660 142270 671900
rect 142510 671660 142600 671900
rect 142840 671660 142950 671900
rect 143190 671660 143280 671900
rect 143520 671660 143610 671900
rect 143850 671660 143940 671900
rect 144180 671660 144290 671900
rect 144530 671660 144550 671900
rect 133550 671550 144550 671660
rect 133550 671310 133570 671550
rect 133810 671310 133900 671550
rect 134140 671310 134230 671550
rect 134470 671310 134560 671550
rect 134800 671310 134910 671550
rect 135150 671310 135240 671550
rect 135480 671310 135570 671550
rect 135810 671310 135900 671550
rect 136140 671310 136250 671550
rect 136490 671310 136580 671550
rect 136820 671310 136910 671550
rect 137150 671310 137240 671550
rect 137480 671310 137590 671550
rect 137830 671310 137920 671550
rect 138160 671310 138250 671550
rect 138490 671310 138580 671550
rect 138820 671310 138930 671550
rect 139170 671310 139260 671550
rect 139500 671310 139590 671550
rect 139830 671310 139920 671550
rect 140160 671310 140270 671550
rect 140510 671310 140600 671550
rect 140840 671310 140930 671550
rect 141170 671310 141260 671550
rect 141500 671310 141610 671550
rect 141850 671310 141940 671550
rect 142180 671310 142270 671550
rect 142510 671310 142600 671550
rect 142840 671310 142950 671550
rect 143190 671310 143280 671550
rect 143520 671310 143610 671550
rect 143850 671310 143940 671550
rect 144180 671310 144290 671550
rect 144530 671310 144550 671550
rect 133550 671220 144550 671310
rect 133550 670980 133570 671220
rect 133810 670980 133900 671220
rect 134140 670980 134230 671220
rect 134470 670980 134560 671220
rect 134800 670980 134910 671220
rect 135150 670980 135240 671220
rect 135480 670980 135570 671220
rect 135810 670980 135900 671220
rect 136140 670980 136250 671220
rect 136490 670980 136580 671220
rect 136820 670980 136910 671220
rect 137150 670980 137240 671220
rect 137480 670980 137590 671220
rect 137830 670980 137920 671220
rect 138160 670980 138250 671220
rect 138490 670980 138580 671220
rect 138820 670980 138930 671220
rect 139170 670980 139260 671220
rect 139500 670980 139590 671220
rect 139830 670980 139920 671220
rect 140160 670980 140270 671220
rect 140510 670980 140600 671220
rect 140840 670980 140930 671220
rect 141170 670980 141260 671220
rect 141500 670980 141610 671220
rect 141850 670980 141940 671220
rect 142180 670980 142270 671220
rect 142510 670980 142600 671220
rect 142840 670980 142950 671220
rect 143190 670980 143280 671220
rect 143520 670980 143610 671220
rect 143850 670980 143940 671220
rect 144180 670980 144290 671220
rect 144530 670980 144550 671220
rect 133550 670890 144550 670980
rect 133550 670650 133570 670890
rect 133810 670650 133900 670890
rect 134140 670650 134230 670890
rect 134470 670650 134560 670890
rect 134800 670650 134910 670890
rect 135150 670650 135240 670890
rect 135480 670650 135570 670890
rect 135810 670650 135900 670890
rect 136140 670650 136250 670890
rect 136490 670650 136580 670890
rect 136820 670650 136910 670890
rect 137150 670650 137240 670890
rect 137480 670650 137590 670890
rect 137830 670650 137920 670890
rect 138160 670650 138250 670890
rect 138490 670650 138580 670890
rect 138820 670650 138930 670890
rect 139170 670650 139260 670890
rect 139500 670650 139590 670890
rect 139830 670650 139920 670890
rect 140160 670650 140270 670890
rect 140510 670650 140600 670890
rect 140840 670650 140930 670890
rect 141170 670650 141260 670890
rect 141500 670650 141610 670890
rect 141850 670650 141940 670890
rect 142180 670650 142270 670890
rect 142510 670650 142600 670890
rect 142840 670650 142950 670890
rect 143190 670650 143280 670890
rect 143520 670650 143610 670890
rect 143850 670650 143940 670890
rect 144180 670650 144290 670890
rect 144530 670650 144550 670890
rect 133550 670560 144550 670650
rect 133550 670320 133570 670560
rect 133810 670320 133900 670560
rect 134140 670320 134230 670560
rect 134470 670320 134560 670560
rect 134800 670320 134910 670560
rect 135150 670320 135240 670560
rect 135480 670320 135570 670560
rect 135810 670320 135900 670560
rect 136140 670320 136250 670560
rect 136490 670320 136580 670560
rect 136820 670320 136910 670560
rect 137150 670320 137240 670560
rect 137480 670320 137590 670560
rect 137830 670320 137920 670560
rect 138160 670320 138250 670560
rect 138490 670320 138580 670560
rect 138820 670320 138930 670560
rect 139170 670320 139260 670560
rect 139500 670320 139590 670560
rect 139830 670320 139920 670560
rect 140160 670320 140270 670560
rect 140510 670320 140600 670560
rect 140840 670320 140930 670560
rect 141170 670320 141260 670560
rect 141500 670320 141610 670560
rect 141850 670320 141940 670560
rect 142180 670320 142270 670560
rect 142510 670320 142600 670560
rect 142840 670320 142950 670560
rect 143190 670320 143280 670560
rect 143520 670320 143610 670560
rect 143850 670320 143940 670560
rect 144180 670320 144290 670560
rect 144530 670320 144550 670560
rect 133550 670210 144550 670320
rect 133550 669970 133570 670210
rect 133810 669970 133900 670210
rect 134140 669970 134230 670210
rect 134470 669970 134560 670210
rect 134800 669970 134910 670210
rect 135150 669970 135240 670210
rect 135480 669970 135570 670210
rect 135810 669970 135900 670210
rect 136140 669970 136250 670210
rect 136490 669970 136580 670210
rect 136820 669970 136910 670210
rect 137150 669970 137240 670210
rect 137480 669970 137590 670210
rect 137830 669970 137920 670210
rect 138160 669970 138250 670210
rect 138490 669970 138580 670210
rect 138820 669970 138930 670210
rect 139170 669970 139260 670210
rect 139500 669970 139590 670210
rect 139830 669970 139920 670210
rect 140160 669970 140270 670210
rect 140510 669970 140600 670210
rect 140840 669970 140930 670210
rect 141170 669970 141260 670210
rect 141500 669970 141610 670210
rect 141850 669970 141940 670210
rect 142180 669970 142270 670210
rect 142510 669970 142600 670210
rect 142840 669970 142950 670210
rect 143190 669970 143280 670210
rect 143520 669970 143610 670210
rect 143850 669970 143940 670210
rect 144180 669970 144290 670210
rect 144530 669970 144550 670210
rect 133550 669880 144550 669970
rect 133550 669640 133570 669880
rect 133810 669640 133900 669880
rect 134140 669640 134230 669880
rect 134470 669640 134560 669880
rect 134800 669640 134910 669880
rect 135150 669640 135240 669880
rect 135480 669640 135570 669880
rect 135810 669640 135900 669880
rect 136140 669640 136250 669880
rect 136490 669640 136580 669880
rect 136820 669640 136910 669880
rect 137150 669640 137240 669880
rect 137480 669640 137590 669880
rect 137830 669640 137920 669880
rect 138160 669640 138250 669880
rect 138490 669640 138580 669880
rect 138820 669640 138930 669880
rect 139170 669640 139260 669880
rect 139500 669640 139590 669880
rect 139830 669640 139920 669880
rect 140160 669640 140270 669880
rect 140510 669640 140600 669880
rect 140840 669640 140930 669880
rect 141170 669640 141260 669880
rect 141500 669640 141610 669880
rect 141850 669640 141940 669880
rect 142180 669640 142270 669880
rect 142510 669640 142600 669880
rect 142840 669640 142950 669880
rect 143190 669640 143280 669880
rect 143520 669640 143610 669880
rect 143850 669640 143940 669880
rect 144180 669640 144290 669880
rect 144530 669640 144550 669880
rect 133550 669550 144550 669640
rect 133550 669310 133570 669550
rect 133810 669310 133900 669550
rect 134140 669310 134230 669550
rect 134470 669310 134560 669550
rect 134800 669310 134910 669550
rect 135150 669310 135240 669550
rect 135480 669310 135570 669550
rect 135810 669310 135900 669550
rect 136140 669310 136250 669550
rect 136490 669310 136580 669550
rect 136820 669310 136910 669550
rect 137150 669310 137240 669550
rect 137480 669310 137590 669550
rect 137830 669310 137920 669550
rect 138160 669310 138250 669550
rect 138490 669310 138580 669550
rect 138820 669310 138930 669550
rect 139170 669310 139260 669550
rect 139500 669310 139590 669550
rect 139830 669310 139920 669550
rect 140160 669310 140270 669550
rect 140510 669310 140600 669550
rect 140840 669310 140930 669550
rect 141170 669310 141260 669550
rect 141500 669310 141610 669550
rect 141850 669310 141940 669550
rect 142180 669310 142270 669550
rect 142510 669310 142600 669550
rect 142840 669310 142950 669550
rect 143190 669310 143280 669550
rect 143520 669310 143610 669550
rect 143850 669310 143940 669550
rect 144180 669310 144290 669550
rect 144530 669310 144550 669550
rect 133550 669220 144550 669310
rect 133550 668980 133570 669220
rect 133810 668980 133900 669220
rect 134140 668980 134230 669220
rect 134470 668980 134560 669220
rect 134800 668980 134910 669220
rect 135150 668980 135240 669220
rect 135480 668980 135570 669220
rect 135810 668980 135900 669220
rect 136140 668980 136250 669220
rect 136490 668980 136580 669220
rect 136820 668980 136910 669220
rect 137150 668980 137240 669220
rect 137480 668980 137590 669220
rect 137830 668980 137920 669220
rect 138160 668980 138250 669220
rect 138490 668980 138580 669220
rect 138820 668980 138930 669220
rect 139170 668980 139260 669220
rect 139500 668980 139590 669220
rect 139830 668980 139920 669220
rect 140160 668980 140270 669220
rect 140510 668980 140600 669220
rect 140840 668980 140930 669220
rect 141170 668980 141260 669220
rect 141500 668980 141610 669220
rect 141850 668980 141940 669220
rect 142180 668980 142270 669220
rect 142510 668980 142600 669220
rect 142840 668980 142950 669220
rect 143190 668980 143280 669220
rect 143520 668980 143610 669220
rect 143850 668980 143940 669220
rect 144180 668980 144290 669220
rect 144530 668980 144550 669220
rect 133550 668870 144550 668980
rect 133550 668630 133570 668870
rect 133810 668630 133900 668870
rect 134140 668630 134230 668870
rect 134470 668630 134560 668870
rect 134800 668630 134910 668870
rect 135150 668630 135240 668870
rect 135480 668630 135570 668870
rect 135810 668630 135900 668870
rect 136140 668630 136250 668870
rect 136490 668630 136580 668870
rect 136820 668630 136910 668870
rect 137150 668630 137240 668870
rect 137480 668630 137590 668870
rect 137830 668630 137920 668870
rect 138160 668630 138250 668870
rect 138490 668630 138580 668870
rect 138820 668630 138930 668870
rect 139170 668630 139260 668870
rect 139500 668630 139590 668870
rect 139830 668630 139920 668870
rect 140160 668630 140270 668870
rect 140510 668630 140600 668870
rect 140840 668630 140930 668870
rect 141170 668630 141260 668870
rect 141500 668630 141610 668870
rect 141850 668630 141940 668870
rect 142180 668630 142270 668870
rect 142510 668630 142600 668870
rect 142840 668630 142950 668870
rect 143190 668630 143280 668870
rect 143520 668630 143610 668870
rect 143850 668630 143940 668870
rect 144180 668630 144290 668870
rect 144530 668630 144550 668870
rect 133550 668540 144550 668630
rect 133550 668300 133570 668540
rect 133810 668300 133900 668540
rect 134140 668300 134230 668540
rect 134470 668300 134560 668540
rect 134800 668300 134910 668540
rect 135150 668300 135240 668540
rect 135480 668300 135570 668540
rect 135810 668300 135900 668540
rect 136140 668300 136250 668540
rect 136490 668300 136580 668540
rect 136820 668300 136910 668540
rect 137150 668300 137240 668540
rect 137480 668300 137590 668540
rect 137830 668300 137920 668540
rect 138160 668300 138250 668540
rect 138490 668300 138580 668540
rect 138820 668300 138930 668540
rect 139170 668300 139260 668540
rect 139500 668300 139590 668540
rect 139830 668300 139920 668540
rect 140160 668300 140270 668540
rect 140510 668300 140600 668540
rect 140840 668300 140930 668540
rect 141170 668300 141260 668540
rect 141500 668300 141610 668540
rect 141850 668300 141940 668540
rect 142180 668300 142270 668540
rect 142510 668300 142600 668540
rect 142840 668300 142950 668540
rect 143190 668300 143280 668540
rect 143520 668300 143610 668540
rect 143850 668300 143940 668540
rect 144180 668300 144290 668540
rect 144530 668300 144550 668540
rect 133550 668210 144550 668300
rect 133550 667970 133570 668210
rect 133810 667970 133900 668210
rect 134140 667970 134230 668210
rect 134470 667970 134560 668210
rect 134800 667970 134910 668210
rect 135150 667970 135240 668210
rect 135480 667970 135570 668210
rect 135810 667970 135900 668210
rect 136140 667970 136250 668210
rect 136490 667970 136580 668210
rect 136820 667970 136910 668210
rect 137150 667970 137240 668210
rect 137480 667970 137590 668210
rect 137830 667970 137920 668210
rect 138160 667970 138250 668210
rect 138490 667970 138580 668210
rect 138820 667970 138930 668210
rect 139170 667970 139260 668210
rect 139500 667970 139590 668210
rect 139830 667970 139920 668210
rect 140160 667970 140270 668210
rect 140510 667970 140600 668210
rect 140840 667970 140930 668210
rect 141170 667970 141260 668210
rect 141500 667970 141610 668210
rect 141850 667970 141940 668210
rect 142180 667970 142270 668210
rect 142510 667970 142600 668210
rect 142840 667970 142950 668210
rect 143190 667970 143280 668210
rect 143520 667970 143610 668210
rect 143850 667970 143940 668210
rect 144180 667970 144290 668210
rect 144530 667970 144550 668210
rect 133550 667880 144550 667970
rect 133550 667640 133570 667880
rect 133810 667640 133900 667880
rect 134140 667640 134230 667880
rect 134470 667640 134560 667880
rect 134800 667640 134910 667880
rect 135150 667640 135240 667880
rect 135480 667640 135570 667880
rect 135810 667640 135900 667880
rect 136140 667640 136250 667880
rect 136490 667640 136580 667880
rect 136820 667640 136910 667880
rect 137150 667640 137240 667880
rect 137480 667640 137590 667880
rect 137830 667640 137920 667880
rect 138160 667640 138250 667880
rect 138490 667640 138580 667880
rect 138820 667640 138930 667880
rect 139170 667640 139260 667880
rect 139500 667640 139590 667880
rect 139830 667640 139920 667880
rect 140160 667640 140270 667880
rect 140510 667640 140600 667880
rect 140840 667640 140930 667880
rect 141170 667640 141260 667880
rect 141500 667640 141610 667880
rect 141850 667640 141940 667880
rect 142180 667640 142270 667880
rect 142510 667640 142600 667880
rect 142840 667640 142950 667880
rect 143190 667640 143280 667880
rect 143520 667640 143610 667880
rect 143850 667640 143940 667880
rect 144180 667640 144290 667880
rect 144530 667640 144550 667880
rect 133550 667530 144550 667640
rect 133550 667290 133570 667530
rect 133810 667290 133900 667530
rect 134140 667290 134230 667530
rect 134470 667290 134560 667530
rect 134800 667290 134910 667530
rect 135150 667290 135240 667530
rect 135480 667290 135570 667530
rect 135810 667290 135900 667530
rect 136140 667290 136250 667530
rect 136490 667290 136580 667530
rect 136820 667290 136910 667530
rect 137150 667290 137240 667530
rect 137480 667290 137590 667530
rect 137830 667290 137920 667530
rect 138160 667290 138250 667530
rect 138490 667290 138580 667530
rect 138820 667290 138930 667530
rect 139170 667290 139260 667530
rect 139500 667290 139590 667530
rect 139830 667290 139920 667530
rect 140160 667290 140270 667530
rect 140510 667290 140600 667530
rect 140840 667290 140930 667530
rect 141170 667290 141260 667530
rect 141500 667290 141610 667530
rect 141850 667290 141940 667530
rect 142180 667290 142270 667530
rect 142510 667290 142600 667530
rect 142840 667290 142950 667530
rect 143190 667290 143280 667530
rect 143520 667290 143610 667530
rect 143850 667290 143940 667530
rect 144180 667290 144290 667530
rect 144530 667290 144550 667530
rect 133550 667200 144550 667290
rect 133550 666960 133570 667200
rect 133810 666960 133900 667200
rect 134140 666960 134230 667200
rect 134470 666960 134560 667200
rect 134800 666960 134910 667200
rect 135150 666960 135240 667200
rect 135480 666960 135570 667200
rect 135810 666960 135900 667200
rect 136140 666960 136250 667200
rect 136490 666960 136580 667200
rect 136820 666960 136910 667200
rect 137150 666960 137240 667200
rect 137480 666960 137590 667200
rect 137830 666960 137920 667200
rect 138160 666960 138250 667200
rect 138490 666960 138580 667200
rect 138820 666960 138930 667200
rect 139170 666960 139260 667200
rect 139500 666960 139590 667200
rect 139830 666960 139920 667200
rect 140160 666960 140270 667200
rect 140510 666960 140600 667200
rect 140840 666960 140930 667200
rect 141170 666960 141260 667200
rect 141500 666960 141610 667200
rect 141850 666960 141940 667200
rect 142180 666960 142270 667200
rect 142510 666960 142600 667200
rect 142840 666960 142950 667200
rect 143190 666960 143280 667200
rect 143520 666960 143610 667200
rect 143850 666960 143940 667200
rect 144180 666960 144290 667200
rect 144530 666960 144550 667200
rect 133550 666870 144550 666960
rect 133550 666630 133570 666870
rect 133810 666630 133900 666870
rect 134140 666630 134230 666870
rect 134470 666630 134560 666870
rect 134800 666630 134910 666870
rect 135150 666630 135240 666870
rect 135480 666630 135570 666870
rect 135810 666630 135900 666870
rect 136140 666630 136250 666870
rect 136490 666630 136580 666870
rect 136820 666630 136910 666870
rect 137150 666630 137240 666870
rect 137480 666630 137590 666870
rect 137830 666630 137920 666870
rect 138160 666630 138250 666870
rect 138490 666630 138580 666870
rect 138820 666630 138930 666870
rect 139170 666630 139260 666870
rect 139500 666630 139590 666870
rect 139830 666630 139920 666870
rect 140160 666630 140270 666870
rect 140510 666630 140600 666870
rect 140840 666630 140930 666870
rect 141170 666630 141260 666870
rect 141500 666630 141610 666870
rect 141850 666630 141940 666870
rect 142180 666630 142270 666870
rect 142510 666630 142600 666870
rect 142840 666630 142950 666870
rect 143190 666630 143280 666870
rect 143520 666630 143610 666870
rect 143850 666630 143940 666870
rect 144180 666630 144290 666870
rect 144530 666630 144550 666870
rect 133550 666540 144550 666630
rect 133550 666300 133570 666540
rect 133810 666300 133900 666540
rect 134140 666300 134230 666540
rect 134470 666300 134560 666540
rect 134800 666300 134910 666540
rect 135150 666300 135240 666540
rect 135480 666300 135570 666540
rect 135810 666300 135900 666540
rect 136140 666300 136250 666540
rect 136490 666300 136580 666540
rect 136820 666300 136910 666540
rect 137150 666300 137240 666540
rect 137480 666300 137590 666540
rect 137830 666300 137920 666540
rect 138160 666300 138250 666540
rect 138490 666300 138580 666540
rect 138820 666300 138930 666540
rect 139170 666300 139260 666540
rect 139500 666300 139590 666540
rect 139830 666300 139920 666540
rect 140160 666300 140270 666540
rect 140510 666300 140600 666540
rect 140840 666300 140930 666540
rect 141170 666300 141260 666540
rect 141500 666300 141610 666540
rect 141850 666300 141940 666540
rect 142180 666300 142270 666540
rect 142510 666300 142600 666540
rect 142840 666300 142950 666540
rect 143190 666300 143280 666540
rect 143520 666300 143610 666540
rect 143850 666300 143940 666540
rect 144180 666300 144290 666540
rect 144530 666300 144550 666540
rect 133550 666190 144550 666300
rect 133550 665950 133570 666190
rect 133810 665950 133900 666190
rect 134140 665950 134230 666190
rect 134470 665950 134560 666190
rect 134800 665950 134910 666190
rect 135150 665950 135240 666190
rect 135480 665950 135570 666190
rect 135810 665950 135900 666190
rect 136140 665950 136250 666190
rect 136490 665950 136580 666190
rect 136820 665950 136910 666190
rect 137150 665950 137240 666190
rect 137480 665950 137590 666190
rect 137830 665950 137920 666190
rect 138160 665950 138250 666190
rect 138490 665950 138580 666190
rect 138820 665950 138930 666190
rect 139170 665950 139260 666190
rect 139500 665950 139590 666190
rect 139830 665950 139920 666190
rect 140160 665950 140270 666190
rect 140510 665950 140600 666190
rect 140840 665950 140930 666190
rect 141170 665950 141260 666190
rect 141500 665950 141610 666190
rect 141850 665950 141940 666190
rect 142180 665950 142270 666190
rect 142510 665950 142600 666190
rect 142840 665950 142950 666190
rect 143190 665950 143280 666190
rect 143520 665950 143610 666190
rect 143850 665950 143940 666190
rect 144180 665950 144290 666190
rect 144530 665950 144550 666190
rect 133550 665860 144550 665950
rect 133550 665620 133570 665860
rect 133810 665620 133900 665860
rect 134140 665620 134230 665860
rect 134470 665620 134560 665860
rect 134800 665620 134910 665860
rect 135150 665620 135240 665860
rect 135480 665620 135570 665860
rect 135810 665620 135900 665860
rect 136140 665620 136250 665860
rect 136490 665620 136580 665860
rect 136820 665620 136910 665860
rect 137150 665620 137240 665860
rect 137480 665620 137590 665860
rect 137830 665620 137920 665860
rect 138160 665620 138250 665860
rect 138490 665620 138580 665860
rect 138820 665620 138930 665860
rect 139170 665620 139260 665860
rect 139500 665620 139590 665860
rect 139830 665620 139920 665860
rect 140160 665620 140270 665860
rect 140510 665620 140600 665860
rect 140840 665620 140930 665860
rect 141170 665620 141260 665860
rect 141500 665620 141610 665860
rect 141850 665620 141940 665860
rect 142180 665620 142270 665860
rect 142510 665620 142600 665860
rect 142840 665620 142950 665860
rect 143190 665620 143280 665860
rect 143520 665620 143610 665860
rect 143850 665620 143940 665860
rect 144180 665620 144290 665860
rect 144530 665620 144550 665860
rect 133550 665530 144550 665620
rect 133550 665290 133570 665530
rect 133810 665290 133900 665530
rect 134140 665290 134230 665530
rect 134470 665290 134560 665530
rect 134800 665290 134910 665530
rect 135150 665290 135240 665530
rect 135480 665290 135570 665530
rect 135810 665290 135900 665530
rect 136140 665290 136250 665530
rect 136490 665290 136580 665530
rect 136820 665290 136910 665530
rect 137150 665290 137240 665530
rect 137480 665290 137590 665530
rect 137830 665290 137920 665530
rect 138160 665290 138250 665530
rect 138490 665290 138580 665530
rect 138820 665290 138930 665530
rect 139170 665290 139260 665530
rect 139500 665290 139590 665530
rect 139830 665290 139920 665530
rect 140160 665290 140270 665530
rect 140510 665290 140600 665530
rect 140840 665290 140930 665530
rect 141170 665290 141260 665530
rect 141500 665290 141610 665530
rect 141850 665290 141940 665530
rect 142180 665290 142270 665530
rect 142510 665290 142600 665530
rect 142840 665290 142950 665530
rect 143190 665290 143280 665530
rect 143520 665290 143610 665530
rect 143850 665290 143940 665530
rect 144180 665290 144290 665530
rect 144530 665290 144550 665530
rect 133550 665200 144550 665290
rect 133550 664960 133570 665200
rect 133810 664960 133900 665200
rect 134140 664960 134230 665200
rect 134470 664960 134560 665200
rect 134800 664960 134910 665200
rect 135150 664960 135240 665200
rect 135480 664960 135570 665200
rect 135810 664960 135900 665200
rect 136140 664960 136250 665200
rect 136490 664960 136580 665200
rect 136820 664960 136910 665200
rect 137150 664960 137240 665200
rect 137480 664960 137590 665200
rect 137830 664960 137920 665200
rect 138160 664960 138250 665200
rect 138490 664960 138580 665200
rect 138820 664960 138930 665200
rect 139170 664960 139260 665200
rect 139500 664960 139590 665200
rect 139830 664960 139920 665200
rect 140160 664960 140270 665200
rect 140510 664960 140600 665200
rect 140840 664960 140930 665200
rect 141170 664960 141260 665200
rect 141500 664960 141610 665200
rect 141850 664960 141940 665200
rect 142180 664960 142270 665200
rect 142510 664960 142600 665200
rect 142840 664960 142950 665200
rect 143190 664960 143280 665200
rect 143520 664960 143610 665200
rect 143850 664960 143940 665200
rect 144180 664960 144290 665200
rect 144530 664960 144550 665200
rect 133550 664850 144550 664960
rect 133550 664610 133570 664850
rect 133810 664610 133900 664850
rect 134140 664610 134230 664850
rect 134470 664610 134560 664850
rect 134800 664610 134910 664850
rect 135150 664610 135240 664850
rect 135480 664610 135570 664850
rect 135810 664610 135900 664850
rect 136140 664610 136250 664850
rect 136490 664610 136580 664850
rect 136820 664610 136910 664850
rect 137150 664610 137240 664850
rect 137480 664610 137590 664850
rect 137830 664610 137920 664850
rect 138160 664610 138250 664850
rect 138490 664610 138580 664850
rect 138820 664610 138930 664850
rect 139170 664610 139260 664850
rect 139500 664610 139590 664850
rect 139830 664610 139920 664850
rect 140160 664610 140270 664850
rect 140510 664610 140600 664850
rect 140840 664610 140930 664850
rect 141170 664610 141260 664850
rect 141500 664610 141610 664850
rect 141850 664610 141940 664850
rect 142180 664610 142270 664850
rect 142510 664610 142600 664850
rect 142840 664610 142950 664850
rect 143190 664610 143280 664850
rect 143520 664610 143610 664850
rect 143850 664610 143940 664850
rect 144180 664610 144290 664850
rect 144530 664610 144550 664850
rect 133550 664520 144550 664610
rect 133550 664280 133570 664520
rect 133810 664280 133900 664520
rect 134140 664280 134230 664520
rect 134470 664280 134560 664520
rect 134800 664280 134910 664520
rect 135150 664280 135240 664520
rect 135480 664280 135570 664520
rect 135810 664280 135900 664520
rect 136140 664280 136250 664520
rect 136490 664280 136580 664520
rect 136820 664280 136910 664520
rect 137150 664280 137240 664520
rect 137480 664280 137590 664520
rect 137830 664280 137920 664520
rect 138160 664280 138250 664520
rect 138490 664280 138580 664520
rect 138820 664280 138930 664520
rect 139170 664280 139260 664520
rect 139500 664280 139590 664520
rect 139830 664280 139920 664520
rect 140160 664280 140270 664520
rect 140510 664280 140600 664520
rect 140840 664280 140930 664520
rect 141170 664280 141260 664520
rect 141500 664280 141610 664520
rect 141850 664280 141940 664520
rect 142180 664280 142270 664520
rect 142510 664280 142600 664520
rect 142840 664280 142950 664520
rect 143190 664280 143280 664520
rect 143520 664280 143610 664520
rect 143850 664280 143940 664520
rect 144180 664280 144290 664520
rect 144530 664280 144550 664520
rect 133550 664190 144550 664280
rect 133550 663950 133570 664190
rect 133810 663950 133900 664190
rect 134140 663950 134230 664190
rect 134470 663950 134560 664190
rect 134800 663950 134910 664190
rect 135150 663950 135240 664190
rect 135480 663950 135570 664190
rect 135810 663950 135900 664190
rect 136140 663950 136250 664190
rect 136490 663950 136580 664190
rect 136820 663950 136910 664190
rect 137150 663950 137240 664190
rect 137480 663950 137590 664190
rect 137830 663950 137920 664190
rect 138160 663950 138250 664190
rect 138490 663950 138580 664190
rect 138820 663950 138930 664190
rect 139170 663950 139260 664190
rect 139500 663950 139590 664190
rect 139830 663950 139920 664190
rect 140160 663950 140270 664190
rect 140510 663950 140600 664190
rect 140840 663950 140930 664190
rect 141170 663950 141260 664190
rect 141500 663950 141610 664190
rect 141850 663950 141940 664190
rect 142180 663950 142270 664190
rect 142510 663950 142600 664190
rect 142840 663950 142950 664190
rect 143190 663950 143280 664190
rect 143520 663950 143610 664190
rect 143850 663950 143940 664190
rect 144180 663950 144290 664190
rect 144530 663950 144550 664190
rect 133550 663860 144550 663950
rect 133550 663620 133570 663860
rect 133810 663620 133900 663860
rect 134140 663620 134230 663860
rect 134470 663620 134560 663860
rect 134800 663620 134910 663860
rect 135150 663620 135240 663860
rect 135480 663620 135570 663860
rect 135810 663620 135900 663860
rect 136140 663620 136250 663860
rect 136490 663620 136580 663860
rect 136820 663620 136910 663860
rect 137150 663620 137240 663860
rect 137480 663620 137590 663860
rect 137830 663620 137920 663860
rect 138160 663620 138250 663860
rect 138490 663620 138580 663860
rect 138820 663620 138930 663860
rect 139170 663620 139260 663860
rect 139500 663620 139590 663860
rect 139830 663620 139920 663860
rect 140160 663620 140270 663860
rect 140510 663620 140600 663860
rect 140840 663620 140930 663860
rect 141170 663620 141260 663860
rect 141500 663620 141610 663860
rect 141850 663620 141940 663860
rect 142180 663620 142270 663860
rect 142510 663620 142600 663860
rect 142840 663620 142950 663860
rect 143190 663620 143280 663860
rect 143520 663620 143610 663860
rect 143850 663620 143940 663860
rect 144180 663620 144290 663860
rect 144530 663620 144550 663860
rect 133550 663510 144550 663620
rect 133550 663270 133570 663510
rect 133810 663270 133900 663510
rect 134140 663270 134230 663510
rect 134470 663270 134560 663510
rect 134800 663270 134910 663510
rect 135150 663270 135240 663510
rect 135480 663270 135570 663510
rect 135810 663270 135900 663510
rect 136140 663270 136250 663510
rect 136490 663270 136580 663510
rect 136820 663270 136910 663510
rect 137150 663270 137240 663510
rect 137480 663270 137590 663510
rect 137830 663270 137920 663510
rect 138160 663270 138250 663510
rect 138490 663270 138580 663510
rect 138820 663270 138930 663510
rect 139170 663270 139260 663510
rect 139500 663270 139590 663510
rect 139830 663270 139920 663510
rect 140160 663270 140270 663510
rect 140510 663270 140600 663510
rect 140840 663270 140930 663510
rect 141170 663270 141260 663510
rect 141500 663270 141610 663510
rect 141850 663270 141940 663510
rect 142180 663270 142270 663510
rect 142510 663270 142600 663510
rect 142840 663270 142950 663510
rect 143190 663270 143280 663510
rect 143520 663270 143610 663510
rect 143850 663270 143940 663510
rect 144180 663270 144290 663510
rect 144530 663270 144550 663510
rect 133550 663180 144550 663270
rect 133550 662940 133570 663180
rect 133810 662940 133900 663180
rect 134140 662940 134230 663180
rect 134470 662940 134560 663180
rect 134800 662940 134910 663180
rect 135150 662940 135240 663180
rect 135480 662940 135570 663180
rect 135810 662940 135900 663180
rect 136140 662940 136250 663180
rect 136490 662940 136580 663180
rect 136820 662940 136910 663180
rect 137150 662940 137240 663180
rect 137480 662940 137590 663180
rect 137830 662940 137920 663180
rect 138160 662940 138250 663180
rect 138490 662940 138580 663180
rect 138820 662940 138930 663180
rect 139170 662940 139260 663180
rect 139500 662940 139590 663180
rect 139830 662940 139920 663180
rect 140160 662940 140270 663180
rect 140510 662940 140600 663180
rect 140840 662940 140930 663180
rect 141170 662940 141260 663180
rect 141500 662940 141610 663180
rect 141850 662940 141940 663180
rect 142180 662940 142270 663180
rect 142510 662940 142600 663180
rect 142840 662940 142950 663180
rect 143190 662940 143280 663180
rect 143520 662940 143610 663180
rect 143850 662940 143940 663180
rect 144180 662940 144290 663180
rect 144530 662940 144550 663180
rect 133550 662850 144550 662940
rect 133550 662610 133570 662850
rect 133810 662610 133900 662850
rect 134140 662610 134230 662850
rect 134470 662610 134560 662850
rect 134800 662610 134910 662850
rect 135150 662610 135240 662850
rect 135480 662610 135570 662850
rect 135810 662610 135900 662850
rect 136140 662610 136250 662850
rect 136490 662610 136580 662850
rect 136820 662610 136910 662850
rect 137150 662610 137240 662850
rect 137480 662610 137590 662850
rect 137830 662610 137920 662850
rect 138160 662610 138250 662850
rect 138490 662610 138580 662850
rect 138820 662610 138930 662850
rect 139170 662610 139260 662850
rect 139500 662610 139590 662850
rect 139830 662610 139920 662850
rect 140160 662610 140270 662850
rect 140510 662610 140600 662850
rect 140840 662610 140930 662850
rect 141170 662610 141260 662850
rect 141500 662610 141610 662850
rect 141850 662610 141940 662850
rect 142180 662610 142270 662850
rect 142510 662610 142600 662850
rect 142840 662610 142950 662850
rect 143190 662610 143280 662850
rect 143520 662610 143610 662850
rect 143850 662610 143940 662850
rect 144180 662610 144290 662850
rect 144530 662610 144550 662850
rect 133550 662520 144550 662610
rect 133550 662280 133570 662520
rect 133810 662280 133900 662520
rect 134140 662280 134230 662520
rect 134470 662280 134560 662520
rect 134800 662280 134910 662520
rect 135150 662280 135240 662520
rect 135480 662280 135570 662520
rect 135810 662280 135900 662520
rect 136140 662280 136250 662520
rect 136490 662280 136580 662520
rect 136820 662280 136910 662520
rect 137150 662280 137240 662520
rect 137480 662280 137590 662520
rect 137830 662280 137920 662520
rect 138160 662280 138250 662520
rect 138490 662280 138580 662520
rect 138820 662280 138930 662520
rect 139170 662280 139260 662520
rect 139500 662280 139590 662520
rect 139830 662280 139920 662520
rect 140160 662280 140270 662520
rect 140510 662280 140600 662520
rect 140840 662280 140930 662520
rect 141170 662280 141260 662520
rect 141500 662280 141610 662520
rect 141850 662280 141940 662520
rect 142180 662280 142270 662520
rect 142510 662280 142600 662520
rect 142840 662280 142950 662520
rect 143190 662280 143280 662520
rect 143520 662280 143610 662520
rect 143850 662280 143940 662520
rect 144180 662280 144290 662520
rect 144530 662280 144550 662520
rect 133550 662170 144550 662280
rect 133550 661930 133570 662170
rect 133810 661930 133900 662170
rect 134140 661930 134230 662170
rect 134470 661930 134560 662170
rect 134800 661930 134910 662170
rect 135150 661930 135240 662170
rect 135480 661930 135570 662170
rect 135810 661930 135900 662170
rect 136140 661930 136250 662170
rect 136490 661930 136580 662170
rect 136820 661930 136910 662170
rect 137150 661930 137240 662170
rect 137480 661930 137590 662170
rect 137830 661930 137920 662170
rect 138160 661930 138250 662170
rect 138490 661930 138580 662170
rect 138820 661930 138930 662170
rect 139170 661930 139260 662170
rect 139500 661930 139590 662170
rect 139830 661930 139920 662170
rect 140160 661930 140270 662170
rect 140510 661930 140600 662170
rect 140840 661930 140930 662170
rect 141170 661930 141260 662170
rect 141500 661930 141610 662170
rect 141850 661930 141940 662170
rect 142180 661930 142270 662170
rect 142510 661930 142600 662170
rect 142840 661930 142950 662170
rect 143190 661930 143280 662170
rect 143520 661930 143610 662170
rect 143850 661930 143940 662170
rect 144180 661930 144290 662170
rect 144530 661930 144550 662170
rect 133550 661840 144550 661930
rect 133550 661600 133570 661840
rect 133810 661600 133900 661840
rect 134140 661600 134230 661840
rect 134470 661600 134560 661840
rect 134800 661600 134910 661840
rect 135150 661600 135240 661840
rect 135480 661600 135570 661840
rect 135810 661600 135900 661840
rect 136140 661600 136250 661840
rect 136490 661600 136580 661840
rect 136820 661600 136910 661840
rect 137150 661600 137240 661840
rect 137480 661600 137590 661840
rect 137830 661600 137920 661840
rect 138160 661600 138250 661840
rect 138490 661600 138580 661840
rect 138820 661600 138930 661840
rect 139170 661600 139260 661840
rect 139500 661600 139590 661840
rect 139830 661600 139920 661840
rect 140160 661600 140270 661840
rect 140510 661600 140600 661840
rect 140840 661600 140930 661840
rect 141170 661600 141260 661840
rect 141500 661600 141610 661840
rect 141850 661600 141940 661840
rect 142180 661600 142270 661840
rect 142510 661600 142600 661840
rect 142840 661600 142950 661840
rect 143190 661600 143280 661840
rect 143520 661600 143610 661840
rect 143850 661600 143940 661840
rect 144180 661600 144290 661840
rect 144530 661600 144550 661840
rect 133550 661510 144550 661600
rect 133550 661270 133570 661510
rect 133810 661270 133900 661510
rect 134140 661270 134230 661510
rect 134470 661270 134560 661510
rect 134800 661270 134910 661510
rect 135150 661270 135240 661510
rect 135480 661270 135570 661510
rect 135810 661270 135900 661510
rect 136140 661270 136250 661510
rect 136490 661270 136580 661510
rect 136820 661270 136910 661510
rect 137150 661270 137240 661510
rect 137480 661270 137590 661510
rect 137830 661270 137920 661510
rect 138160 661270 138250 661510
rect 138490 661270 138580 661510
rect 138820 661270 138930 661510
rect 139170 661270 139260 661510
rect 139500 661270 139590 661510
rect 139830 661270 139920 661510
rect 140160 661270 140270 661510
rect 140510 661270 140600 661510
rect 140840 661270 140930 661510
rect 141170 661270 141260 661510
rect 141500 661270 141610 661510
rect 141850 661270 141940 661510
rect 142180 661270 142270 661510
rect 142510 661270 142600 661510
rect 142840 661270 142950 661510
rect 143190 661270 143280 661510
rect 143520 661270 143610 661510
rect 143850 661270 143940 661510
rect 144180 661270 144290 661510
rect 144530 661270 144550 661510
rect 133550 661180 144550 661270
rect 133550 660940 133570 661180
rect 133810 660940 133900 661180
rect 134140 660940 134230 661180
rect 134470 660940 134560 661180
rect 134800 660940 134910 661180
rect 135150 660940 135240 661180
rect 135480 660940 135570 661180
rect 135810 660940 135900 661180
rect 136140 660940 136250 661180
rect 136490 660940 136580 661180
rect 136820 660940 136910 661180
rect 137150 660940 137240 661180
rect 137480 660940 137590 661180
rect 137830 660940 137920 661180
rect 138160 660940 138250 661180
rect 138490 660940 138580 661180
rect 138820 660940 138930 661180
rect 139170 660940 139260 661180
rect 139500 660940 139590 661180
rect 139830 660940 139920 661180
rect 140160 660940 140270 661180
rect 140510 660940 140600 661180
rect 140840 660940 140930 661180
rect 141170 660940 141260 661180
rect 141500 660940 141610 661180
rect 141850 660940 141940 661180
rect 142180 660940 142270 661180
rect 142510 660940 142600 661180
rect 142840 660940 142950 661180
rect 143190 660940 143280 661180
rect 143520 660940 143610 661180
rect 143850 660940 143940 661180
rect 144180 660940 144290 661180
rect 144530 660940 144550 661180
rect 133550 660920 144550 660940
rect 144930 671900 155930 671920
rect 144930 671660 144950 671900
rect 145190 671660 145280 671900
rect 145520 671660 145610 671900
rect 145850 671660 145940 671900
rect 146180 671660 146290 671900
rect 146530 671660 146620 671900
rect 146860 671660 146950 671900
rect 147190 671660 147280 671900
rect 147520 671660 147630 671900
rect 147870 671660 147960 671900
rect 148200 671660 148290 671900
rect 148530 671660 148620 671900
rect 148860 671660 148970 671900
rect 149210 671660 149300 671900
rect 149540 671660 149630 671900
rect 149870 671660 149960 671900
rect 150200 671660 150310 671900
rect 150550 671660 150640 671900
rect 150880 671660 150970 671900
rect 151210 671660 151300 671900
rect 151540 671660 151650 671900
rect 151890 671660 151980 671900
rect 152220 671660 152310 671900
rect 152550 671660 152640 671900
rect 152880 671660 152990 671900
rect 153230 671660 153320 671900
rect 153560 671660 153650 671900
rect 153890 671660 153980 671900
rect 154220 671660 154330 671900
rect 154570 671660 154660 671900
rect 154900 671660 154990 671900
rect 155230 671660 155320 671900
rect 155560 671660 155670 671900
rect 155910 671660 155930 671900
rect 144930 671550 155930 671660
rect 144930 671310 144950 671550
rect 145190 671310 145280 671550
rect 145520 671310 145610 671550
rect 145850 671310 145940 671550
rect 146180 671310 146290 671550
rect 146530 671310 146620 671550
rect 146860 671310 146950 671550
rect 147190 671310 147280 671550
rect 147520 671310 147630 671550
rect 147870 671310 147960 671550
rect 148200 671310 148290 671550
rect 148530 671310 148620 671550
rect 148860 671310 148970 671550
rect 149210 671310 149300 671550
rect 149540 671310 149630 671550
rect 149870 671310 149960 671550
rect 150200 671310 150310 671550
rect 150550 671310 150640 671550
rect 150880 671310 150970 671550
rect 151210 671310 151300 671550
rect 151540 671310 151650 671550
rect 151890 671310 151980 671550
rect 152220 671310 152310 671550
rect 152550 671310 152640 671550
rect 152880 671310 152990 671550
rect 153230 671310 153320 671550
rect 153560 671310 153650 671550
rect 153890 671310 153980 671550
rect 154220 671310 154330 671550
rect 154570 671310 154660 671550
rect 154900 671310 154990 671550
rect 155230 671310 155320 671550
rect 155560 671310 155670 671550
rect 155910 671310 155930 671550
rect 144930 671220 155930 671310
rect 144930 670980 144950 671220
rect 145190 670980 145280 671220
rect 145520 670980 145610 671220
rect 145850 670980 145940 671220
rect 146180 670980 146290 671220
rect 146530 670980 146620 671220
rect 146860 670980 146950 671220
rect 147190 670980 147280 671220
rect 147520 670980 147630 671220
rect 147870 670980 147960 671220
rect 148200 670980 148290 671220
rect 148530 670980 148620 671220
rect 148860 670980 148970 671220
rect 149210 670980 149300 671220
rect 149540 670980 149630 671220
rect 149870 670980 149960 671220
rect 150200 670980 150310 671220
rect 150550 670980 150640 671220
rect 150880 670980 150970 671220
rect 151210 670980 151300 671220
rect 151540 670980 151650 671220
rect 151890 670980 151980 671220
rect 152220 670980 152310 671220
rect 152550 670980 152640 671220
rect 152880 670980 152990 671220
rect 153230 670980 153320 671220
rect 153560 670980 153650 671220
rect 153890 670980 153980 671220
rect 154220 670980 154330 671220
rect 154570 670980 154660 671220
rect 154900 670980 154990 671220
rect 155230 670980 155320 671220
rect 155560 670980 155670 671220
rect 155910 670980 155930 671220
rect 144930 670890 155930 670980
rect 144930 670650 144950 670890
rect 145190 670650 145280 670890
rect 145520 670650 145610 670890
rect 145850 670650 145940 670890
rect 146180 670650 146290 670890
rect 146530 670650 146620 670890
rect 146860 670650 146950 670890
rect 147190 670650 147280 670890
rect 147520 670650 147630 670890
rect 147870 670650 147960 670890
rect 148200 670650 148290 670890
rect 148530 670650 148620 670890
rect 148860 670650 148970 670890
rect 149210 670650 149300 670890
rect 149540 670650 149630 670890
rect 149870 670650 149960 670890
rect 150200 670650 150310 670890
rect 150550 670650 150640 670890
rect 150880 670650 150970 670890
rect 151210 670650 151300 670890
rect 151540 670650 151650 670890
rect 151890 670650 151980 670890
rect 152220 670650 152310 670890
rect 152550 670650 152640 670890
rect 152880 670650 152990 670890
rect 153230 670650 153320 670890
rect 153560 670650 153650 670890
rect 153890 670650 153980 670890
rect 154220 670650 154330 670890
rect 154570 670650 154660 670890
rect 154900 670650 154990 670890
rect 155230 670650 155320 670890
rect 155560 670650 155670 670890
rect 155910 670650 155930 670890
rect 144930 670560 155930 670650
rect 144930 670320 144950 670560
rect 145190 670320 145280 670560
rect 145520 670320 145610 670560
rect 145850 670320 145940 670560
rect 146180 670320 146290 670560
rect 146530 670320 146620 670560
rect 146860 670320 146950 670560
rect 147190 670320 147280 670560
rect 147520 670320 147630 670560
rect 147870 670320 147960 670560
rect 148200 670320 148290 670560
rect 148530 670320 148620 670560
rect 148860 670320 148970 670560
rect 149210 670320 149300 670560
rect 149540 670320 149630 670560
rect 149870 670320 149960 670560
rect 150200 670320 150310 670560
rect 150550 670320 150640 670560
rect 150880 670320 150970 670560
rect 151210 670320 151300 670560
rect 151540 670320 151650 670560
rect 151890 670320 151980 670560
rect 152220 670320 152310 670560
rect 152550 670320 152640 670560
rect 152880 670320 152990 670560
rect 153230 670320 153320 670560
rect 153560 670320 153650 670560
rect 153890 670320 153980 670560
rect 154220 670320 154330 670560
rect 154570 670320 154660 670560
rect 154900 670320 154990 670560
rect 155230 670320 155320 670560
rect 155560 670320 155670 670560
rect 155910 670320 155930 670560
rect 144930 670210 155930 670320
rect 144930 669970 144950 670210
rect 145190 669970 145280 670210
rect 145520 669970 145610 670210
rect 145850 669970 145940 670210
rect 146180 669970 146290 670210
rect 146530 669970 146620 670210
rect 146860 669970 146950 670210
rect 147190 669970 147280 670210
rect 147520 669970 147630 670210
rect 147870 669970 147960 670210
rect 148200 669970 148290 670210
rect 148530 669970 148620 670210
rect 148860 669970 148970 670210
rect 149210 669970 149300 670210
rect 149540 669970 149630 670210
rect 149870 669970 149960 670210
rect 150200 669970 150310 670210
rect 150550 669970 150640 670210
rect 150880 669970 150970 670210
rect 151210 669970 151300 670210
rect 151540 669970 151650 670210
rect 151890 669970 151980 670210
rect 152220 669970 152310 670210
rect 152550 669970 152640 670210
rect 152880 669970 152990 670210
rect 153230 669970 153320 670210
rect 153560 669970 153650 670210
rect 153890 669970 153980 670210
rect 154220 669970 154330 670210
rect 154570 669970 154660 670210
rect 154900 669970 154990 670210
rect 155230 669970 155320 670210
rect 155560 669970 155670 670210
rect 155910 669970 155930 670210
rect 144930 669880 155930 669970
rect 144930 669640 144950 669880
rect 145190 669640 145280 669880
rect 145520 669640 145610 669880
rect 145850 669640 145940 669880
rect 146180 669640 146290 669880
rect 146530 669640 146620 669880
rect 146860 669640 146950 669880
rect 147190 669640 147280 669880
rect 147520 669640 147630 669880
rect 147870 669640 147960 669880
rect 148200 669640 148290 669880
rect 148530 669640 148620 669880
rect 148860 669640 148970 669880
rect 149210 669640 149300 669880
rect 149540 669640 149630 669880
rect 149870 669640 149960 669880
rect 150200 669640 150310 669880
rect 150550 669640 150640 669880
rect 150880 669640 150970 669880
rect 151210 669640 151300 669880
rect 151540 669640 151650 669880
rect 151890 669640 151980 669880
rect 152220 669640 152310 669880
rect 152550 669640 152640 669880
rect 152880 669640 152990 669880
rect 153230 669640 153320 669880
rect 153560 669640 153650 669880
rect 153890 669640 153980 669880
rect 154220 669640 154330 669880
rect 154570 669640 154660 669880
rect 154900 669640 154990 669880
rect 155230 669640 155320 669880
rect 155560 669640 155670 669880
rect 155910 669640 155930 669880
rect 144930 669550 155930 669640
rect 144930 669310 144950 669550
rect 145190 669310 145280 669550
rect 145520 669310 145610 669550
rect 145850 669310 145940 669550
rect 146180 669310 146290 669550
rect 146530 669310 146620 669550
rect 146860 669310 146950 669550
rect 147190 669310 147280 669550
rect 147520 669310 147630 669550
rect 147870 669310 147960 669550
rect 148200 669310 148290 669550
rect 148530 669310 148620 669550
rect 148860 669310 148970 669550
rect 149210 669310 149300 669550
rect 149540 669310 149630 669550
rect 149870 669310 149960 669550
rect 150200 669310 150310 669550
rect 150550 669310 150640 669550
rect 150880 669310 150970 669550
rect 151210 669310 151300 669550
rect 151540 669310 151650 669550
rect 151890 669310 151980 669550
rect 152220 669310 152310 669550
rect 152550 669310 152640 669550
rect 152880 669310 152990 669550
rect 153230 669310 153320 669550
rect 153560 669310 153650 669550
rect 153890 669310 153980 669550
rect 154220 669310 154330 669550
rect 154570 669310 154660 669550
rect 154900 669310 154990 669550
rect 155230 669310 155320 669550
rect 155560 669310 155670 669550
rect 155910 669310 155930 669550
rect 144930 669220 155930 669310
rect 144930 668980 144950 669220
rect 145190 668980 145280 669220
rect 145520 668980 145610 669220
rect 145850 668980 145940 669220
rect 146180 668980 146290 669220
rect 146530 668980 146620 669220
rect 146860 668980 146950 669220
rect 147190 668980 147280 669220
rect 147520 668980 147630 669220
rect 147870 668980 147960 669220
rect 148200 668980 148290 669220
rect 148530 668980 148620 669220
rect 148860 668980 148970 669220
rect 149210 668980 149300 669220
rect 149540 668980 149630 669220
rect 149870 668980 149960 669220
rect 150200 668980 150310 669220
rect 150550 668980 150640 669220
rect 150880 668980 150970 669220
rect 151210 668980 151300 669220
rect 151540 668980 151650 669220
rect 151890 668980 151980 669220
rect 152220 668980 152310 669220
rect 152550 668980 152640 669220
rect 152880 668980 152990 669220
rect 153230 668980 153320 669220
rect 153560 668980 153650 669220
rect 153890 668980 153980 669220
rect 154220 668980 154330 669220
rect 154570 668980 154660 669220
rect 154900 668980 154990 669220
rect 155230 668980 155320 669220
rect 155560 668980 155670 669220
rect 155910 668980 155930 669220
rect 144930 668870 155930 668980
rect 144930 668630 144950 668870
rect 145190 668630 145280 668870
rect 145520 668630 145610 668870
rect 145850 668630 145940 668870
rect 146180 668630 146290 668870
rect 146530 668630 146620 668870
rect 146860 668630 146950 668870
rect 147190 668630 147280 668870
rect 147520 668630 147630 668870
rect 147870 668630 147960 668870
rect 148200 668630 148290 668870
rect 148530 668630 148620 668870
rect 148860 668630 148970 668870
rect 149210 668630 149300 668870
rect 149540 668630 149630 668870
rect 149870 668630 149960 668870
rect 150200 668630 150310 668870
rect 150550 668630 150640 668870
rect 150880 668630 150970 668870
rect 151210 668630 151300 668870
rect 151540 668630 151650 668870
rect 151890 668630 151980 668870
rect 152220 668630 152310 668870
rect 152550 668630 152640 668870
rect 152880 668630 152990 668870
rect 153230 668630 153320 668870
rect 153560 668630 153650 668870
rect 153890 668630 153980 668870
rect 154220 668630 154330 668870
rect 154570 668630 154660 668870
rect 154900 668630 154990 668870
rect 155230 668630 155320 668870
rect 155560 668630 155670 668870
rect 155910 668630 155930 668870
rect 144930 668540 155930 668630
rect 144930 668300 144950 668540
rect 145190 668300 145280 668540
rect 145520 668300 145610 668540
rect 145850 668300 145940 668540
rect 146180 668300 146290 668540
rect 146530 668300 146620 668540
rect 146860 668300 146950 668540
rect 147190 668300 147280 668540
rect 147520 668300 147630 668540
rect 147870 668300 147960 668540
rect 148200 668300 148290 668540
rect 148530 668300 148620 668540
rect 148860 668300 148970 668540
rect 149210 668300 149300 668540
rect 149540 668300 149630 668540
rect 149870 668300 149960 668540
rect 150200 668300 150310 668540
rect 150550 668300 150640 668540
rect 150880 668300 150970 668540
rect 151210 668300 151300 668540
rect 151540 668300 151650 668540
rect 151890 668300 151980 668540
rect 152220 668300 152310 668540
rect 152550 668300 152640 668540
rect 152880 668300 152990 668540
rect 153230 668300 153320 668540
rect 153560 668300 153650 668540
rect 153890 668300 153980 668540
rect 154220 668300 154330 668540
rect 154570 668300 154660 668540
rect 154900 668300 154990 668540
rect 155230 668300 155320 668540
rect 155560 668300 155670 668540
rect 155910 668300 155930 668540
rect 144930 668210 155930 668300
rect 144930 667970 144950 668210
rect 145190 667970 145280 668210
rect 145520 667970 145610 668210
rect 145850 667970 145940 668210
rect 146180 667970 146290 668210
rect 146530 667970 146620 668210
rect 146860 667970 146950 668210
rect 147190 667970 147280 668210
rect 147520 667970 147630 668210
rect 147870 667970 147960 668210
rect 148200 667970 148290 668210
rect 148530 667970 148620 668210
rect 148860 667970 148970 668210
rect 149210 667970 149300 668210
rect 149540 667970 149630 668210
rect 149870 667970 149960 668210
rect 150200 667970 150310 668210
rect 150550 667970 150640 668210
rect 150880 667970 150970 668210
rect 151210 667970 151300 668210
rect 151540 667970 151650 668210
rect 151890 667970 151980 668210
rect 152220 667970 152310 668210
rect 152550 667970 152640 668210
rect 152880 667970 152990 668210
rect 153230 667970 153320 668210
rect 153560 667970 153650 668210
rect 153890 667970 153980 668210
rect 154220 667970 154330 668210
rect 154570 667970 154660 668210
rect 154900 667970 154990 668210
rect 155230 667970 155320 668210
rect 155560 667970 155670 668210
rect 155910 667970 155930 668210
rect 144930 667880 155930 667970
rect 144930 667640 144950 667880
rect 145190 667640 145280 667880
rect 145520 667640 145610 667880
rect 145850 667640 145940 667880
rect 146180 667640 146290 667880
rect 146530 667640 146620 667880
rect 146860 667640 146950 667880
rect 147190 667640 147280 667880
rect 147520 667640 147630 667880
rect 147870 667640 147960 667880
rect 148200 667640 148290 667880
rect 148530 667640 148620 667880
rect 148860 667640 148970 667880
rect 149210 667640 149300 667880
rect 149540 667640 149630 667880
rect 149870 667640 149960 667880
rect 150200 667640 150310 667880
rect 150550 667640 150640 667880
rect 150880 667640 150970 667880
rect 151210 667640 151300 667880
rect 151540 667640 151650 667880
rect 151890 667640 151980 667880
rect 152220 667640 152310 667880
rect 152550 667640 152640 667880
rect 152880 667640 152990 667880
rect 153230 667640 153320 667880
rect 153560 667640 153650 667880
rect 153890 667640 153980 667880
rect 154220 667640 154330 667880
rect 154570 667640 154660 667880
rect 154900 667640 154990 667880
rect 155230 667640 155320 667880
rect 155560 667640 155670 667880
rect 155910 667640 155930 667880
rect 144930 667530 155930 667640
rect 144930 667290 144950 667530
rect 145190 667290 145280 667530
rect 145520 667290 145610 667530
rect 145850 667290 145940 667530
rect 146180 667290 146290 667530
rect 146530 667290 146620 667530
rect 146860 667290 146950 667530
rect 147190 667290 147280 667530
rect 147520 667290 147630 667530
rect 147870 667290 147960 667530
rect 148200 667290 148290 667530
rect 148530 667290 148620 667530
rect 148860 667290 148970 667530
rect 149210 667290 149300 667530
rect 149540 667290 149630 667530
rect 149870 667290 149960 667530
rect 150200 667290 150310 667530
rect 150550 667290 150640 667530
rect 150880 667290 150970 667530
rect 151210 667290 151300 667530
rect 151540 667290 151650 667530
rect 151890 667290 151980 667530
rect 152220 667290 152310 667530
rect 152550 667290 152640 667530
rect 152880 667290 152990 667530
rect 153230 667290 153320 667530
rect 153560 667290 153650 667530
rect 153890 667290 153980 667530
rect 154220 667290 154330 667530
rect 154570 667290 154660 667530
rect 154900 667290 154990 667530
rect 155230 667290 155320 667530
rect 155560 667290 155670 667530
rect 155910 667290 155930 667530
rect 144930 667200 155930 667290
rect 144930 666960 144950 667200
rect 145190 666960 145280 667200
rect 145520 666960 145610 667200
rect 145850 666960 145940 667200
rect 146180 666960 146290 667200
rect 146530 666960 146620 667200
rect 146860 666960 146950 667200
rect 147190 666960 147280 667200
rect 147520 666960 147630 667200
rect 147870 666960 147960 667200
rect 148200 666960 148290 667200
rect 148530 666960 148620 667200
rect 148860 666960 148970 667200
rect 149210 666960 149300 667200
rect 149540 666960 149630 667200
rect 149870 666960 149960 667200
rect 150200 666960 150310 667200
rect 150550 666960 150640 667200
rect 150880 666960 150970 667200
rect 151210 666960 151300 667200
rect 151540 666960 151650 667200
rect 151890 666960 151980 667200
rect 152220 666960 152310 667200
rect 152550 666960 152640 667200
rect 152880 666960 152990 667200
rect 153230 666960 153320 667200
rect 153560 666960 153650 667200
rect 153890 666960 153980 667200
rect 154220 666960 154330 667200
rect 154570 666960 154660 667200
rect 154900 666960 154990 667200
rect 155230 666960 155320 667200
rect 155560 666960 155670 667200
rect 155910 666960 155930 667200
rect 144930 666870 155930 666960
rect 144930 666630 144950 666870
rect 145190 666630 145280 666870
rect 145520 666630 145610 666870
rect 145850 666630 145940 666870
rect 146180 666630 146290 666870
rect 146530 666630 146620 666870
rect 146860 666630 146950 666870
rect 147190 666630 147280 666870
rect 147520 666630 147630 666870
rect 147870 666630 147960 666870
rect 148200 666630 148290 666870
rect 148530 666630 148620 666870
rect 148860 666630 148970 666870
rect 149210 666630 149300 666870
rect 149540 666630 149630 666870
rect 149870 666630 149960 666870
rect 150200 666630 150310 666870
rect 150550 666630 150640 666870
rect 150880 666630 150970 666870
rect 151210 666630 151300 666870
rect 151540 666630 151650 666870
rect 151890 666630 151980 666870
rect 152220 666630 152310 666870
rect 152550 666630 152640 666870
rect 152880 666630 152990 666870
rect 153230 666630 153320 666870
rect 153560 666630 153650 666870
rect 153890 666630 153980 666870
rect 154220 666630 154330 666870
rect 154570 666630 154660 666870
rect 154900 666630 154990 666870
rect 155230 666630 155320 666870
rect 155560 666630 155670 666870
rect 155910 666630 155930 666870
rect 144930 666540 155930 666630
rect 144930 666300 144950 666540
rect 145190 666300 145280 666540
rect 145520 666300 145610 666540
rect 145850 666300 145940 666540
rect 146180 666300 146290 666540
rect 146530 666300 146620 666540
rect 146860 666300 146950 666540
rect 147190 666300 147280 666540
rect 147520 666300 147630 666540
rect 147870 666300 147960 666540
rect 148200 666300 148290 666540
rect 148530 666300 148620 666540
rect 148860 666300 148970 666540
rect 149210 666300 149300 666540
rect 149540 666300 149630 666540
rect 149870 666300 149960 666540
rect 150200 666300 150310 666540
rect 150550 666300 150640 666540
rect 150880 666300 150970 666540
rect 151210 666300 151300 666540
rect 151540 666300 151650 666540
rect 151890 666300 151980 666540
rect 152220 666300 152310 666540
rect 152550 666300 152640 666540
rect 152880 666300 152990 666540
rect 153230 666300 153320 666540
rect 153560 666300 153650 666540
rect 153890 666300 153980 666540
rect 154220 666300 154330 666540
rect 154570 666300 154660 666540
rect 154900 666300 154990 666540
rect 155230 666300 155320 666540
rect 155560 666300 155670 666540
rect 155910 666300 155930 666540
rect 144930 666190 155930 666300
rect 144930 665950 144950 666190
rect 145190 665950 145280 666190
rect 145520 665950 145610 666190
rect 145850 665950 145940 666190
rect 146180 665950 146290 666190
rect 146530 665950 146620 666190
rect 146860 665950 146950 666190
rect 147190 665950 147280 666190
rect 147520 665950 147630 666190
rect 147870 665950 147960 666190
rect 148200 665950 148290 666190
rect 148530 665950 148620 666190
rect 148860 665950 148970 666190
rect 149210 665950 149300 666190
rect 149540 665950 149630 666190
rect 149870 665950 149960 666190
rect 150200 665950 150310 666190
rect 150550 665950 150640 666190
rect 150880 665950 150970 666190
rect 151210 665950 151300 666190
rect 151540 665950 151650 666190
rect 151890 665950 151980 666190
rect 152220 665950 152310 666190
rect 152550 665950 152640 666190
rect 152880 665950 152990 666190
rect 153230 665950 153320 666190
rect 153560 665950 153650 666190
rect 153890 665950 153980 666190
rect 154220 665950 154330 666190
rect 154570 665950 154660 666190
rect 154900 665950 154990 666190
rect 155230 665950 155320 666190
rect 155560 665950 155670 666190
rect 155910 665950 155930 666190
rect 144930 665860 155930 665950
rect 144930 665620 144950 665860
rect 145190 665620 145280 665860
rect 145520 665620 145610 665860
rect 145850 665620 145940 665860
rect 146180 665620 146290 665860
rect 146530 665620 146620 665860
rect 146860 665620 146950 665860
rect 147190 665620 147280 665860
rect 147520 665620 147630 665860
rect 147870 665620 147960 665860
rect 148200 665620 148290 665860
rect 148530 665620 148620 665860
rect 148860 665620 148970 665860
rect 149210 665620 149300 665860
rect 149540 665620 149630 665860
rect 149870 665620 149960 665860
rect 150200 665620 150310 665860
rect 150550 665620 150640 665860
rect 150880 665620 150970 665860
rect 151210 665620 151300 665860
rect 151540 665620 151650 665860
rect 151890 665620 151980 665860
rect 152220 665620 152310 665860
rect 152550 665620 152640 665860
rect 152880 665620 152990 665860
rect 153230 665620 153320 665860
rect 153560 665620 153650 665860
rect 153890 665620 153980 665860
rect 154220 665620 154330 665860
rect 154570 665620 154660 665860
rect 154900 665620 154990 665860
rect 155230 665620 155320 665860
rect 155560 665620 155670 665860
rect 155910 665620 155930 665860
rect 144930 665530 155930 665620
rect 144930 665290 144950 665530
rect 145190 665290 145280 665530
rect 145520 665290 145610 665530
rect 145850 665290 145940 665530
rect 146180 665290 146290 665530
rect 146530 665290 146620 665530
rect 146860 665290 146950 665530
rect 147190 665290 147280 665530
rect 147520 665290 147630 665530
rect 147870 665290 147960 665530
rect 148200 665290 148290 665530
rect 148530 665290 148620 665530
rect 148860 665290 148970 665530
rect 149210 665290 149300 665530
rect 149540 665290 149630 665530
rect 149870 665290 149960 665530
rect 150200 665290 150310 665530
rect 150550 665290 150640 665530
rect 150880 665290 150970 665530
rect 151210 665290 151300 665530
rect 151540 665290 151650 665530
rect 151890 665290 151980 665530
rect 152220 665290 152310 665530
rect 152550 665290 152640 665530
rect 152880 665290 152990 665530
rect 153230 665290 153320 665530
rect 153560 665290 153650 665530
rect 153890 665290 153980 665530
rect 154220 665290 154330 665530
rect 154570 665290 154660 665530
rect 154900 665290 154990 665530
rect 155230 665290 155320 665530
rect 155560 665290 155670 665530
rect 155910 665290 155930 665530
rect 144930 665200 155930 665290
rect 144930 664960 144950 665200
rect 145190 664960 145280 665200
rect 145520 664960 145610 665200
rect 145850 664960 145940 665200
rect 146180 664960 146290 665200
rect 146530 664960 146620 665200
rect 146860 664960 146950 665200
rect 147190 664960 147280 665200
rect 147520 664960 147630 665200
rect 147870 664960 147960 665200
rect 148200 664960 148290 665200
rect 148530 664960 148620 665200
rect 148860 664960 148970 665200
rect 149210 664960 149300 665200
rect 149540 664960 149630 665200
rect 149870 664960 149960 665200
rect 150200 664960 150310 665200
rect 150550 664960 150640 665200
rect 150880 664960 150970 665200
rect 151210 664960 151300 665200
rect 151540 664960 151650 665200
rect 151890 664960 151980 665200
rect 152220 664960 152310 665200
rect 152550 664960 152640 665200
rect 152880 664960 152990 665200
rect 153230 664960 153320 665200
rect 153560 664960 153650 665200
rect 153890 664960 153980 665200
rect 154220 664960 154330 665200
rect 154570 664960 154660 665200
rect 154900 664960 154990 665200
rect 155230 664960 155320 665200
rect 155560 664960 155670 665200
rect 155910 664960 155930 665200
rect 144930 664850 155930 664960
rect 144930 664610 144950 664850
rect 145190 664610 145280 664850
rect 145520 664610 145610 664850
rect 145850 664610 145940 664850
rect 146180 664610 146290 664850
rect 146530 664610 146620 664850
rect 146860 664610 146950 664850
rect 147190 664610 147280 664850
rect 147520 664610 147630 664850
rect 147870 664610 147960 664850
rect 148200 664610 148290 664850
rect 148530 664610 148620 664850
rect 148860 664610 148970 664850
rect 149210 664610 149300 664850
rect 149540 664610 149630 664850
rect 149870 664610 149960 664850
rect 150200 664610 150310 664850
rect 150550 664610 150640 664850
rect 150880 664610 150970 664850
rect 151210 664610 151300 664850
rect 151540 664610 151650 664850
rect 151890 664610 151980 664850
rect 152220 664610 152310 664850
rect 152550 664610 152640 664850
rect 152880 664610 152990 664850
rect 153230 664610 153320 664850
rect 153560 664610 153650 664850
rect 153890 664610 153980 664850
rect 154220 664610 154330 664850
rect 154570 664610 154660 664850
rect 154900 664610 154990 664850
rect 155230 664610 155320 664850
rect 155560 664610 155670 664850
rect 155910 664610 155930 664850
rect 144930 664520 155930 664610
rect 144930 664280 144950 664520
rect 145190 664280 145280 664520
rect 145520 664280 145610 664520
rect 145850 664280 145940 664520
rect 146180 664280 146290 664520
rect 146530 664280 146620 664520
rect 146860 664280 146950 664520
rect 147190 664280 147280 664520
rect 147520 664280 147630 664520
rect 147870 664280 147960 664520
rect 148200 664280 148290 664520
rect 148530 664280 148620 664520
rect 148860 664280 148970 664520
rect 149210 664280 149300 664520
rect 149540 664280 149630 664520
rect 149870 664280 149960 664520
rect 150200 664280 150310 664520
rect 150550 664280 150640 664520
rect 150880 664280 150970 664520
rect 151210 664280 151300 664520
rect 151540 664280 151650 664520
rect 151890 664280 151980 664520
rect 152220 664280 152310 664520
rect 152550 664280 152640 664520
rect 152880 664280 152990 664520
rect 153230 664280 153320 664520
rect 153560 664280 153650 664520
rect 153890 664280 153980 664520
rect 154220 664280 154330 664520
rect 154570 664280 154660 664520
rect 154900 664280 154990 664520
rect 155230 664280 155320 664520
rect 155560 664280 155670 664520
rect 155910 664280 155930 664520
rect 144930 664190 155930 664280
rect 144930 663950 144950 664190
rect 145190 663950 145280 664190
rect 145520 663950 145610 664190
rect 145850 663950 145940 664190
rect 146180 663950 146290 664190
rect 146530 663950 146620 664190
rect 146860 663950 146950 664190
rect 147190 663950 147280 664190
rect 147520 663950 147630 664190
rect 147870 663950 147960 664190
rect 148200 663950 148290 664190
rect 148530 663950 148620 664190
rect 148860 663950 148970 664190
rect 149210 663950 149300 664190
rect 149540 663950 149630 664190
rect 149870 663950 149960 664190
rect 150200 663950 150310 664190
rect 150550 663950 150640 664190
rect 150880 663950 150970 664190
rect 151210 663950 151300 664190
rect 151540 663950 151650 664190
rect 151890 663950 151980 664190
rect 152220 663950 152310 664190
rect 152550 663950 152640 664190
rect 152880 663950 152990 664190
rect 153230 663950 153320 664190
rect 153560 663950 153650 664190
rect 153890 663950 153980 664190
rect 154220 663950 154330 664190
rect 154570 663950 154660 664190
rect 154900 663950 154990 664190
rect 155230 663950 155320 664190
rect 155560 663950 155670 664190
rect 155910 663950 155930 664190
rect 144930 663860 155930 663950
rect 144930 663620 144950 663860
rect 145190 663620 145280 663860
rect 145520 663620 145610 663860
rect 145850 663620 145940 663860
rect 146180 663620 146290 663860
rect 146530 663620 146620 663860
rect 146860 663620 146950 663860
rect 147190 663620 147280 663860
rect 147520 663620 147630 663860
rect 147870 663620 147960 663860
rect 148200 663620 148290 663860
rect 148530 663620 148620 663860
rect 148860 663620 148970 663860
rect 149210 663620 149300 663860
rect 149540 663620 149630 663860
rect 149870 663620 149960 663860
rect 150200 663620 150310 663860
rect 150550 663620 150640 663860
rect 150880 663620 150970 663860
rect 151210 663620 151300 663860
rect 151540 663620 151650 663860
rect 151890 663620 151980 663860
rect 152220 663620 152310 663860
rect 152550 663620 152640 663860
rect 152880 663620 152990 663860
rect 153230 663620 153320 663860
rect 153560 663620 153650 663860
rect 153890 663620 153980 663860
rect 154220 663620 154330 663860
rect 154570 663620 154660 663860
rect 154900 663620 154990 663860
rect 155230 663620 155320 663860
rect 155560 663620 155670 663860
rect 155910 663620 155930 663860
rect 144930 663510 155930 663620
rect 144930 663270 144950 663510
rect 145190 663270 145280 663510
rect 145520 663270 145610 663510
rect 145850 663270 145940 663510
rect 146180 663270 146290 663510
rect 146530 663270 146620 663510
rect 146860 663270 146950 663510
rect 147190 663270 147280 663510
rect 147520 663270 147630 663510
rect 147870 663270 147960 663510
rect 148200 663270 148290 663510
rect 148530 663270 148620 663510
rect 148860 663270 148970 663510
rect 149210 663270 149300 663510
rect 149540 663270 149630 663510
rect 149870 663270 149960 663510
rect 150200 663270 150310 663510
rect 150550 663270 150640 663510
rect 150880 663270 150970 663510
rect 151210 663270 151300 663510
rect 151540 663270 151650 663510
rect 151890 663270 151980 663510
rect 152220 663270 152310 663510
rect 152550 663270 152640 663510
rect 152880 663270 152990 663510
rect 153230 663270 153320 663510
rect 153560 663270 153650 663510
rect 153890 663270 153980 663510
rect 154220 663270 154330 663510
rect 154570 663270 154660 663510
rect 154900 663270 154990 663510
rect 155230 663270 155320 663510
rect 155560 663270 155670 663510
rect 155910 663270 155930 663510
rect 144930 663180 155930 663270
rect 144930 662940 144950 663180
rect 145190 662940 145280 663180
rect 145520 662940 145610 663180
rect 145850 662940 145940 663180
rect 146180 662940 146290 663180
rect 146530 662940 146620 663180
rect 146860 662940 146950 663180
rect 147190 662940 147280 663180
rect 147520 662940 147630 663180
rect 147870 662940 147960 663180
rect 148200 662940 148290 663180
rect 148530 662940 148620 663180
rect 148860 662940 148970 663180
rect 149210 662940 149300 663180
rect 149540 662940 149630 663180
rect 149870 662940 149960 663180
rect 150200 662940 150310 663180
rect 150550 662940 150640 663180
rect 150880 662940 150970 663180
rect 151210 662940 151300 663180
rect 151540 662940 151650 663180
rect 151890 662940 151980 663180
rect 152220 662940 152310 663180
rect 152550 662940 152640 663180
rect 152880 662940 152990 663180
rect 153230 662940 153320 663180
rect 153560 662940 153650 663180
rect 153890 662940 153980 663180
rect 154220 662940 154330 663180
rect 154570 662940 154660 663180
rect 154900 662940 154990 663180
rect 155230 662940 155320 663180
rect 155560 662940 155670 663180
rect 155910 662940 155930 663180
rect 144930 662850 155930 662940
rect 144930 662610 144950 662850
rect 145190 662610 145280 662850
rect 145520 662610 145610 662850
rect 145850 662610 145940 662850
rect 146180 662610 146290 662850
rect 146530 662610 146620 662850
rect 146860 662610 146950 662850
rect 147190 662610 147280 662850
rect 147520 662610 147630 662850
rect 147870 662610 147960 662850
rect 148200 662610 148290 662850
rect 148530 662610 148620 662850
rect 148860 662610 148970 662850
rect 149210 662610 149300 662850
rect 149540 662610 149630 662850
rect 149870 662610 149960 662850
rect 150200 662610 150310 662850
rect 150550 662610 150640 662850
rect 150880 662610 150970 662850
rect 151210 662610 151300 662850
rect 151540 662610 151650 662850
rect 151890 662610 151980 662850
rect 152220 662610 152310 662850
rect 152550 662610 152640 662850
rect 152880 662610 152990 662850
rect 153230 662610 153320 662850
rect 153560 662610 153650 662850
rect 153890 662610 153980 662850
rect 154220 662610 154330 662850
rect 154570 662610 154660 662850
rect 154900 662610 154990 662850
rect 155230 662610 155320 662850
rect 155560 662610 155670 662850
rect 155910 662610 155930 662850
rect 144930 662520 155930 662610
rect 144930 662280 144950 662520
rect 145190 662280 145280 662520
rect 145520 662280 145610 662520
rect 145850 662280 145940 662520
rect 146180 662280 146290 662520
rect 146530 662280 146620 662520
rect 146860 662280 146950 662520
rect 147190 662280 147280 662520
rect 147520 662280 147630 662520
rect 147870 662280 147960 662520
rect 148200 662280 148290 662520
rect 148530 662280 148620 662520
rect 148860 662280 148970 662520
rect 149210 662280 149300 662520
rect 149540 662280 149630 662520
rect 149870 662280 149960 662520
rect 150200 662280 150310 662520
rect 150550 662280 150640 662520
rect 150880 662280 150970 662520
rect 151210 662280 151300 662520
rect 151540 662280 151650 662520
rect 151890 662280 151980 662520
rect 152220 662280 152310 662520
rect 152550 662280 152640 662520
rect 152880 662280 152990 662520
rect 153230 662280 153320 662520
rect 153560 662280 153650 662520
rect 153890 662280 153980 662520
rect 154220 662280 154330 662520
rect 154570 662280 154660 662520
rect 154900 662280 154990 662520
rect 155230 662280 155320 662520
rect 155560 662280 155670 662520
rect 155910 662280 155930 662520
rect 144930 662170 155930 662280
rect 144930 661930 144950 662170
rect 145190 661930 145280 662170
rect 145520 661930 145610 662170
rect 145850 661930 145940 662170
rect 146180 661930 146290 662170
rect 146530 661930 146620 662170
rect 146860 661930 146950 662170
rect 147190 661930 147280 662170
rect 147520 661930 147630 662170
rect 147870 661930 147960 662170
rect 148200 661930 148290 662170
rect 148530 661930 148620 662170
rect 148860 661930 148970 662170
rect 149210 661930 149300 662170
rect 149540 661930 149630 662170
rect 149870 661930 149960 662170
rect 150200 661930 150310 662170
rect 150550 661930 150640 662170
rect 150880 661930 150970 662170
rect 151210 661930 151300 662170
rect 151540 661930 151650 662170
rect 151890 661930 151980 662170
rect 152220 661930 152310 662170
rect 152550 661930 152640 662170
rect 152880 661930 152990 662170
rect 153230 661930 153320 662170
rect 153560 661930 153650 662170
rect 153890 661930 153980 662170
rect 154220 661930 154330 662170
rect 154570 661930 154660 662170
rect 154900 661930 154990 662170
rect 155230 661930 155320 662170
rect 155560 661930 155670 662170
rect 155910 661930 155930 662170
rect 144930 661840 155930 661930
rect 144930 661600 144950 661840
rect 145190 661600 145280 661840
rect 145520 661600 145610 661840
rect 145850 661600 145940 661840
rect 146180 661600 146290 661840
rect 146530 661600 146620 661840
rect 146860 661600 146950 661840
rect 147190 661600 147280 661840
rect 147520 661600 147630 661840
rect 147870 661600 147960 661840
rect 148200 661600 148290 661840
rect 148530 661600 148620 661840
rect 148860 661600 148970 661840
rect 149210 661600 149300 661840
rect 149540 661600 149630 661840
rect 149870 661600 149960 661840
rect 150200 661600 150310 661840
rect 150550 661600 150640 661840
rect 150880 661600 150970 661840
rect 151210 661600 151300 661840
rect 151540 661600 151650 661840
rect 151890 661600 151980 661840
rect 152220 661600 152310 661840
rect 152550 661600 152640 661840
rect 152880 661600 152990 661840
rect 153230 661600 153320 661840
rect 153560 661600 153650 661840
rect 153890 661600 153980 661840
rect 154220 661600 154330 661840
rect 154570 661600 154660 661840
rect 154900 661600 154990 661840
rect 155230 661600 155320 661840
rect 155560 661600 155670 661840
rect 155910 661600 155930 661840
rect 144930 661510 155930 661600
rect 144930 661270 144950 661510
rect 145190 661270 145280 661510
rect 145520 661270 145610 661510
rect 145850 661270 145940 661510
rect 146180 661270 146290 661510
rect 146530 661270 146620 661510
rect 146860 661270 146950 661510
rect 147190 661270 147280 661510
rect 147520 661270 147630 661510
rect 147870 661270 147960 661510
rect 148200 661270 148290 661510
rect 148530 661270 148620 661510
rect 148860 661270 148970 661510
rect 149210 661270 149300 661510
rect 149540 661270 149630 661510
rect 149870 661270 149960 661510
rect 150200 661270 150310 661510
rect 150550 661270 150640 661510
rect 150880 661270 150970 661510
rect 151210 661270 151300 661510
rect 151540 661270 151650 661510
rect 151890 661270 151980 661510
rect 152220 661270 152310 661510
rect 152550 661270 152640 661510
rect 152880 661270 152990 661510
rect 153230 661270 153320 661510
rect 153560 661270 153650 661510
rect 153890 661270 153980 661510
rect 154220 661270 154330 661510
rect 154570 661270 154660 661510
rect 154900 661270 154990 661510
rect 155230 661270 155320 661510
rect 155560 661270 155670 661510
rect 155910 661270 155930 661510
rect 144930 661180 155930 661270
rect 144930 660940 144950 661180
rect 145190 660940 145280 661180
rect 145520 660940 145610 661180
rect 145850 660940 145940 661180
rect 146180 660940 146290 661180
rect 146530 660940 146620 661180
rect 146860 660940 146950 661180
rect 147190 660940 147280 661180
rect 147520 660940 147630 661180
rect 147870 660940 147960 661180
rect 148200 660940 148290 661180
rect 148530 660940 148620 661180
rect 148860 660940 148970 661180
rect 149210 660940 149300 661180
rect 149540 660940 149630 661180
rect 149870 660940 149960 661180
rect 150200 660940 150310 661180
rect 150550 660940 150640 661180
rect 150880 660940 150970 661180
rect 151210 660940 151300 661180
rect 151540 660940 151650 661180
rect 151890 660940 151980 661180
rect 152220 660940 152310 661180
rect 152550 660940 152640 661180
rect 152880 660940 152990 661180
rect 153230 660940 153320 661180
rect 153560 660940 153650 661180
rect 153890 660940 153980 661180
rect 154220 660940 154330 661180
rect 154570 660940 154660 661180
rect 154900 660940 154990 661180
rect 155230 660940 155320 661180
rect 155560 660940 155670 661180
rect 155910 660940 155930 661180
rect 144930 660920 155930 660940
rect 110790 660340 121790 660360
rect 110790 660100 110810 660340
rect 111050 660100 111160 660340
rect 111400 660100 111490 660340
rect 111730 660100 111820 660340
rect 112060 660100 112150 660340
rect 112390 660100 112500 660340
rect 112740 660100 112830 660340
rect 113070 660100 113160 660340
rect 113400 660100 113490 660340
rect 113730 660100 113840 660340
rect 114080 660100 114170 660340
rect 114410 660100 114500 660340
rect 114740 660100 114830 660340
rect 115070 660100 115180 660340
rect 115420 660100 115510 660340
rect 115750 660100 115840 660340
rect 116080 660100 116170 660340
rect 116410 660100 116520 660340
rect 116760 660100 116850 660340
rect 117090 660100 117180 660340
rect 117420 660100 117510 660340
rect 117750 660100 117860 660340
rect 118100 660100 118190 660340
rect 118430 660100 118520 660340
rect 118760 660100 118850 660340
rect 119090 660100 119200 660340
rect 119440 660100 119530 660340
rect 119770 660100 119860 660340
rect 120100 660100 120190 660340
rect 120430 660100 120540 660340
rect 120780 660100 120870 660340
rect 121110 660100 121200 660340
rect 121440 660100 121530 660340
rect 121770 660100 121790 660340
rect 110790 660010 121790 660100
rect 110790 659770 110810 660010
rect 111050 659770 111160 660010
rect 111400 659770 111490 660010
rect 111730 659770 111820 660010
rect 112060 659770 112150 660010
rect 112390 659770 112500 660010
rect 112740 659770 112830 660010
rect 113070 659770 113160 660010
rect 113400 659770 113490 660010
rect 113730 659770 113840 660010
rect 114080 659770 114170 660010
rect 114410 659770 114500 660010
rect 114740 659770 114830 660010
rect 115070 659770 115180 660010
rect 115420 659770 115510 660010
rect 115750 659770 115840 660010
rect 116080 659770 116170 660010
rect 116410 659770 116520 660010
rect 116760 659770 116850 660010
rect 117090 659770 117180 660010
rect 117420 659770 117510 660010
rect 117750 659770 117860 660010
rect 118100 659770 118190 660010
rect 118430 659770 118520 660010
rect 118760 659770 118850 660010
rect 119090 659770 119200 660010
rect 119440 659770 119530 660010
rect 119770 659770 119860 660010
rect 120100 659770 120190 660010
rect 120430 659770 120540 660010
rect 120780 659770 120870 660010
rect 121110 659770 121200 660010
rect 121440 659770 121530 660010
rect 121770 659770 121790 660010
rect 110790 659680 121790 659770
rect 110790 659440 110810 659680
rect 111050 659440 111160 659680
rect 111400 659440 111490 659680
rect 111730 659440 111820 659680
rect 112060 659440 112150 659680
rect 112390 659440 112500 659680
rect 112740 659440 112830 659680
rect 113070 659440 113160 659680
rect 113400 659440 113490 659680
rect 113730 659440 113840 659680
rect 114080 659440 114170 659680
rect 114410 659440 114500 659680
rect 114740 659440 114830 659680
rect 115070 659440 115180 659680
rect 115420 659440 115510 659680
rect 115750 659440 115840 659680
rect 116080 659440 116170 659680
rect 116410 659440 116520 659680
rect 116760 659440 116850 659680
rect 117090 659440 117180 659680
rect 117420 659440 117510 659680
rect 117750 659440 117860 659680
rect 118100 659440 118190 659680
rect 118430 659440 118520 659680
rect 118760 659440 118850 659680
rect 119090 659440 119200 659680
rect 119440 659440 119530 659680
rect 119770 659440 119860 659680
rect 120100 659440 120190 659680
rect 120430 659440 120540 659680
rect 120780 659440 120870 659680
rect 121110 659440 121200 659680
rect 121440 659440 121530 659680
rect 121770 659440 121790 659680
rect 110790 659350 121790 659440
rect 110790 659110 110810 659350
rect 111050 659110 111160 659350
rect 111400 659110 111490 659350
rect 111730 659110 111820 659350
rect 112060 659110 112150 659350
rect 112390 659110 112500 659350
rect 112740 659110 112830 659350
rect 113070 659110 113160 659350
rect 113400 659110 113490 659350
rect 113730 659110 113840 659350
rect 114080 659110 114170 659350
rect 114410 659110 114500 659350
rect 114740 659110 114830 659350
rect 115070 659110 115180 659350
rect 115420 659110 115510 659350
rect 115750 659110 115840 659350
rect 116080 659110 116170 659350
rect 116410 659110 116520 659350
rect 116760 659110 116850 659350
rect 117090 659110 117180 659350
rect 117420 659110 117510 659350
rect 117750 659110 117860 659350
rect 118100 659110 118190 659350
rect 118430 659110 118520 659350
rect 118760 659110 118850 659350
rect 119090 659110 119200 659350
rect 119440 659110 119530 659350
rect 119770 659110 119860 659350
rect 120100 659110 120190 659350
rect 120430 659110 120540 659350
rect 120780 659110 120870 659350
rect 121110 659110 121200 659350
rect 121440 659110 121530 659350
rect 121770 659110 121790 659350
rect 110790 659000 121790 659110
rect 110790 658760 110810 659000
rect 111050 658760 111160 659000
rect 111400 658760 111490 659000
rect 111730 658760 111820 659000
rect 112060 658760 112150 659000
rect 112390 658760 112500 659000
rect 112740 658760 112830 659000
rect 113070 658760 113160 659000
rect 113400 658760 113490 659000
rect 113730 658760 113840 659000
rect 114080 658760 114170 659000
rect 114410 658760 114500 659000
rect 114740 658760 114830 659000
rect 115070 658760 115180 659000
rect 115420 658760 115510 659000
rect 115750 658760 115840 659000
rect 116080 658760 116170 659000
rect 116410 658760 116520 659000
rect 116760 658760 116850 659000
rect 117090 658760 117180 659000
rect 117420 658760 117510 659000
rect 117750 658760 117860 659000
rect 118100 658760 118190 659000
rect 118430 658760 118520 659000
rect 118760 658760 118850 659000
rect 119090 658760 119200 659000
rect 119440 658760 119530 659000
rect 119770 658760 119860 659000
rect 120100 658760 120190 659000
rect 120430 658760 120540 659000
rect 120780 658760 120870 659000
rect 121110 658760 121200 659000
rect 121440 658760 121530 659000
rect 121770 658760 121790 659000
rect 110790 658670 121790 658760
rect 110790 658430 110810 658670
rect 111050 658430 111160 658670
rect 111400 658430 111490 658670
rect 111730 658430 111820 658670
rect 112060 658430 112150 658670
rect 112390 658430 112500 658670
rect 112740 658430 112830 658670
rect 113070 658430 113160 658670
rect 113400 658430 113490 658670
rect 113730 658430 113840 658670
rect 114080 658430 114170 658670
rect 114410 658430 114500 658670
rect 114740 658430 114830 658670
rect 115070 658430 115180 658670
rect 115420 658430 115510 658670
rect 115750 658430 115840 658670
rect 116080 658430 116170 658670
rect 116410 658430 116520 658670
rect 116760 658430 116850 658670
rect 117090 658430 117180 658670
rect 117420 658430 117510 658670
rect 117750 658430 117860 658670
rect 118100 658430 118190 658670
rect 118430 658430 118520 658670
rect 118760 658430 118850 658670
rect 119090 658430 119200 658670
rect 119440 658430 119530 658670
rect 119770 658430 119860 658670
rect 120100 658430 120190 658670
rect 120430 658430 120540 658670
rect 120780 658430 120870 658670
rect 121110 658430 121200 658670
rect 121440 658430 121530 658670
rect 121770 658430 121790 658670
rect 110790 658340 121790 658430
rect 110790 658100 110810 658340
rect 111050 658100 111160 658340
rect 111400 658100 111490 658340
rect 111730 658100 111820 658340
rect 112060 658100 112150 658340
rect 112390 658100 112500 658340
rect 112740 658100 112830 658340
rect 113070 658100 113160 658340
rect 113400 658100 113490 658340
rect 113730 658100 113840 658340
rect 114080 658100 114170 658340
rect 114410 658100 114500 658340
rect 114740 658100 114830 658340
rect 115070 658100 115180 658340
rect 115420 658100 115510 658340
rect 115750 658100 115840 658340
rect 116080 658100 116170 658340
rect 116410 658100 116520 658340
rect 116760 658100 116850 658340
rect 117090 658100 117180 658340
rect 117420 658100 117510 658340
rect 117750 658100 117860 658340
rect 118100 658100 118190 658340
rect 118430 658100 118520 658340
rect 118760 658100 118850 658340
rect 119090 658100 119200 658340
rect 119440 658100 119530 658340
rect 119770 658100 119860 658340
rect 120100 658100 120190 658340
rect 120430 658100 120540 658340
rect 120780 658100 120870 658340
rect 121110 658100 121200 658340
rect 121440 658100 121530 658340
rect 121770 658100 121790 658340
rect 110790 658010 121790 658100
rect 110790 657770 110810 658010
rect 111050 657770 111160 658010
rect 111400 657770 111490 658010
rect 111730 657770 111820 658010
rect 112060 657770 112150 658010
rect 112390 657770 112500 658010
rect 112740 657770 112830 658010
rect 113070 657770 113160 658010
rect 113400 657770 113490 658010
rect 113730 657770 113840 658010
rect 114080 657770 114170 658010
rect 114410 657770 114500 658010
rect 114740 657770 114830 658010
rect 115070 657770 115180 658010
rect 115420 657770 115510 658010
rect 115750 657770 115840 658010
rect 116080 657770 116170 658010
rect 116410 657770 116520 658010
rect 116760 657770 116850 658010
rect 117090 657770 117180 658010
rect 117420 657770 117510 658010
rect 117750 657770 117860 658010
rect 118100 657770 118190 658010
rect 118430 657770 118520 658010
rect 118760 657770 118850 658010
rect 119090 657770 119200 658010
rect 119440 657770 119530 658010
rect 119770 657770 119860 658010
rect 120100 657770 120190 658010
rect 120430 657770 120540 658010
rect 120780 657770 120870 658010
rect 121110 657770 121200 658010
rect 121440 657770 121530 658010
rect 121770 657770 121790 658010
rect 110790 657660 121790 657770
rect 110790 657420 110810 657660
rect 111050 657420 111160 657660
rect 111400 657420 111490 657660
rect 111730 657420 111820 657660
rect 112060 657420 112150 657660
rect 112390 657420 112500 657660
rect 112740 657420 112830 657660
rect 113070 657420 113160 657660
rect 113400 657420 113490 657660
rect 113730 657420 113840 657660
rect 114080 657420 114170 657660
rect 114410 657420 114500 657660
rect 114740 657420 114830 657660
rect 115070 657420 115180 657660
rect 115420 657420 115510 657660
rect 115750 657420 115840 657660
rect 116080 657420 116170 657660
rect 116410 657420 116520 657660
rect 116760 657420 116850 657660
rect 117090 657420 117180 657660
rect 117420 657420 117510 657660
rect 117750 657420 117860 657660
rect 118100 657420 118190 657660
rect 118430 657420 118520 657660
rect 118760 657420 118850 657660
rect 119090 657420 119200 657660
rect 119440 657420 119530 657660
rect 119770 657420 119860 657660
rect 120100 657420 120190 657660
rect 120430 657420 120540 657660
rect 120780 657420 120870 657660
rect 121110 657420 121200 657660
rect 121440 657420 121530 657660
rect 121770 657420 121790 657660
rect 110790 657330 121790 657420
rect 110790 657090 110810 657330
rect 111050 657090 111160 657330
rect 111400 657090 111490 657330
rect 111730 657090 111820 657330
rect 112060 657090 112150 657330
rect 112390 657090 112500 657330
rect 112740 657090 112830 657330
rect 113070 657090 113160 657330
rect 113400 657090 113490 657330
rect 113730 657090 113840 657330
rect 114080 657090 114170 657330
rect 114410 657090 114500 657330
rect 114740 657090 114830 657330
rect 115070 657090 115180 657330
rect 115420 657090 115510 657330
rect 115750 657090 115840 657330
rect 116080 657090 116170 657330
rect 116410 657090 116520 657330
rect 116760 657090 116850 657330
rect 117090 657090 117180 657330
rect 117420 657090 117510 657330
rect 117750 657090 117860 657330
rect 118100 657090 118190 657330
rect 118430 657090 118520 657330
rect 118760 657090 118850 657330
rect 119090 657090 119200 657330
rect 119440 657090 119530 657330
rect 119770 657090 119860 657330
rect 120100 657090 120190 657330
rect 120430 657090 120540 657330
rect 120780 657090 120870 657330
rect 121110 657090 121200 657330
rect 121440 657090 121530 657330
rect 121770 657090 121790 657330
rect 110790 657000 121790 657090
rect 110790 656760 110810 657000
rect 111050 656760 111160 657000
rect 111400 656760 111490 657000
rect 111730 656760 111820 657000
rect 112060 656760 112150 657000
rect 112390 656760 112500 657000
rect 112740 656760 112830 657000
rect 113070 656760 113160 657000
rect 113400 656760 113490 657000
rect 113730 656760 113840 657000
rect 114080 656760 114170 657000
rect 114410 656760 114500 657000
rect 114740 656760 114830 657000
rect 115070 656760 115180 657000
rect 115420 656760 115510 657000
rect 115750 656760 115840 657000
rect 116080 656760 116170 657000
rect 116410 656760 116520 657000
rect 116760 656760 116850 657000
rect 117090 656760 117180 657000
rect 117420 656760 117510 657000
rect 117750 656760 117860 657000
rect 118100 656760 118190 657000
rect 118430 656760 118520 657000
rect 118760 656760 118850 657000
rect 119090 656760 119200 657000
rect 119440 656760 119530 657000
rect 119770 656760 119860 657000
rect 120100 656760 120190 657000
rect 120430 656760 120540 657000
rect 120780 656760 120870 657000
rect 121110 656760 121200 657000
rect 121440 656760 121530 657000
rect 121770 656760 121790 657000
rect 110790 656670 121790 656760
rect 110790 656430 110810 656670
rect 111050 656430 111160 656670
rect 111400 656430 111490 656670
rect 111730 656430 111820 656670
rect 112060 656430 112150 656670
rect 112390 656430 112500 656670
rect 112740 656430 112830 656670
rect 113070 656430 113160 656670
rect 113400 656430 113490 656670
rect 113730 656430 113840 656670
rect 114080 656430 114170 656670
rect 114410 656430 114500 656670
rect 114740 656430 114830 656670
rect 115070 656430 115180 656670
rect 115420 656430 115510 656670
rect 115750 656430 115840 656670
rect 116080 656430 116170 656670
rect 116410 656430 116520 656670
rect 116760 656430 116850 656670
rect 117090 656430 117180 656670
rect 117420 656430 117510 656670
rect 117750 656430 117860 656670
rect 118100 656430 118190 656670
rect 118430 656430 118520 656670
rect 118760 656430 118850 656670
rect 119090 656430 119200 656670
rect 119440 656430 119530 656670
rect 119770 656430 119860 656670
rect 120100 656430 120190 656670
rect 120430 656430 120540 656670
rect 120780 656430 120870 656670
rect 121110 656430 121200 656670
rect 121440 656430 121530 656670
rect 121770 656430 121790 656670
rect 110790 656320 121790 656430
rect 110790 656080 110810 656320
rect 111050 656080 111160 656320
rect 111400 656080 111490 656320
rect 111730 656080 111820 656320
rect 112060 656080 112150 656320
rect 112390 656080 112500 656320
rect 112740 656080 112830 656320
rect 113070 656080 113160 656320
rect 113400 656080 113490 656320
rect 113730 656080 113840 656320
rect 114080 656080 114170 656320
rect 114410 656080 114500 656320
rect 114740 656080 114830 656320
rect 115070 656080 115180 656320
rect 115420 656080 115510 656320
rect 115750 656080 115840 656320
rect 116080 656080 116170 656320
rect 116410 656080 116520 656320
rect 116760 656080 116850 656320
rect 117090 656080 117180 656320
rect 117420 656080 117510 656320
rect 117750 656080 117860 656320
rect 118100 656080 118190 656320
rect 118430 656080 118520 656320
rect 118760 656080 118850 656320
rect 119090 656080 119200 656320
rect 119440 656080 119530 656320
rect 119770 656080 119860 656320
rect 120100 656080 120190 656320
rect 120430 656080 120540 656320
rect 120780 656080 120870 656320
rect 121110 656080 121200 656320
rect 121440 656080 121530 656320
rect 121770 656080 121790 656320
rect 110790 655990 121790 656080
rect 110790 655750 110810 655990
rect 111050 655750 111160 655990
rect 111400 655750 111490 655990
rect 111730 655750 111820 655990
rect 112060 655750 112150 655990
rect 112390 655750 112500 655990
rect 112740 655750 112830 655990
rect 113070 655750 113160 655990
rect 113400 655750 113490 655990
rect 113730 655750 113840 655990
rect 114080 655750 114170 655990
rect 114410 655750 114500 655990
rect 114740 655750 114830 655990
rect 115070 655750 115180 655990
rect 115420 655750 115510 655990
rect 115750 655750 115840 655990
rect 116080 655750 116170 655990
rect 116410 655750 116520 655990
rect 116760 655750 116850 655990
rect 117090 655750 117180 655990
rect 117420 655750 117510 655990
rect 117750 655750 117860 655990
rect 118100 655750 118190 655990
rect 118430 655750 118520 655990
rect 118760 655750 118850 655990
rect 119090 655750 119200 655990
rect 119440 655750 119530 655990
rect 119770 655750 119860 655990
rect 120100 655750 120190 655990
rect 120430 655750 120540 655990
rect 120780 655750 120870 655990
rect 121110 655750 121200 655990
rect 121440 655750 121530 655990
rect 121770 655750 121790 655990
rect 110790 655660 121790 655750
rect 110790 655420 110810 655660
rect 111050 655420 111160 655660
rect 111400 655420 111490 655660
rect 111730 655420 111820 655660
rect 112060 655420 112150 655660
rect 112390 655420 112500 655660
rect 112740 655420 112830 655660
rect 113070 655420 113160 655660
rect 113400 655420 113490 655660
rect 113730 655420 113840 655660
rect 114080 655420 114170 655660
rect 114410 655420 114500 655660
rect 114740 655420 114830 655660
rect 115070 655420 115180 655660
rect 115420 655420 115510 655660
rect 115750 655420 115840 655660
rect 116080 655420 116170 655660
rect 116410 655420 116520 655660
rect 116760 655420 116850 655660
rect 117090 655420 117180 655660
rect 117420 655420 117510 655660
rect 117750 655420 117860 655660
rect 118100 655420 118190 655660
rect 118430 655420 118520 655660
rect 118760 655420 118850 655660
rect 119090 655420 119200 655660
rect 119440 655420 119530 655660
rect 119770 655420 119860 655660
rect 120100 655420 120190 655660
rect 120430 655420 120540 655660
rect 120780 655420 120870 655660
rect 121110 655420 121200 655660
rect 121440 655420 121530 655660
rect 121770 655420 121790 655660
rect 110790 655330 121790 655420
rect 110790 655090 110810 655330
rect 111050 655090 111160 655330
rect 111400 655090 111490 655330
rect 111730 655090 111820 655330
rect 112060 655090 112150 655330
rect 112390 655090 112500 655330
rect 112740 655090 112830 655330
rect 113070 655090 113160 655330
rect 113400 655090 113490 655330
rect 113730 655090 113840 655330
rect 114080 655090 114170 655330
rect 114410 655090 114500 655330
rect 114740 655090 114830 655330
rect 115070 655090 115180 655330
rect 115420 655090 115510 655330
rect 115750 655090 115840 655330
rect 116080 655090 116170 655330
rect 116410 655090 116520 655330
rect 116760 655090 116850 655330
rect 117090 655090 117180 655330
rect 117420 655090 117510 655330
rect 117750 655090 117860 655330
rect 118100 655090 118190 655330
rect 118430 655090 118520 655330
rect 118760 655090 118850 655330
rect 119090 655090 119200 655330
rect 119440 655090 119530 655330
rect 119770 655090 119860 655330
rect 120100 655090 120190 655330
rect 120430 655090 120540 655330
rect 120780 655090 120870 655330
rect 121110 655090 121200 655330
rect 121440 655090 121530 655330
rect 121770 655090 121790 655330
rect 110790 654980 121790 655090
rect 110790 654740 110810 654980
rect 111050 654740 111160 654980
rect 111400 654740 111490 654980
rect 111730 654740 111820 654980
rect 112060 654740 112150 654980
rect 112390 654740 112500 654980
rect 112740 654740 112830 654980
rect 113070 654740 113160 654980
rect 113400 654740 113490 654980
rect 113730 654740 113840 654980
rect 114080 654740 114170 654980
rect 114410 654740 114500 654980
rect 114740 654740 114830 654980
rect 115070 654740 115180 654980
rect 115420 654740 115510 654980
rect 115750 654740 115840 654980
rect 116080 654740 116170 654980
rect 116410 654740 116520 654980
rect 116760 654740 116850 654980
rect 117090 654740 117180 654980
rect 117420 654740 117510 654980
rect 117750 654740 117860 654980
rect 118100 654740 118190 654980
rect 118430 654740 118520 654980
rect 118760 654740 118850 654980
rect 119090 654740 119200 654980
rect 119440 654740 119530 654980
rect 119770 654740 119860 654980
rect 120100 654740 120190 654980
rect 120430 654740 120540 654980
rect 120780 654740 120870 654980
rect 121110 654740 121200 654980
rect 121440 654740 121530 654980
rect 121770 654740 121790 654980
rect 110790 654650 121790 654740
rect 110790 654410 110810 654650
rect 111050 654410 111160 654650
rect 111400 654410 111490 654650
rect 111730 654410 111820 654650
rect 112060 654410 112150 654650
rect 112390 654410 112500 654650
rect 112740 654410 112830 654650
rect 113070 654410 113160 654650
rect 113400 654410 113490 654650
rect 113730 654410 113840 654650
rect 114080 654410 114170 654650
rect 114410 654410 114500 654650
rect 114740 654410 114830 654650
rect 115070 654410 115180 654650
rect 115420 654410 115510 654650
rect 115750 654410 115840 654650
rect 116080 654410 116170 654650
rect 116410 654410 116520 654650
rect 116760 654410 116850 654650
rect 117090 654410 117180 654650
rect 117420 654410 117510 654650
rect 117750 654410 117860 654650
rect 118100 654410 118190 654650
rect 118430 654410 118520 654650
rect 118760 654410 118850 654650
rect 119090 654410 119200 654650
rect 119440 654410 119530 654650
rect 119770 654410 119860 654650
rect 120100 654410 120190 654650
rect 120430 654410 120540 654650
rect 120780 654410 120870 654650
rect 121110 654410 121200 654650
rect 121440 654410 121530 654650
rect 121770 654410 121790 654650
rect 110790 654320 121790 654410
rect 110790 654080 110810 654320
rect 111050 654080 111160 654320
rect 111400 654080 111490 654320
rect 111730 654080 111820 654320
rect 112060 654080 112150 654320
rect 112390 654080 112500 654320
rect 112740 654080 112830 654320
rect 113070 654080 113160 654320
rect 113400 654080 113490 654320
rect 113730 654080 113840 654320
rect 114080 654080 114170 654320
rect 114410 654080 114500 654320
rect 114740 654080 114830 654320
rect 115070 654080 115180 654320
rect 115420 654080 115510 654320
rect 115750 654080 115840 654320
rect 116080 654080 116170 654320
rect 116410 654080 116520 654320
rect 116760 654080 116850 654320
rect 117090 654080 117180 654320
rect 117420 654080 117510 654320
rect 117750 654080 117860 654320
rect 118100 654080 118190 654320
rect 118430 654080 118520 654320
rect 118760 654080 118850 654320
rect 119090 654080 119200 654320
rect 119440 654080 119530 654320
rect 119770 654080 119860 654320
rect 120100 654080 120190 654320
rect 120430 654080 120540 654320
rect 120780 654080 120870 654320
rect 121110 654080 121200 654320
rect 121440 654080 121530 654320
rect 121770 654080 121790 654320
rect 110790 653990 121790 654080
rect 110790 653750 110810 653990
rect 111050 653750 111160 653990
rect 111400 653750 111490 653990
rect 111730 653750 111820 653990
rect 112060 653750 112150 653990
rect 112390 653750 112500 653990
rect 112740 653750 112830 653990
rect 113070 653750 113160 653990
rect 113400 653750 113490 653990
rect 113730 653750 113840 653990
rect 114080 653750 114170 653990
rect 114410 653750 114500 653990
rect 114740 653750 114830 653990
rect 115070 653750 115180 653990
rect 115420 653750 115510 653990
rect 115750 653750 115840 653990
rect 116080 653750 116170 653990
rect 116410 653750 116520 653990
rect 116760 653750 116850 653990
rect 117090 653750 117180 653990
rect 117420 653750 117510 653990
rect 117750 653750 117860 653990
rect 118100 653750 118190 653990
rect 118430 653750 118520 653990
rect 118760 653750 118850 653990
rect 119090 653750 119200 653990
rect 119440 653750 119530 653990
rect 119770 653750 119860 653990
rect 120100 653750 120190 653990
rect 120430 653750 120540 653990
rect 120780 653750 120870 653990
rect 121110 653750 121200 653990
rect 121440 653750 121530 653990
rect 121770 653750 121790 653990
rect 110790 653640 121790 653750
rect 110790 653400 110810 653640
rect 111050 653400 111160 653640
rect 111400 653400 111490 653640
rect 111730 653400 111820 653640
rect 112060 653400 112150 653640
rect 112390 653400 112500 653640
rect 112740 653400 112830 653640
rect 113070 653400 113160 653640
rect 113400 653400 113490 653640
rect 113730 653400 113840 653640
rect 114080 653400 114170 653640
rect 114410 653400 114500 653640
rect 114740 653400 114830 653640
rect 115070 653400 115180 653640
rect 115420 653400 115510 653640
rect 115750 653400 115840 653640
rect 116080 653400 116170 653640
rect 116410 653400 116520 653640
rect 116760 653400 116850 653640
rect 117090 653400 117180 653640
rect 117420 653400 117510 653640
rect 117750 653400 117860 653640
rect 118100 653400 118190 653640
rect 118430 653400 118520 653640
rect 118760 653400 118850 653640
rect 119090 653400 119200 653640
rect 119440 653400 119530 653640
rect 119770 653400 119860 653640
rect 120100 653400 120190 653640
rect 120430 653400 120540 653640
rect 120780 653400 120870 653640
rect 121110 653400 121200 653640
rect 121440 653400 121530 653640
rect 121770 653400 121790 653640
rect 110790 653310 121790 653400
rect 110790 653070 110810 653310
rect 111050 653070 111160 653310
rect 111400 653070 111490 653310
rect 111730 653070 111820 653310
rect 112060 653070 112150 653310
rect 112390 653070 112500 653310
rect 112740 653070 112830 653310
rect 113070 653070 113160 653310
rect 113400 653070 113490 653310
rect 113730 653070 113840 653310
rect 114080 653070 114170 653310
rect 114410 653070 114500 653310
rect 114740 653070 114830 653310
rect 115070 653070 115180 653310
rect 115420 653070 115510 653310
rect 115750 653070 115840 653310
rect 116080 653070 116170 653310
rect 116410 653070 116520 653310
rect 116760 653070 116850 653310
rect 117090 653070 117180 653310
rect 117420 653070 117510 653310
rect 117750 653070 117860 653310
rect 118100 653070 118190 653310
rect 118430 653070 118520 653310
rect 118760 653070 118850 653310
rect 119090 653070 119200 653310
rect 119440 653070 119530 653310
rect 119770 653070 119860 653310
rect 120100 653070 120190 653310
rect 120430 653070 120540 653310
rect 120780 653070 120870 653310
rect 121110 653070 121200 653310
rect 121440 653070 121530 653310
rect 121770 653070 121790 653310
rect 110790 652980 121790 653070
rect 110790 652740 110810 652980
rect 111050 652740 111160 652980
rect 111400 652740 111490 652980
rect 111730 652740 111820 652980
rect 112060 652740 112150 652980
rect 112390 652740 112500 652980
rect 112740 652740 112830 652980
rect 113070 652740 113160 652980
rect 113400 652740 113490 652980
rect 113730 652740 113840 652980
rect 114080 652740 114170 652980
rect 114410 652740 114500 652980
rect 114740 652740 114830 652980
rect 115070 652740 115180 652980
rect 115420 652740 115510 652980
rect 115750 652740 115840 652980
rect 116080 652740 116170 652980
rect 116410 652740 116520 652980
rect 116760 652740 116850 652980
rect 117090 652740 117180 652980
rect 117420 652740 117510 652980
rect 117750 652740 117860 652980
rect 118100 652740 118190 652980
rect 118430 652740 118520 652980
rect 118760 652740 118850 652980
rect 119090 652740 119200 652980
rect 119440 652740 119530 652980
rect 119770 652740 119860 652980
rect 120100 652740 120190 652980
rect 120430 652740 120540 652980
rect 120780 652740 120870 652980
rect 121110 652740 121200 652980
rect 121440 652740 121530 652980
rect 121770 652740 121790 652980
rect 110790 652650 121790 652740
rect 110790 652410 110810 652650
rect 111050 652410 111160 652650
rect 111400 652410 111490 652650
rect 111730 652410 111820 652650
rect 112060 652410 112150 652650
rect 112390 652410 112500 652650
rect 112740 652410 112830 652650
rect 113070 652410 113160 652650
rect 113400 652410 113490 652650
rect 113730 652410 113840 652650
rect 114080 652410 114170 652650
rect 114410 652410 114500 652650
rect 114740 652410 114830 652650
rect 115070 652410 115180 652650
rect 115420 652410 115510 652650
rect 115750 652410 115840 652650
rect 116080 652410 116170 652650
rect 116410 652410 116520 652650
rect 116760 652410 116850 652650
rect 117090 652410 117180 652650
rect 117420 652410 117510 652650
rect 117750 652410 117860 652650
rect 118100 652410 118190 652650
rect 118430 652410 118520 652650
rect 118760 652410 118850 652650
rect 119090 652410 119200 652650
rect 119440 652410 119530 652650
rect 119770 652410 119860 652650
rect 120100 652410 120190 652650
rect 120430 652410 120540 652650
rect 120780 652410 120870 652650
rect 121110 652410 121200 652650
rect 121440 652410 121530 652650
rect 121770 652410 121790 652650
rect 110790 652300 121790 652410
rect 110790 652060 110810 652300
rect 111050 652060 111160 652300
rect 111400 652060 111490 652300
rect 111730 652060 111820 652300
rect 112060 652060 112150 652300
rect 112390 652060 112500 652300
rect 112740 652060 112830 652300
rect 113070 652060 113160 652300
rect 113400 652060 113490 652300
rect 113730 652060 113840 652300
rect 114080 652060 114170 652300
rect 114410 652060 114500 652300
rect 114740 652060 114830 652300
rect 115070 652060 115180 652300
rect 115420 652060 115510 652300
rect 115750 652060 115840 652300
rect 116080 652060 116170 652300
rect 116410 652060 116520 652300
rect 116760 652060 116850 652300
rect 117090 652060 117180 652300
rect 117420 652060 117510 652300
rect 117750 652060 117860 652300
rect 118100 652060 118190 652300
rect 118430 652060 118520 652300
rect 118760 652060 118850 652300
rect 119090 652060 119200 652300
rect 119440 652060 119530 652300
rect 119770 652060 119860 652300
rect 120100 652060 120190 652300
rect 120430 652060 120540 652300
rect 120780 652060 120870 652300
rect 121110 652060 121200 652300
rect 121440 652060 121530 652300
rect 121770 652060 121790 652300
rect 110790 651970 121790 652060
rect 110790 651730 110810 651970
rect 111050 651730 111160 651970
rect 111400 651730 111490 651970
rect 111730 651730 111820 651970
rect 112060 651730 112150 651970
rect 112390 651730 112500 651970
rect 112740 651730 112830 651970
rect 113070 651730 113160 651970
rect 113400 651730 113490 651970
rect 113730 651730 113840 651970
rect 114080 651730 114170 651970
rect 114410 651730 114500 651970
rect 114740 651730 114830 651970
rect 115070 651730 115180 651970
rect 115420 651730 115510 651970
rect 115750 651730 115840 651970
rect 116080 651730 116170 651970
rect 116410 651730 116520 651970
rect 116760 651730 116850 651970
rect 117090 651730 117180 651970
rect 117420 651730 117510 651970
rect 117750 651730 117860 651970
rect 118100 651730 118190 651970
rect 118430 651730 118520 651970
rect 118760 651730 118850 651970
rect 119090 651730 119200 651970
rect 119440 651730 119530 651970
rect 119770 651730 119860 651970
rect 120100 651730 120190 651970
rect 120430 651730 120540 651970
rect 120780 651730 120870 651970
rect 121110 651730 121200 651970
rect 121440 651730 121530 651970
rect 121770 651730 121790 651970
rect 110790 651640 121790 651730
rect 110790 651400 110810 651640
rect 111050 651400 111160 651640
rect 111400 651400 111490 651640
rect 111730 651400 111820 651640
rect 112060 651400 112150 651640
rect 112390 651400 112500 651640
rect 112740 651400 112830 651640
rect 113070 651400 113160 651640
rect 113400 651400 113490 651640
rect 113730 651400 113840 651640
rect 114080 651400 114170 651640
rect 114410 651400 114500 651640
rect 114740 651400 114830 651640
rect 115070 651400 115180 651640
rect 115420 651400 115510 651640
rect 115750 651400 115840 651640
rect 116080 651400 116170 651640
rect 116410 651400 116520 651640
rect 116760 651400 116850 651640
rect 117090 651400 117180 651640
rect 117420 651400 117510 651640
rect 117750 651400 117860 651640
rect 118100 651400 118190 651640
rect 118430 651400 118520 651640
rect 118760 651400 118850 651640
rect 119090 651400 119200 651640
rect 119440 651400 119530 651640
rect 119770 651400 119860 651640
rect 120100 651400 120190 651640
rect 120430 651400 120540 651640
rect 120780 651400 120870 651640
rect 121110 651400 121200 651640
rect 121440 651400 121530 651640
rect 121770 651400 121790 651640
rect 110790 651310 121790 651400
rect 110790 651070 110810 651310
rect 111050 651070 111160 651310
rect 111400 651070 111490 651310
rect 111730 651070 111820 651310
rect 112060 651070 112150 651310
rect 112390 651070 112500 651310
rect 112740 651070 112830 651310
rect 113070 651070 113160 651310
rect 113400 651070 113490 651310
rect 113730 651070 113840 651310
rect 114080 651070 114170 651310
rect 114410 651070 114500 651310
rect 114740 651070 114830 651310
rect 115070 651070 115180 651310
rect 115420 651070 115510 651310
rect 115750 651070 115840 651310
rect 116080 651070 116170 651310
rect 116410 651070 116520 651310
rect 116760 651070 116850 651310
rect 117090 651070 117180 651310
rect 117420 651070 117510 651310
rect 117750 651070 117860 651310
rect 118100 651070 118190 651310
rect 118430 651070 118520 651310
rect 118760 651070 118850 651310
rect 119090 651070 119200 651310
rect 119440 651070 119530 651310
rect 119770 651070 119860 651310
rect 120100 651070 120190 651310
rect 120430 651070 120540 651310
rect 120780 651070 120870 651310
rect 121110 651070 121200 651310
rect 121440 651070 121530 651310
rect 121770 651070 121790 651310
rect 110790 650960 121790 651070
rect 110790 650720 110810 650960
rect 111050 650720 111160 650960
rect 111400 650720 111490 650960
rect 111730 650720 111820 650960
rect 112060 650720 112150 650960
rect 112390 650720 112500 650960
rect 112740 650720 112830 650960
rect 113070 650720 113160 650960
rect 113400 650720 113490 650960
rect 113730 650720 113840 650960
rect 114080 650720 114170 650960
rect 114410 650720 114500 650960
rect 114740 650720 114830 650960
rect 115070 650720 115180 650960
rect 115420 650720 115510 650960
rect 115750 650720 115840 650960
rect 116080 650720 116170 650960
rect 116410 650720 116520 650960
rect 116760 650720 116850 650960
rect 117090 650720 117180 650960
rect 117420 650720 117510 650960
rect 117750 650720 117860 650960
rect 118100 650720 118190 650960
rect 118430 650720 118520 650960
rect 118760 650720 118850 650960
rect 119090 650720 119200 650960
rect 119440 650720 119530 650960
rect 119770 650720 119860 650960
rect 120100 650720 120190 650960
rect 120430 650720 120540 650960
rect 120780 650720 120870 650960
rect 121110 650720 121200 650960
rect 121440 650720 121530 650960
rect 121770 650720 121790 650960
rect 110790 650630 121790 650720
rect 110790 650390 110810 650630
rect 111050 650390 111160 650630
rect 111400 650390 111490 650630
rect 111730 650390 111820 650630
rect 112060 650390 112150 650630
rect 112390 650390 112500 650630
rect 112740 650390 112830 650630
rect 113070 650390 113160 650630
rect 113400 650390 113490 650630
rect 113730 650390 113840 650630
rect 114080 650390 114170 650630
rect 114410 650390 114500 650630
rect 114740 650390 114830 650630
rect 115070 650390 115180 650630
rect 115420 650390 115510 650630
rect 115750 650390 115840 650630
rect 116080 650390 116170 650630
rect 116410 650390 116520 650630
rect 116760 650390 116850 650630
rect 117090 650390 117180 650630
rect 117420 650390 117510 650630
rect 117750 650390 117860 650630
rect 118100 650390 118190 650630
rect 118430 650390 118520 650630
rect 118760 650390 118850 650630
rect 119090 650390 119200 650630
rect 119440 650390 119530 650630
rect 119770 650390 119860 650630
rect 120100 650390 120190 650630
rect 120430 650390 120540 650630
rect 120780 650390 120870 650630
rect 121110 650390 121200 650630
rect 121440 650390 121530 650630
rect 121770 650390 121790 650630
rect 110790 650300 121790 650390
rect 110790 650060 110810 650300
rect 111050 650060 111160 650300
rect 111400 650060 111490 650300
rect 111730 650060 111820 650300
rect 112060 650060 112150 650300
rect 112390 650060 112500 650300
rect 112740 650060 112830 650300
rect 113070 650060 113160 650300
rect 113400 650060 113490 650300
rect 113730 650060 113840 650300
rect 114080 650060 114170 650300
rect 114410 650060 114500 650300
rect 114740 650060 114830 650300
rect 115070 650060 115180 650300
rect 115420 650060 115510 650300
rect 115750 650060 115840 650300
rect 116080 650060 116170 650300
rect 116410 650060 116520 650300
rect 116760 650060 116850 650300
rect 117090 650060 117180 650300
rect 117420 650060 117510 650300
rect 117750 650060 117860 650300
rect 118100 650060 118190 650300
rect 118430 650060 118520 650300
rect 118760 650060 118850 650300
rect 119090 650060 119200 650300
rect 119440 650060 119530 650300
rect 119770 650060 119860 650300
rect 120100 650060 120190 650300
rect 120430 650060 120540 650300
rect 120780 650060 120870 650300
rect 121110 650060 121200 650300
rect 121440 650060 121530 650300
rect 121770 650060 121790 650300
rect 110790 649970 121790 650060
rect 110790 649730 110810 649970
rect 111050 649730 111160 649970
rect 111400 649730 111490 649970
rect 111730 649730 111820 649970
rect 112060 649730 112150 649970
rect 112390 649730 112500 649970
rect 112740 649730 112830 649970
rect 113070 649730 113160 649970
rect 113400 649730 113490 649970
rect 113730 649730 113840 649970
rect 114080 649730 114170 649970
rect 114410 649730 114500 649970
rect 114740 649730 114830 649970
rect 115070 649730 115180 649970
rect 115420 649730 115510 649970
rect 115750 649730 115840 649970
rect 116080 649730 116170 649970
rect 116410 649730 116520 649970
rect 116760 649730 116850 649970
rect 117090 649730 117180 649970
rect 117420 649730 117510 649970
rect 117750 649730 117860 649970
rect 118100 649730 118190 649970
rect 118430 649730 118520 649970
rect 118760 649730 118850 649970
rect 119090 649730 119200 649970
rect 119440 649730 119530 649970
rect 119770 649730 119860 649970
rect 120100 649730 120190 649970
rect 120430 649730 120540 649970
rect 120780 649730 120870 649970
rect 121110 649730 121200 649970
rect 121440 649730 121530 649970
rect 121770 649730 121790 649970
rect 110790 649620 121790 649730
rect 110790 649380 110810 649620
rect 111050 649380 111160 649620
rect 111400 649380 111490 649620
rect 111730 649380 111820 649620
rect 112060 649380 112150 649620
rect 112390 649380 112500 649620
rect 112740 649380 112830 649620
rect 113070 649380 113160 649620
rect 113400 649380 113490 649620
rect 113730 649380 113840 649620
rect 114080 649380 114170 649620
rect 114410 649380 114500 649620
rect 114740 649380 114830 649620
rect 115070 649380 115180 649620
rect 115420 649380 115510 649620
rect 115750 649380 115840 649620
rect 116080 649380 116170 649620
rect 116410 649380 116520 649620
rect 116760 649380 116850 649620
rect 117090 649380 117180 649620
rect 117420 649380 117510 649620
rect 117750 649380 117860 649620
rect 118100 649380 118190 649620
rect 118430 649380 118520 649620
rect 118760 649380 118850 649620
rect 119090 649380 119200 649620
rect 119440 649380 119530 649620
rect 119770 649380 119860 649620
rect 120100 649380 120190 649620
rect 120430 649380 120540 649620
rect 120780 649380 120870 649620
rect 121110 649380 121200 649620
rect 121440 649380 121530 649620
rect 121770 649380 121790 649620
rect 110790 649360 121790 649380
rect 122170 660340 133170 660360
rect 122170 660100 122190 660340
rect 122430 660100 122540 660340
rect 122780 660100 122870 660340
rect 123110 660100 123200 660340
rect 123440 660100 123530 660340
rect 123770 660100 123880 660340
rect 124120 660100 124210 660340
rect 124450 660100 124540 660340
rect 124780 660100 124870 660340
rect 125110 660100 125220 660340
rect 125460 660100 125550 660340
rect 125790 660100 125880 660340
rect 126120 660100 126210 660340
rect 126450 660100 126560 660340
rect 126800 660100 126890 660340
rect 127130 660100 127220 660340
rect 127460 660100 127550 660340
rect 127790 660100 127900 660340
rect 128140 660100 128230 660340
rect 128470 660100 128560 660340
rect 128800 660100 128890 660340
rect 129130 660100 129240 660340
rect 129480 660100 129570 660340
rect 129810 660100 129900 660340
rect 130140 660100 130230 660340
rect 130470 660100 130580 660340
rect 130820 660100 130910 660340
rect 131150 660100 131240 660340
rect 131480 660100 131570 660340
rect 131810 660100 131920 660340
rect 132160 660100 132250 660340
rect 132490 660100 132580 660340
rect 132820 660100 132910 660340
rect 133150 660100 133170 660340
rect 122170 660010 133170 660100
rect 122170 659770 122190 660010
rect 122430 659770 122540 660010
rect 122780 659770 122870 660010
rect 123110 659770 123200 660010
rect 123440 659770 123530 660010
rect 123770 659770 123880 660010
rect 124120 659770 124210 660010
rect 124450 659770 124540 660010
rect 124780 659770 124870 660010
rect 125110 659770 125220 660010
rect 125460 659770 125550 660010
rect 125790 659770 125880 660010
rect 126120 659770 126210 660010
rect 126450 659770 126560 660010
rect 126800 659770 126890 660010
rect 127130 659770 127220 660010
rect 127460 659770 127550 660010
rect 127790 659770 127900 660010
rect 128140 659770 128230 660010
rect 128470 659770 128560 660010
rect 128800 659770 128890 660010
rect 129130 659770 129240 660010
rect 129480 659770 129570 660010
rect 129810 659770 129900 660010
rect 130140 659770 130230 660010
rect 130470 659770 130580 660010
rect 130820 659770 130910 660010
rect 131150 659770 131240 660010
rect 131480 659770 131570 660010
rect 131810 659770 131920 660010
rect 132160 659770 132250 660010
rect 132490 659770 132580 660010
rect 132820 659770 132910 660010
rect 133150 659770 133170 660010
rect 122170 659680 133170 659770
rect 122170 659440 122190 659680
rect 122430 659440 122540 659680
rect 122780 659440 122870 659680
rect 123110 659440 123200 659680
rect 123440 659440 123530 659680
rect 123770 659440 123880 659680
rect 124120 659440 124210 659680
rect 124450 659440 124540 659680
rect 124780 659440 124870 659680
rect 125110 659440 125220 659680
rect 125460 659440 125550 659680
rect 125790 659440 125880 659680
rect 126120 659440 126210 659680
rect 126450 659440 126560 659680
rect 126800 659440 126890 659680
rect 127130 659440 127220 659680
rect 127460 659440 127550 659680
rect 127790 659440 127900 659680
rect 128140 659440 128230 659680
rect 128470 659440 128560 659680
rect 128800 659440 128890 659680
rect 129130 659440 129240 659680
rect 129480 659440 129570 659680
rect 129810 659440 129900 659680
rect 130140 659440 130230 659680
rect 130470 659440 130580 659680
rect 130820 659440 130910 659680
rect 131150 659440 131240 659680
rect 131480 659440 131570 659680
rect 131810 659440 131920 659680
rect 132160 659440 132250 659680
rect 132490 659440 132580 659680
rect 132820 659440 132910 659680
rect 133150 659440 133170 659680
rect 122170 659350 133170 659440
rect 122170 659110 122190 659350
rect 122430 659110 122540 659350
rect 122780 659110 122870 659350
rect 123110 659110 123200 659350
rect 123440 659110 123530 659350
rect 123770 659110 123880 659350
rect 124120 659110 124210 659350
rect 124450 659110 124540 659350
rect 124780 659110 124870 659350
rect 125110 659110 125220 659350
rect 125460 659110 125550 659350
rect 125790 659110 125880 659350
rect 126120 659110 126210 659350
rect 126450 659110 126560 659350
rect 126800 659110 126890 659350
rect 127130 659110 127220 659350
rect 127460 659110 127550 659350
rect 127790 659110 127900 659350
rect 128140 659110 128230 659350
rect 128470 659110 128560 659350
rect 128800 659110 128890 659350
rect 129130 659110 129240 659350
rect 129480 659110 129570 659350
rect 129810 659110 129900 659350
rect 130140 659110 130230 659350
rect 130470 659110 130580 659350
rect 130820 659110 130910 659350
rect 131150 659110 131240 659350
rect 131480 659110 131570 659350
rect 131810 659110 131920 659350
rect 132160 659110 132250 659350
rect 132490 659110 132580 659350
rect 132820 659110 132910 659350
rect 133150 659110 133170 659350
rect 122170 659000 133170 659110
rect 122170 658760 122190 659000
rect 122430 658760 122540 659000
rect 122780 658760 122870 659000
rect 123110 658760 123200 659000
rect 123440 658760 123530 659000
rect 123770 658760 123880 659000
rect 124120 658760 124210 659000
rect 124450 658760 124540 659000
rect 124780 658760 124870 659000
rect 125110 658760 125220 659000
rect 125460 658760 125550 659000
rect 125790 658760 125880 659000
rect 126120 658760 126210 659000
rect 126450 658760 126560 659000
rect 126800 658760 126890 659000
rect 127130 658760 127220 659000
rect 127460 658760 127550 659000
rect 127790 658760 127900 659000
rect 128140 658760 128230 659000
rect 128470 658760 128560 659000
rect 128800 658760 128890 659000
rect 129130 658760 129240 659000
rect 129480 658760 129570 659000
rect 129810 658760 129900 659000
rect 130140 658760 130230 659000
rect 130470 658760 130580 659000
rect 130820 658760 130910 659000
rect 131150 658760 131240 659000
rect 131480 658760 131570 659000
rect 131810 658760 131920 659000
rect 132160 658760 132250 659000
rect 132490 658760 132580 659000
rect 132820 658760 132910 659000
rect 133150 658760 133170 659000
rect 122170 658670 133170 658760
rect 122170 658430 122190 658670
rect 122430 658430 122540 658670
rect 122780 658430 122870 658670
rect 123110 658430 123200 658670
rect 123440 658430 123530 658670
rect 123770 658430 123880 658670
rect 124120 658430 124210 658670
rect 124450 658430 124540 658670
rect 124780 658430 124870 658670
rect 125110 658430 125220 658670
rect 125460 658430 125550 658670
rect 125790 658430 125880 658670
rect 126120 658430 126210 658670
rect 126450 658430 126560 658670
rect 126800 658430 126890 658670
rect 127130 658430 127220 658670
rect 127460 658430 127550 658670
rect 127790 658430 127900 658670
rect 128140 658430 128230 658670
rect 128470 658430 128560 658670
rect 128800 658430 128890 658670
rect 129130 658430 129240 658670
rect 129480 658430 129570 658670
rect 129810 658430 129900 658670
rect 130140 658430 130230 658670
rect 130470 658430 130580 658670
rect 130820 658430 130910 658670
rect 131150 658430 131240 658670
rect 131480 658430 131570 658670
rect 131810 658430 131920 658670
rect 132160 658430 132250 658670
rect 132490 658430 132580 658670
rect 132820 658430 132910 658670
rect 133150 658430 133170 658670
rect 122170 658340 133170 658430
rect 122170 658100 122190 658340
rect 122430 658100 122540 658340
rect 122780 658100 122870 658340
rect 123110 658100 123200 658340
rect 123440 658100 123530 658340
rect 123770 658100 123880 658340
rect 124120 658100 124210 658340
rect 124450 658100 124540 658340
rect 124780 658100 124870 658340
rect 125110 658100 125220 658340
rect 125460 658100 125550 658340
rect 125790 658100 125880 658340
rect 126120 658100 126210 658340
rect 126450 658100 126560 658340
rect 126800 658100 126890 658340
rect 127130 658100 127220 658340
rect 127460 658100 127550 658340
rect 127790 658100 127900 658340
rect 128140 658100 128230 658340
rect 128470 658100 128560 658340
rect 128800 658100 128890 658340
rect 129130 658100 129240 658340
rect 129480 658100 129570 658340
rect 129810 658100 129900 658340
rect 130140 658100 130230 658340
rect 130470 658100 130580 658340
rect 130820 658100 130910 658340
rect 131150 658100 131240 658340
rect 131480 658100 131570 658340
rect 131810 658100 131920 658340
rect 132160 658100 132250 658340
rect 132490 658100 132580 658340
rect 132820 658100 132910 658340
rect 133150 658100 133170 658340
rect 122170 658010 133170 658100
rect 122170 657770 122190 658010
rect 122430 657770 122540 658010
rect 122780 657770 122870 658010
rect 123110 657770 123200 658010
rect 123440 657770 123530 658010
rect 123770 657770 123880 658010
rect 124120 657770 124210 658010
rect 124450 657770 124540 658010
rect 124780 657770 124870 658010
rect 125110 657770 125220 658010
rect 125460 657770 125550 658010
rect 125790 657770 125880 658010
rect 126120 657770 126210 658010
rect 126450 657770 126560 658010
rect 126800 657770 126890 658010
rect 127130 657770 127220 658010
rect 127460 657770 127550 658010
rect 127790 657770 127900 658010
rect 128140 657770 128230 658010
rect 128470 657770 128560 658010
rect 128800 657770 128890 658010
rect 129130 657770 129240 658010
rect 129480 657770 129570 658010
rect 129810 657770 129900 658010
rect 130140 657770 130230 658010
rect 130470 657770 130580 658010
rect 130820 657770 130910 658010
rect 131150 657770 131240 658010
rect 131480 657770 131570 658010
rect 131810 657770 131920 658010
rect 132160 657770 132250 658010
rect 132490 657770 132580 658010
rect 132820 657770 132910 658010
rect 133150 657770 133170 658010
rect 122170 657660 133170 657770
rect 122170 657420 122190 657660
rect 122430 657420 122540 657660
rect 122780 657420 122870 657660
rect 123110 657420 123200 657660
rect 123440 657420 123530 657660
rect 123770 657420 123880 657660
rect 124120 657420 124210 657660
rect 124450 657420 124540 657660
rect 124780 657420 124870 657660
rect 125110 657420 125220 657660
rect 125460 657420 125550 657660
rect 125790 657420 125880 657660
rect 126120 657420 126210 657660
rect 126450 657420 126560 657660
rect 126800 657420 126890 657660
rect 127130 657420 127220 657660
rect 127460 657420 127550 657660
rect 127790 657420 127900 657660
rect 128140 657420 128230 657660
rect 128470 657420 128560 657660
rect 128800 657420 128890 657660
rect 129130 657420 129240 657660
rect 129480 657420 129570 657660
rect 129810 657420 129900 657660
rect 130140 657420 130230 657660
rect 130470 657420 130580 657660
rect 130820 657420 130910 657660
rect 131150 657420 131240 657660
rect 131480 657420 131570 657660
rect 131810 657420 131920 657660
rect 132160 657420 132250 657660
rect 132490 657420 132580 657660
rect 132820 657420 132910 657660
rect 133150 657420 133170 657660
rect 122170 657330 133170 657420
rect 122170 657090 122190 657330
rect 122430 657090 122540 657330
rect 122780 657090 122870 657330
rect 123110 657090 123200 657330
rect 123440 657090 123530 657330
rect 123770 657090 123880 657330
rect 124120 657090 124210 657330
rect 124450 657090 124540 657330
rect 124780 657090 124870 657330
rect 125110 657090 125220 657330
rect 125460 657090 125550 657330
rect 125790 657090 125880 657330
rect 126120 657090 126210 657330
rect 126450 657090 126560 657330
rect 126800 657090 126890 657330
rect 127130 657090 127220 657330
rect 127460 657090 127550 657330
rect 127790 657090 127900 657330
rect 128140 657090 128230 657330
rect 128470 657090 128560 657330
rect 128800 657090 128890 657330
rect 129130 657090 129240 657330
rect 129480 657090 129570 657330
rect 129810 657090 129900 657330
rect 130140 657090 130230 657330
rect 130470 657090 130580 657330
rect 130820 657090 130910 657330
rect 131150 657090 131240 657330
rect 131480 657090 131570 657330
rect 131810 657090 131920 657330
rect 132160 657090 132250 657330
rect 132490 657090 132580 657330
rect 132820 657090 132910 657330
rect 133150 657090 133170 657330
rect 122170 657000 133170 657090
rect 122170 656760 122190 657000
rect 122430 656760 122540 657000
rect 122780 656760 122870 657000
rect 123110 656760 123200 657000
rect 123440 656760 123530 657000
rect 123770 656760 123880 657000
rect 124120 656760 124210 657000
rect 124450 656760 124540 657000
rect 124780 656760 124870 657000
rect 125110 656760 125220 657000
rect 125460 656760 125550 657000
rect 125790 656760 125880 657000
rect 126120 656760 126210 657000
rect 126450 656760 126560 657000
rect 126800 656760 126890 657000
rect 127130 656760 127220 657000
rect 127460 656760 127550 657000
rect 127790 656760 127900 657000
rect 128140 656760 128230 657000
rect 128470 656760 128560 657000
rect 128800 656760 128890 657000
rect 129130 656760 129240 657000
rect 129480 656760 129570 657000
rect 129810 656760 129900 657000
rect 130140 656760 130230 657000
rect 130470 656760 130580 657000
rect 130820 656760 130910 657000
rect 131150 656760 131240 657000
rect 131480 656760 131570 657000
rect 131810 656760 131920 657000
rect 132160 656760 132250 657000
rect 132490 656760 132580 657000
rect 132820 656760 132910 657000
rect 133150 656760 133170 657000
rect 122170 656670 133170 656760
rect 122170 656430 122190 656670
rect 122430 656430 122540 656670
rect 122780 656430 122870 656670
rect 123110 656430 123200 656670
rect 123440 656430 123530 656670
rect 123770 656430 123880 656670
rect 124120 656430 124210 656670
rect 124450 656430 124540 656670
rect 124780 656430 124870 656670
rect 125110 656430 125220 656670
rect 125460 656430 125550 656670
rect 125790 656430 125880 656670
rect 126120 656430 126210 656670
rect 126450 656430 126560 656670
rect 126800 656430 126890 656670
rect 127130 656430 127220 656670
rect 127460 656430 127550 656670
rect 127790 656430 127900 656670
rect 128140 656430 128230 656670
rect 128470 656430 128560 656670
rect 128800 656430 128890 656670
rect 129130 656430 129240 656670
rect 129480 656430 129570 656670
rect 129810 656430 129900 656670
rect 130140 656430 130230 656670
rect 130470 656430 130580 656670
rect 130820 656430 130910 656670
rect 131150 656430 131240 656670
rect 131480 656430 131570 656670
rect 131810 656430 131920 656670
rect 132160 656430 132250 656670
rect 132490 656430 132580 656670
rect 132820 656430 132910 656670
rect 133150 656430 133170 656670
rect 122170 656320 133170 656430
rect 122170 656080 122190 656320
rect 122430 656080 122540 656320
rect 122780 656080 122870 656320
rect 123110 656080 123200 656320
rect 123440 656080 123530 656320
rect 123770 656080 123880 656320
rect 124120 656080 124210 656320
rect 124450 656080 124540 656320
rect 124780 656080 124870 656320
rect 125110 656080 125220 656320
rect 125460 656080 125550 656320
rect 125790 656080 125880 656320
rect 126120 656080 126210 656320
rect 126450 656080 126560 656320
rect 126800 656080 126890 656320
rect 127130 656080 127220 656320
rect 127460 656080 127550 656320
rect 127790 656080 127900 656320
rect 128140 656080 128230 656320
rect 128470 656080 128560 656320
rect 128800 656080 128890 656320
rect 129130 656080 129240 656320
rect 129480 656080 129570 656320
rect 129810 656080 129900 656320
rect 130140 656080 130230 656320
rect 130470 656080 130580 656320
rect 130820 656080 130910 656320
rect 131150 656080 131240 656320
rect 131480 656080 131570 656320
rect 131810 656080 131920 656320
rect 132160 656080 132250 656320
rect 132490 656080 132580 656320
rect 132820 656080 132910 656320
rect 133150 656080 133170 656320
rect 122170 655990 133170 656080
rect 122170 655750 122190 655990
rect 122430 655750 122540 655990
rect 122780 655750 122870 655990
rect 123110 655750 123200 655990
rect 123440 655750 123530 655990
rect 123770 655750 123880 655990
rect 124120 655750 124210 655990
rect 124450 655750 124540 655990
rect 124780 655750 124870 655990
rect 125110 655750 125220 655990
rect 125460 655750 125550 655990
rect 125790 655750 125880 655990
rect 126120 655750 126210 655990
rect 126450 655750 126560 655990
rect 126800 655750 126890 655990
rect 127130 655750 127220 655990
rect 127460 655750 127550 655990
rect 127790 655750 127900 655990
rect 128140 655750 128230 655990
rect 128470 655750 128560 655990
rect 128800 655750 128890 655990
rect 129130 655750 129240 655990
rect 129480 655750 129570 655990
rect 129810 655750 129900 655990
rect 130140 655750 130230 655990
rect 130470 655750 130580 655990
rect 130820 655750 130910 655990
rect 131150 655750 131240 655990
rect 131480 655750 131570 655990
rect 131810 655750 131920 655990
rect 132160 655750 132250 655990
rect 132490 655750 132580 655990
rect 132820 655750 132910 655990
rect 133150 655750 133170 655990
rect 122170 655660 133170 655750
rect 122170 655420 122190 655660
rect 122430 655420 122540 655660
rect 122780 655420 122870 655660
rect 123110 655420 123200 655660
rect 123440 655420 123530 655660
rect 123770 655420 123880 655660
rect 124120 655420 124210 655660
rect 124450 655420 124540 655660
rect 124780 655420 124870 655660
rect 125110 655420 125220 655660
rect 125460 655420 125550 655660
rect 125790 655420 125880 655660
rect 126120 655420 126210 655660
rect 126450 655420 126560 655660
rect 126800 655420 126890 655660
rect 127130 655420 127220 655660
rect 127460 655420 127550 655660
rect 127790 655420 127900 655660
rect 128140 655420 128230 655660
rect 128470 655420 128560 655660
rect 128800 655420 128890 655660
rect 129130 655420 129240 655660
rect 129480 655420 129570 655660
rect 129810 655420 129900 655660
rect 130140 655420 130230 655660
rect 130470 655420 130580 655660
rect 130820 655420 130910 655660
rect 131150 655420 131240 655660
rect 131480 655420 131570 655660
rect 131810 655420 131920 655660
rect 132160 655420 132250 655660
rect 132490 655420 132580 655660
rect 132820 655420 132910 655660
rect 133150 655420 133170 655660
rect 122170 655330 133170 655420
rect 122170 655090 122190 655330
rect 122430 655090 122540 655330
rect 122780 655090 122870 655330
rect 123110 655090 123200 655330
rect 123440 655090 123530 655330
rect 123770 655090 123880 655330
rect 124120 655090 124210 655330
rect 124450 655090 124540 655330
rect 124780 655090 124870 655330
rect 125110 655090 125220 655330
rect 125460 655090 125550 655330
rect 125790 655090 125880 655330
rect 126120 655090 126210 655330
rect 126450 655090 126560 655330
rect 126800 655090 126890 655330
rect 127130 655090 127220 655330
rect 127460 655090 127550 655330
rect 127790 655090 127900 655330
rect 128140 655090 128230 655330
rect 128470 655090 128560 655330
rect 128800 655090 128890 655330
rect 129130 655090 129240 655330
rect 129480 655090 129570 655330
rect 129810 655090 129900 655330
rect 130140 655090 130230 655330
rect 130470 655090 130580 655330
rect 130820 655090 130910 655330
rect 131150 655090 131240 655330
rect 131480 655090 131570 655330
rect 131810 655090 131920 655330
rect 132160 655090 132250 655330
rect 132490 655090 132580 655330
rect 132820 655090 132910 655330
rect 133150 655090 133170 655330
rect 122170 654980 133170 655090
rect 122170 654740 122190 654980
rect 122430 654740 122540 654980
rect 122780 654740 122870 654980
rect 123110 654740 123200 654980
rect 123440 654740 123530 654980
rect 123770 654740 123880 654980
rect 124120 654740 124210 654980
rect 124450 654740 124540 654980
rect 124780 654740 124870 654980
rect 125110 654740 125220 654980
rect 125460 654740 125550 654980
rect 125790 654740 125880 654980
rect 126120 654740 126210 654980
rect 126450 654740 126560 654980
rect 126800 654740 126890 654980
rect 127130 654740 127220 654980
rect 127460 654740 127550 654980
rect 127790 654740 127900 654980
rect 128140 654740 128230 654980
rect 128470 654740 128560 654980
rect 128800 654740 128890 654980
rect 129130 654740 129240 654980
rect 129480 654740 129570 654980
rect 129810 654740 129900 654980
rect 130140 654740 130230 654980
rect 130470 654740 130580 654980
rect 130820 654740 130910 654980
rect 131150 654740 131240 654980
rect 131480 654740 131570 654980
rect 131810 654740 131920 654980
rect 132160 654740 132250 654980
rect 132490 654740 132580 654980
rect 132820 654740 132910 654980
rect 133150 654740 133170 654980
rect 122170 654650 133170 654740
rect 122170 654410 122190 654650
rect 122430 654410 122540 654650
rect 122780 654410 122870 654650
rect 123110 654410 123200 654650
rect 123440 654410 123530 654650
rect 123770 654410 123880 654650
rect 124120 654410 124210 654650
rect 124450 654410 124540 654650
rect 124780 654410 124870 654650
rect 125110 654410 125220 654650
rect 125460 654410 125550 654650
rect 125790 654410 125880 654650
rect 126120 654410 126210 654650
rect 126450 654410 126560 654650
rect 126800 654410 126890 654650
rect 127130 654410 127220 654650
rect 127460 654410 127550 654650
rect 127790 654410 127900 654650
rect 128140 654410 128230 654650
rect 128470 654410 128560 654650
rect 128800 654410 128890 654650
rect 129130 654410 129240 654650
rect 129480 654410 129570 654650
rect 129810 654410 129900 654650
rect 130140 654410 130230 654650
rect 130470 654410 130580 654650
rect 130820 654410 130910 654650
rect 131150 654410 131240 654650
rect 131480 654410 131570 654650
rect 131810 654410 131920 654650
rect 132160 654410 132250 654650
rect 132490 654410 132580 654650
rect 132820 654410 132910 654650
rect 133150 654410 133170 654650
rect 122170 654320 133170 654410
rect 122170 654080 122190 654320
rect 122430 654080 122540 654320
rect 122780 654080 122870 654320
rect 123110 654080 123200 654320
rect 123440 654080 123530 654320
rect 123770 654080 123880 654320
rect 124120 654080 124210 654320
rect 124450 654080 124540 654320
rect 124780 654080 124870 654320
rect 125110 654080 125220 654320
rect 125460 654080 125550 654320
rect 125790 654080 125880 654320
rect 126120 654080 126210 654320
rect 126450 654080 126560 654320
rect 126800 654080 126890 654320
rect 127130 654080 127220 654320
rect 127460 654080 127550 654320
rect 127790 654080 127900 654320
rect 128140 654080 128230 654320
rect 128470 654080 128560 654320
rect 128800 654080 128890 654320
rect 129130 654080 129240 654320
rect 129480 654080 129570 654320
rect 129810 654080 129900 654320
rect 130140 654080 130230 654320
rect 130470 654080 130580 654320
rect 130820 654080 130910 654320
rect 131150 654080 131240 654320
rect 131480 654080 131570 654320
rect 131810 654080 131920 654320
rect 132160 654080 132250 654320
rect 132490 654080 132580 654320
rect 132820 654080 132910 654320
rect 133150 654080 133170 654320
rect 122170 653990 133170 654080
rect 122170 653750 122190 653990
rect 122430 653750 122540 653990
rect 122780 653750 122870 653990
rect 123110 653750 123200 653990
rect 123440 653750 123530 653990
rect 123770 653750 123880 653990
rect 124120 653750 124210 653990
rect 124450 653750 124540 653990
rect 124780 653750 124870 653990
rect 125110 653750 125220 653990
rect 125460 653750 125550 653990
rect 125790 653750 125880 653990
rect 126120 653750 126210 653990
rect 126450 653750 126560 653990
rect 126800 653750 126890 653990
rect 127130 653750 127220 653990
rect 127460 653750 127550 653990
rect 127790 653750 127900 653990
rect 128140 653750 128230 653990
rect 128470 653750 128560 653990
rect 128800 653750 128890 653990
rect 129130 653750 129240 653990
rect 129480 653750 129570 653990
rect 129810 653750 129900 653990
rect 130140 653750 130230 653990
rect 130470 653750 130580 653990
rect 130820 653750 130910 653990
rect 131150 653750 131240 653990
rect 131480 653750 131570 653990
rect 131810 653750 131920 653990
rect 132160 653750 132250 653990
rect 132490 653750 132580 653990
rect 132820 653750 132910 653990
rect 133150 653750 133170 653990
rect 122170 653640 133170 653750
rect 122170 653400 122190 653640
rect 122430 653400 122540 653640
rect 122780 653400 122870 653640
rect 123110 653400 123200 653640
rect 123440 653400 123530 653640
rect 123770 653400 123880 653640
rect 124120 653400 124210 653640
rect 124450 653400 124540 653640
rect 124780 653400 124870 653640
rect 125110 653400 125220 653640
rect 125460 653400 125550 653640
rect 125790 653400 125880 653640
rect 126120 653400 126210 653640
rect 126450 653400 126560 653640
rect 126800 653400 126890 653640
rect 127130 653400 127220 653640
rect 127460 653400 127550 653640
rect 127790 653400 127900 653640
rect 128140 653400 128230 653640
rect 128470 653400 128560 653640
rect 128800 653400 128890 653640
rect 129130 653400 129240 653640
rect 129480 653400 129570 653640
rect 129810 653400 129900 653640
rect 130140 653400 130230 653640
rect 130470 653400 130580 653640
rect 130820 653400 130910 653640
rect 131150 653400 131240 653640
rect 131480 653400 131570 653640
rect 131810 653400 131920 653640
rect 132160 653400 132250 653640
rect 132490 653400 132580 653640
rect 132820 653400 132910 653640
rect 133150 653400 133170 653640
rect 122170 653310 133170 653400
rect 122170 653070 122190 653310
rect 122430 653070 122540 653310
rect 122780 653070 122870 653310
rect 123110 653070 123200 653310
rect 123440 653070 123530 653310
rect 123770 653070 123880 653310
rect 124120 653070 124210 653310
rect 124450 653070 124540 653310
rect 124780 653070 124870 653310
rect 125110 653070 125220 653310
rect 125460 653070 125550 653310
rect 125790 653070 125880 653310
rect 126120 653070 126210 653310
rect 126450 653070 126560 653310
rect 126800 653070 126890 653310
rect 127130 653070 127220 653310
rect 127460 653070 127550 653310
rect 127790 653070 127900 653310
rect 128140 653070 128230 653310
rect 128470 653070 128560 653310
rect 128800 653070 128890 653310
rect 129130 653070 129240 653310
rect 129480 653070 129570 653310
rect 129810 653070 129900 653310
rect 130140 653070 130230 653310
rect 130470 653070 130580 653310
rect 130820 653070 130910 653310
rect 131150 653070 131240 653310
rect 131480 653070 131570 653310
rect 131810 653070 131920 653310
rect 132160 653070 132250 653310
rect 132490 653070 132580 653310
rect 132820 653070 132910 653310
rect 133150 653070 133170 653310
rect 122170 652980 133170 653070
rect 122170 652740 122190 652980
rect 122430 652740 122540 652980
rect 122780 652740 122870 652980
rect 123110 652740 123200 652980
rect 123440 652740 123530 652980
rect 123770 652740 123880 652980
rect 124120 652740 124210 652980
rect 124450 652740 124540 652980
rect 124780 652740 124870 652980
rect 125110 652740 125220 652980
rect 125460 652740 125550 652980
rect 125790 652740 125880 652980
rect 126120 652740 126210 652980
rect 126450 652740 126560 652980
rect 126800 652740 126890 652980
rect 127130 652740 127220 652980
rect 127460 652740 127550 652980
rect 127790 652740 127900 652980
rect 128140 652740 128230 652980
rect 128470 652740 128560 652980
rect 128800 652740 128890 652980
rect 129130 652740 129240 652980
rect 129480 652740 129570 652980
rect 129810 652740 129900 652980
rect 130140 652740 130230 652980
rect 130470 652740 130580 652980
rect 130820 652740 130910 652980
rect 131150 652740 131240 652980
rect 131480 652740 131570 652980
rect 131810 652740 131920 652980
rect 132160 652740 132250 652980
rect 132490 652740 132580 652980
rect 132820 652740 132910 652980
rect 133150 652740 133170 652980
rect 122170 652650 133170 652740
rect 122170 652410 122190 652650
rect 122430 652410 122540 652650
rect 122780 652410 122870 652650
rect 123110 652410 123200 652650
rect 123440 652410 123530 652650
rect 123770 652410 123880 652650
rect 124120 652410 124210 652650
rect 124450 652410 124540 652650
rect 124780 652410 124870 652650
rect 125110 652410 125220 652650
rect 125460 652410 125550 652650
rect 125790 652410 125880 652650
rect 126120 652410 126210 652650
rect 126450 652410 126560 652650
rect 126800 652410 126890 652650
rect 127130 652410 127220 652650
rect 127460 652410 127550 652650
rect 127790 652410 127900 652650
rect 128140 652410 128230 652650
rect 128470 652410 128560 652650
rect 128800 652410 128890 652650
rect 129130 652410 129240 652650
rect 129480 652410 129570 652650
rect 129810 652410 129900 652650
rect 130140 652410 130230 652650
rect 130470 652410 130580 652650
rect 130820 652410 130910 652650
rect 131150 652410 131240 652650
rect 131480 652410 131570 652650
rect 131810 652410 131920 652650
rect 132160 652410 132250 652650
rect 132490 652410 132580 652650
rect 132820 652410 132910 652650
rect 133150 652410 133170 652650
rect 122170 652300 133170 652410
rect 122170 652060 122190 652300
rect 122430 652060 122540 652300
rect 122780 652060 122870 652300
rect 123110 652060 123200 652300
rect 123440 652060 123530 652300
rect 123770 652060 123880 652300
rect 124120 652060 124210 652300
rect 124450 652060 124540 652300
rect 124780 652060 124870 652300
rect 125110 652060 125220 652300
rect 125460 652060 125550 652300
rect 125790 652060 125880 652300
rect 126120 652060 126210 652300
rect 126450 652060 126560 652300
rect 126800 652060 126890 652300
rect 127130 652060 127220 652300
rect 127460 652060 127550 652300
rect 127790 652060 127900 652300
rect 128140 652060 128230 652300
rect 128470 652060 128560 652300
rect 128800 652060 128890 652300
rect 129130 652060 129240 652300
rect 129480 652060 129570 652300
rect 129810 652060 129900 652300
rect 130140 652060 130230 652300
rect 130470 652060 130580 652300
rect 130820 652060 130910 652300
rect 131150 652060 131240 652300
rect 131480 652060 131570 652300
rect 131810 652060 131920 652300
rect 132160 652060 132250 652300
rect 132490 652060 132580 652300
rect 132820 652060 132910 652300
rect 133150 652060 133170 652300
rect 122170 651970 133170 652060
rect 122170 651730 122190 651970
rect 122430 651730 122540 651970
rect 122780 651730 122870 651970
rect 123110 651730 123200 651970
rect 123440 651730 123530 651970
rect 123770 651730 123880 651970
rect 124120 651730 124210 651970
rect 124450 651730 124540 651970
rect 124780 651730 124870 651970
rect 125110 651730 125220 651970
rect 125460 651730 125550 651970
rect 125790 651730 125880 651970
rect 126120 651730 126210 651970
rect 126450 651730 126560 651970
rect 126800 651730 126890 651970
rect 127130 651730 127220 651970
rect 127460 651730 127550 651970
rect 127790 651730 127900 651970
rect 128140 651730 128230 651970
rect 128470 651730 128560 651970
rect 128800 651730 128890 651970
rect 129130 651730 129240 651970
rect 129480 651730 129570 651970
rect 129810 651730 129900 651970
rect 130140 651730 130230 651970
rect 130470 651730 130580 651970
rect 130820 651730 130910 651970
rect 131150 651730 131240 651970
rect 131480 651730 131570 651970
rect 131810 651730 131920 651970
rect 132160 651730 132250 651970
rect 132490 651730 132580 651970
rect 132820 651730 132910 651970
rect 133150 651730 133170 651970
rect 122170 651640 133170 651730
rect 122170 651400 122190 651640
rect 122430 651400 122540 651640
rect 122780 651400 122870 651640
rect 123110 651400 123200 651640
rect 123440 651400 123530 651640
rect 123770 651400 123880 651640
rect 124120 651400 124210 651640
rect 124450 651400 124540 651640
rect 124780 651400 124870 651640
rect 125110 651400 125220 651640
rect 125460 651400 125550 651640
rect 125790 651400 125880 651640
rect 126120 651400 126210 651640
rect 126450 651400 126560 651640
rect 126800 651400 126890 651640
rect 127130 651400 127220 651640
rect 127460 651400 127550 651640
rect 127790 651400 127900 651640
rect 128140 651400 128230 651640
rect 128470 651400 128560 651640
rect 128800 651400 128890 651640
rect 129130 651400 129240 651640
rect 129480 651400 129570 651640
rect 129810 651400 129900 651640
rect 130140 651400 130230 651640
rect 130470 651400 130580 651640
rect 130820 651400 130910 651640
rect 131150 651400 131240 651640
rect 131480 651400 131570 651640
rect 131810 651400 131920 651640
rect 132160 651400 132250 651640
rect 132490 651400 132580 651640
rect 132820 651400 132910 651640
rect 133150 651400 133170 651640
rect 122170 651310 133170 651400
rect 122170 651070 122190 651310
rect 122430 651070 122540 651310
rect 122780 651070 122870 651310
rect 123110 651070 123200 651310
rect 123440 651070 123530 651310
rect 123770 651070 123880 651310
rect 124120 651070 124210 651310
rect 124450 651070 124540 651310
rect 124780 651070 124870 651310
rect 125110 651070 125220 651310
rect 125460 651070 125550 651310
rect 125790 651070 125880 651310
rect 126120 651070 126210 651310
rect 126450 651070 126560 651310
rect 126800 651070 126890 651310
rect 127130 651070 127220 651310
rect 127460 651070 127550 651310
rect 127790 651070 127900 651310
rect 128140 651070 128230 651310
rect 128470 651070 128560 651310
rect 128800 651070 128890 651310
rect 129130 651070 129240 651310
rect 129480 651070 129570 651310
rect 129810 651070 129900 651310
rect 130140 651070 130230 651310
rect 130470 651070 130580 651310
rect 130820 651070 130910 651310
rect 131150 651070 131240 651310
rect 131480 651070 131570 651310
rect 131810 651070 131920 651310
rect 132160 651070 132250 651310
rect 132490 651070 132580 651310
rect 132820 651070 132910 651310
rect 133150 651070 133170 651310
rect 122170 650960 133170 651070
rect 122170 650720 122190 650960
rect 122430 650720 122540 650960
rect 122780 650720 122870 650960
rect 123110 650720 123200 650960
rect 123440 650720 123530 650960
rect 123770 650720 123880 650960
rect 124120 650720 124210 650960
rect 124450 650720 124540 650960
rect 124780 650720 124870 650960
rect 125110 650720 125220 650960
rect 125460 650720 125550 650960
rect 125790 650720 125880 650960
rect 126120 650720 126210 650960
rect 126450 650720 126560 650960
rect 126800 650720 126890 650960
rect 127130 650720 127220 650960
rect 127460 650720 127550 650960
rect 127790 650720 127900 650960
rect 128140 650720 128230 650960
rect 128470 650720 128560 650960
rect 128800 650720 128890 650960
rect 129130 650720 129240 650960
rect 129480 650720 129570 650960
rect 129810 650720 129900 650960
rect 130140 650720 130230 650960
rect 130470 650720 130580 650960
rect 130820 650720 130910 650960
rect 131150 650720 131240 650960
rect 131480 650720 131570 650960
rect 131810 650720 131920 650960
rect 132160 650720 132250 650960
rect 132490 650720 132580 650960
rect 132820 650720 132910 650960
rect 133150 650720 133170 650960
rect 122170 650630 133170 650720
rect 122170 650390 122190 650630
rect 122430 650390 122540 650630
rect 122780 650390 122870 650630
rect 123110 650390 123200 650630
rect 123440 650390 123530 650630
rect 123770 650390 123880 650630
rect 124120 650390 124210 650630
rect 124450 650390 124540 650630
rect 124780 650390 124870 650630
rect 125110 650390 125220 650630
rect 125460 650390 125550 650630
rect 125790 650390 125880 650630
rect 126120 650390 126210 650630
rect 126450 650390 126560 650630
rect 126800 650390 126890 650630
rect 127130 650390 127220 650630
rect 127460 650390 127550 650630
rect 127790 650390 127900 650630
rect 128140 650390 128230 650630
rect 128470 650390 128560 650630
rect 128800 650390 128890 650630
rect 129130 650390 129240 650630
rect 129480 650390 129570 650630
rect 129810 650390 129900 650630
rect 130140 650390 130230 650630
rect 130470 650390 130580 650630
rect 130820 650390 130910 650630
rect 131150 650390 131240 650630
rect 131480 650390 131570 650630
rect 131810 650390 131920 650630
rect 132160 650390 132250 650630
rect 132490 650390 132580 650630
rect 132820 650390 132910 650630
rect 133150 650390 133170 650630
rect 122170 650300 133170 650390
rect 122170 650060 122190 650300
rect 122430 650060 122540 650300
rect 122780 650060 122870 650300
rect 123110 650060 123200 650300
rect 123440 650060 123530 650300
rect 123770 650060 123880 650300
rect 124120 650060 124210 650300
rect 124450 650060 124540 650300
rect 124780 650060 124870 650300
rect 125110 650060 125220 650300
rect 125460 650060 125550 650300
rect 125790 650060 125880 650300
rect 126120 650060 126210 650300
rect 126450 650060 126560 650300
rect 126800 650060 126890 650300
rect 127130 650060 127220 650300
rect 127460 650060 127550 650300
rect 127790 650060 127900 650300
rect 128140 650060 128230 650300
rect 128470 650060 128560 650300
rect 128800 650060 128890 650300
rect 129130 650060 129240 650300
rect 129480 650060 129570 650300
rect 129810 650060 129900 650300
rect 130140 650060 130230 650300
rect 130470 650060 130580 650300
rect 130820 650060 130910 650300
rect 131150 650060 131240 650300
rect 131480 650060 131570 650300
rect 131810 650060 131920 650300
rect 132160 650060 132250 650300
rect 132490 650060 132580 650300
rect 132820 650060 132910 650300
rect 133150 650060 133170 650300
rect 122170 649970 133170 650060
rect 122170 649730 122190 649970
rect 122430 649730 122540 649970
rect 122780 649730 122870 649970
rect 123110 649730 123200 649970
rect 123440 649730 123530 649970
rect 123770 649730 123880 649970
rect 124120 649730 124210 649970
rect 124450 649730 124540 649970
rect 124780 649730 124870 649970
rect 125110 649730 125220 649970
rect 125460 649730 125550 649970
rect 125790 649730 125880 649970
rect 126120 649730 126210 649970
rect 126450 649730 126560 649970
rect 126800 649730 126890 649970
rect 127130 649730 127220 649970
rect 127460 649730 127550 649970
rect 127790 649730 127900 649970
rect 128140 649730 128230 649970
rect 128470 649730 128560 649970
rect 128800 649730 128890 649970
rect 129130 649730 129240 649970
rect 129480 649730 129570 649970
rect 129810 649730 129900 649970
rect 130140 649730 130230 649970
rect 130470 649730 130580 649970
rect 130820 649730 130910 649970
rect 131150 649730 131240 649970
rect 131480 649730 131570 649970
rect 131810 649730 131920 649970
rect 132160 649730 132250 649970
rect 132490 649730 132580 649970
rect 132820 649730 132910 649970
rect 133150 649730 133170 649970
rect 122170 649620 133170 649730
rect 122170 649380 122190 649620
rect 122430 649380 122540 649620
rect 122780 649380 122870 649620
rect 123110 649380 123200 649620
rect 123440 649380 123530 649620
rect 123770 649380 123880 649620
rect 124120 649380 124210 649620
rect 124450 649380 124540 649620
rect 124780 649380 124870 649620
rect 125110 649380 125220 649620
rect 125460 649380 125550 649620
rect 125790 649380 125880 649620
rect 126120 649380 126210 649620
rect 126450 649380 126560 649620
rect 126800 649380 126890 649620
rect 127130 649380 127220 649620
rect 127460 649380 127550 649620
rect 127790 649380 127900 649620
rect 128140 649380 128230 649620
rect 128470 649380 128560 649620
rect 128800 649380 128890 649620
rect 129130 649380 129240 649620
rect 129480 649380 129570 649620
rect 129810 649380 129900 649620
rect 130140 649380 130230 649620
rect 130470 649380 130580 649620
rect 130820 649380 130910 649620
rect 131150 649380 131240 649620
rect 131480 649380 131570 649620
rect 131810 649380 131920 649620
rect 132160 649380 132250 649620
rect 132490 649380 132580 649620
rect 132820 649380 132910 649620
rect 133150 649380 133170 649620
rect 122170 649360 133170 649380
rect 133550 660340 144550 660360
rect 133550 660100 133570 660340
rect 133810 660100 133920 660340
rect 134160 660100 134250 660340
rect 134490 660100 134580 660340
rect 134820 660100 134910 660340
rect 135150 660100 135260 660340
rect 135500 660100 135590 660340
rect 135830 660100 135920 660340
rect 136160 660100 136250 660340
rect 136490 660100 136600 660340
rect 136840 660100 136930 660340
rect 137170 660100 137260 660340
rect 137500 660100 137590 660340
rect 137830 660100 137940 660340
rect 138180 660100 138270 660340
rect 138510 660100 138600 660340
rect 138840 660100 138930 660340
rect 139170 660100 139280 660340
rect 139520 660100 139610 660340
rect 139850 660100 139940 660340
rect 140180 660100 140270 660340
rect 140510 660100 140620 660340
rect 140860 660100 140950 660340
rect 141190 660100 141280 660340
rect 141520 660100 141610 660340
rect 141850 660100 141960 660340
rect 142200 660100 142290 660340
rect 142530 660100 142620 660340
rect 142860 660100 142950 660340
rect 143190 660100 143300 660340
rect 143540 660100 143630 660340
rect 143870 660100 143960 660340
rect 144200 660100 144290 660340
rect 144530 660100 144550 660340
rect 133550 660010 144550 660100
rect 133550 659770 133570 660010
rect 133810 659770 133920 660010
rect 134160 659770 134250 660010
rect 134490 659770 134580 660010
rect 134820 659770 134910 660010
rect 135150 659770 135260 660010
rect 135500 659770 135590 660010
rect 135830 659770 135920 660010
rect 136160 659770 136250 660010
rect 136490 659770 136600 660010
rect 136840 659770 136930 660010
rect 137170 659770 137260 660010
rect 137500 659770 137590 660010
rect 137830 659770 137940 660010
rect 138180 659770 138270 660010
rect 138510 659770 138600 660010
rect 138840 659770 138930 660010
rect 139170 659770 139280 660010
rect 139520 659770 139610 660010
rect 139850 659770 139940 660010
rect 140180 659770 140270 660010
rect 140510 659770 140620 660010
rect 140860 659770 140950 660010
rect 141190 659770 141280 660010
rect 141520 659770 141610 660010
rect 141850 659770 141960 660010
rect 142200 659770 142290 660010
rect 142530 659770 142620 660010
rect 142860 659770 142950 660010
rect 143190 659770 143300 660010
rect 143540 659770 143630 660010
rect 143870 659770 143960 660010
rect 144200 659770 144290 660010
rect 144530 659770 144550 660010
rect 133550 659680 144550 659770
rect 133550 659440 133570 659680
rect 133810 659440 133920 659680
rect 134160 659440 134250 659680
rect 134490 659440 134580 659680
rect 134820 659440 134910 659680
rect 135150 659440 135260 659680
rect 135500 659440 135590 659680
rect 135830 659440 135920 659680
rect 136160 659440 136250 659680
rect 136490 659440 136600 659680
rect 136840 659440 136930 659680
rect 137170 659440 137260 659680
rect 137500 659440 137590 659680
rect 137830 659440 137940 659680
rect 138180 659440 138270 659680
rect 138510 659440 138600 659680
rect 138840 659440 138930 659680
rect 139170 659440 139280 659680
rect 139520 659440 139610 659680
rect 139850 659440 139940 659680
rect 140180 659440 140270 659680
rect 140510 659440 140620 659680
rect 140860 659440 140950 659680
rect 141190 659440 141280 659680
rect 141520 659440 141610 659680
rect 141850 659440 141960 659680
rect 142200 659440 142290 659680
rect 142530 659440 142620 659680
rect 142860 659440 142950 659680
rect 143190 659440 143300 659680
rect 143540 659440 143630 659680
rect 143870 659440 143960 659680
rect 144200 659440 144290 659680
rect 144530 659440 144550 659680
rect 133550 659350 144550 659440
rect 133550 659110 133570 659350
rect 133810 659110 133920 659350
rect 134160 659110 134250 659350
rect 134490 659110 134580 659350
rect 134820 659110 134910 659350
rect 135150 659110 135260 659350
rect 135500 659110 135590 659350
rect 135830 659110 135920 659350
rect 136160 659110 136250 659350
rect 136490 659110 136600 659350
rect 136840 659110 136930 659350
rect 137170 659110 137260 659350
rect 137500 659110 137590 659350
rect 137830 659110 137940 659350
rect 138180 659110 138270 659350
rect 138510 659110 138600 659350
rect 138840 659110 138930 659350
rect 139170 659110 139280 659350
rect 139520 659110 139610 659350
rect 139850 659110 139940 659350
rect 140180 659110 140270 659350
rect 140510 659110 140620 659350
rect 140860 659110 140950 659350
rect 141190 659110 141280 659350
rect 141520 659110 141610 659350
rect 141850 659110 141960 659350
rect 142200 659110 142290 659350
rect 142530 659110 142620 659350
rect 142860 659110 142950 659350
rect 143190 659110 143300 659350
rect 143540 659110 143630 659350
rect 143870 659110 143960 659350
rect 144200 659110 144290 659350
rect 144530 659110 144550 659350
rect 133550 659000 144550 659110
rect 133550 658760 133570 659000
rect 133810 658760 133920 659000
rect 134160 658760 134250 659000
rect 134490 658760 134580 659000
rect 134820 658760 134910 659000
rect 135150 658760 135260 659000
rect 135500 658760 135590 659000
rect 135830 658760 135920 659000
rect 136160 658760 136250 659000
rect 136490 658760 136600 659000
rect 136840 658760 136930 659000
rect 137170 658760 137260 659000
rect 137500 658760 137590 659000
rect 137830 658760 137940 659000
rect 138180 658760 138270 659000
rect 138510 658760 138600 659000
rect 138840 658760 138930 659000
rect 139170 658760 139280 659000
rect 139520 658760 139610 659000
rect 139850 658760 139940 659000
rect 140180 658760 140270 659000
rect 140510 658760 140620 659000
rect 140860 658760 140950 659000
rect 141190 658760 141280 659000
rect 141520 658760 141610 659000
rect 141850 658760 141960 659000
rect 142200 658760 142290 659000
rect 142530 658760 142620 659000
rect 142860 658760 142950 659000
rect 143190 658760 143300 659000
rect 143540 658760 143630 659000
rect 143870 658760 143960 659000
rect 144200 658760 144290 659000
rect 144530 658760 144550 659000
rect 133550 658670 144550 658760
rect 133550 658430 133570 658670
rect 133810 658430 133920 658670
rect 134160 658430 134250 658670
rect 134490 658430 134580 658670
rect 134820 658430 134910 658670
rect 135150 658430 135260 658670
rect 135500 658430 135590 658670
rect 135830 658430 135920 658670
rect 136160 658430 136250 658670
rect 136490 658430 136600 658670
rect 136840 658430 136930 658670
rect 137170 658430 137260 658670
rect 137500 658430 137590 658670
rect 137830 658430 137940 658670
rect 138180 658430 138270 658670
rect 138510 658430 138600 658670
rect 138840 658430 138930 658670
rect 139170 658430 139280 658670
rect 139520 658430 139610 658670
rect 139850 658430 139940 658670
rect 140180 658430 140270 658670
rect 140510 658430 140620 658670
rect 140860 658430 140950 658670
rect 141190 658430 141280 658670
rect 141520 658430 141610 658670
rect 141850 658430 141960 658670
rect 142200 658430 142290 658670
rect 142530 658430 142620 658670
rect 142860 658430 142950 658670
rect 143190 658430 143300 658670
rect 143540 658430 143630 658670
rect 143870 658430 143960 658670
rect 144200 658430 144290 658670
rect 144530 658430 144550 658670
rect 133550 658340 144550 658430
rect 133550 658100 133570 658340
rect 133810 658100 133920 658340
rect 134160 658100 134250 658340
rect 134490 658100 134580 658340
rect 134820 658100 134910 658340
rect 135150 658100 135260 658340
rect 135500 658100 135590 658340
rect 135830 658100 135920 658340
rect 136160 658100 136250 658340
rect 136490 658100 136600 658340
rect 136840 658100 136930 658340
rect 137170 658100 137260 658340
rect 137500 658100 137590 658340
rect 137830 658100 137940 658340
rect 138180 658100 138270 658340
rect 138510 658100 138600 658340
rect 138840 658100 138930 658340
rect 139170 658100 139280 658340
rect 139520 658100 139610 658340
rect 139850 658100 139940 658340
rect 140180 658100 140270 658340
rect 140510 658100 140620 658340
rect 140860 658100 140950 658340
rect 141190 658100 141280 658340
rect 141520 658100 141610 658340
rect 141850 658100 141960 658340
rect 142200 658100 142290 658340
rect 142530 658100 142620 658340
rect 142860 658100 142950 658340
rect 143190 658100 143300 658340
rect 143540 658100 143630 658340
rect 143870 658100 143960 658340
rect 144200 658100 144290 658340
rect 144530 658100 144550 658340
rect 133550 658010 144550 658100
rect 133550 657770 133570 658010
rect 133810 657770 133920 658010
rect 134160 657770 134250 658010
rect 134490 657770 134580 658010
rect 134820 657770 134910 658010
rect 135150 657770 135260 658010
rect 135500 657770 135590 658010
rect 135830 657770 135920 658010
rect 136160 657770 136250 658010
rect 136490 657770 136600 658010
rect 136840 657770 136930 658010
rect 137170 657770 137260 658010
rect 137500 657770 137590 658010
rect 137830 657770 137940 658010
rect 138180 657770 138270 658010
rect 138510 657770 138600 658010
rect 138840 657770 138930 658010
rect 139170 657770 139280 658010
rect 139520 657770 139610 658010
rect 139850 657770 139940 658010
rect 140180 657770 140270 658010
rect 140510 657770 140620 658010
rect 140860 657770 140950 658010
rect 141190 657770 141280 658010
rect 141520 657770 141610 658010
rect 141850 657770 141960 658010
rect 142200 657770 142290 658010
rect 142530 657770 142620 658010
rect 142860 657770 142950 658010
rect 143190 657770 143300 658010
rect 143540 657770 143630 658010
rect 143870 657770 143960 658010
rect 144200 657770 144290 658010
rect 144530 657770 144550 658010
rect 133550 657660 144550 657770
rect 133550 657420 133570 657660
rect 133810 657420 133920 657660
rect 134160 657420 134250 657660
rect 134490 657420 134580 657660
rect 134820 657420 134910 657660
rect 135150 657420 135260 657660
rect 135500 657420 135590 657660
rect 135830 657420 135920 657660
rect 136160 657420 136250 657660
rect 136490 657420 136600 657660
rect 136840 657420 136930 657660
rect 137170 657420 137260 657660
rect 137500 657420 137590 657660
rect 137830 657420 137940 657660
rect 138180 657420 138270 657660
rect 138510 657420 138600 657660
rect 138840 657420 138930 657660
rect 139170 657420 139280 657660
rect 139520 657420 139610 657660
rect 139850 657420 139940 657660
rect 140180 657420 140270 657660
rect 140510 657420 140620 657660
rect 140860 657420 140950 657660
rect 141190 657420 141280 657660
rect 141520 657420 141610 657660
rect 141850 657420 141960 657660
rect 142200 657420 142290 657660
rect 142530 657420 142620 657660
rect 142860 657420 142950 657660
rect 143190 657420 143300 657660
rect 143540 657420 143630 657660
rect 143870 657420 143960 657660
rect 144200 657420 144290 657660
rect 144530 657420 144550 657660
rect 133550 657330 144550 657420
rect 133550 657090 133570 657330
rect 133810 657090 133920 657330
rect 134160 657090 134250 657330
rect 134490 657090 134580 657330
rect 134820 657090 134910 657330
rect 135150 657090 135260 657330
rect 135500 657090 135590 657330
rect 135830 657090 135920 657330
rect 136160 657090 136250 657330
rect 136490 657090 136600 657330
rect 136840 657090 136930 657330
rect 137170 657090 137260 657330
rect 137500 657090 137590 657330
rect 137830 657090 137940 657330
rect 138180 657090 138270 657330
rect 138510 657090 138600 657330
rect 138840 657090 138930 657330
rect 139170 657090 139280 657330
rect 139520 657090 139610 657330
rect 139850 657090 139940 657330
rect 140180 657090 140270 657330
rect 140510 657090 140620 657330
rect 140860 657090 140950 657330
rect 141190 657090 141280 657330
rect 141520 657090 141610 657330
rect 141850 657090 141960 657330
rect 142200 657090 142290 657330
rect 142530 657090 142620 657330
rect 142860 657090 142950 657330
rect 143190 657090 143300 657330
rect 143540 657090 143630 657330
rect 143870 657090 143960 657330
rect 144200 657090 144290 657330
rect 144530 657090 144550 657330
rect 133550 657000 144550 657090
rect 133550 656760 133570 657000
rect 133810 656760 133920 657000
rect 134160 656760 134250 657000
rect 134490 656760 134580 657000
rect 134820 656760 134910 657000
rect 135150 656760 135260 657000
rect 135500 656760 135590 657000
rect 135830 656760 135920 657000
rect 136160 656760 136250 657000
rect 136490 656760 136600 657000
rect 136840 656760 136930 657000
rect 137170 656760 137260 657000
rect 137500 656760 137590 657000
rect 137830 656760 137940 657000
rect 138180 656760 138270 657000
rect 138510 656760 138600 657000
rect 138840 656760 138930 657000
rect 139170 656760 139280 657000
rect 139520 656760 139610 657000
rect 139850 656760 139940 657000
rect 140180 656760 140270 657000
rect 140510 656760 140620 657000
rect 140860 656760 140950 657000
rect 141190 656760 141280 657000
rect 141520 656760 141610 657000
rect 141850 656760 141960 657000
rect 142200 656760 142290 657000
rect 142530 656760 142620 657000
rect 142860 656760 142950 657000
rect 143190 656760 143300 657000
rect 143540 656760 143630 657000
rect 143870 656760 143960 657000
rect 144200 656760 144290 657000
rect 144530 656760 144550 657000
rect 133550 656670 144550 656760
rect 133550 656430 133570 656670
rect 133810 656430 133920 656670
rect 134160 656430 134250 656670
rect 134490 656430 134580 656670
rect 134820 656430 134910 656670
rect 135150 656430 135260 656670
rect 135500 656430 135590 656670
rect 135830 656430 135920 656670
rect 136160 656430 136250 656670
rect 136490 656430 136600 656670
rect 136840 656430 136930 656670
rect 137170 656430 137260 656670
rect 137500 656430 137590 656670
rect 137830 656430 137940 656670
rect 138180 656430 138270 656670
rect 138510 656430 138600 656670
rect 138840 656430 138930 656670
rect 139170 656430 139280 656670
rect 139520 656430 139610 656670
rect 139850 656430 139940 656670
rect 140180 656430 140270 656670
rect 140510 656430 140620 656670
rect 140860 656430 140950 656670
rect 141190 656430 141280 656670
rect 141520 656430 141610 656670
rect 141850 656430 141960 656670
rect 142200 656430 142290 656670
rect 142530 656430 142620 656670
rect 142860 656430 142950 656670
rect 143190 656430 143300 656670
rect 143540 656430 143630 656670
rect 143870 656430 143960 656670
rect 144200 656430 144290 656670
rect 144530 656430 144550 656670
rect 133550 656320 144550 656430
rect 133550 656080 133570 656320
rect 133810 656080 133920 656320
rect 134160 656080 134250 656320
rect 134490 656080 134580 656320
rect 134820 656080 134910 656320
rect 135150 656080 135260 656320
rect 135500 656080 135590 656320
rect 135830 656080 135920 656320
rect 136160 656080 136250 656320
rect 136490 656080 136600 656320
rect 136840 656080 136930 656320
rect 137170 656080 137260 656320
rect 137500 656080 137590 656320
rect 137830 656080 137940 656320
rect 138180 656080 138270 656320
rect 138510 656080 138600 656320
rect 138840 656080 138930 656320
rect 139170 656080 139280 656320
rect 139520 656080 139610 656320
rect 139850 656080 139940 656320
rect 140180 656080 140270 656320
rect 140510 656080 140620 656320
rect 140860 656080 140950 656320
rect 141190 656080 141280 656320
rect 141520 656080 141610 656320
rect 141850 656080 141960 656320
rect 142200 656080 142290 656320
rect 142530 656080 142620 656320
rect 142860 656080 142950 656320
rect 143190 656080 143300 656320
rect 143540 656080 143630 656320
rect 143870 656080 143960 656320
rect 144200 656080 144290 656320
rect 144530 656080 144550 656320
rect 133550 655990 144550 656080
rect 133550 655750 133570 655990
rect 133810 655750 133920 655990
rect 134160 655750 134250 655990
rect 134490 655750 134580 655990
rect 134820 655750 134910 655990
rect 135150 655750 135260 655990
rect 135500 655750 135590 655990
rect 135830 655750 135920 655990
rect 136160 655750 136250 655990
rect 136490 655750 136600 655990
rect 136840 655750 136930 655990
rect 137170 655750 137260 655990
rect 137500 655750 137590 655990
rect 137830 655750 137940 655990
rect 138180 655750 138270 655990
rect 138510 655750 138600 655990
rect 138840 655750 138930 655990
rect 139170 655750 139280 655990
rect 139520 655750 139610 655990
rect 139850 655750 139940 655990
rect 140180 655750 140270 655990
rect 140510 655750 140620 655990
rect 140860 655750 140950 655990
rect 141190 655750 141280 655990
rect 141520 655750 141610 655990
rect 141850 655750 141960 655990
rect 142200 655750 142290 655990
rect 142530 655750 142620 655990
rect 142860 655750 142950 655990
rect 143190 655750 143300 655990
rect 143540 655750 143630 655990
rect 143870 655750 143960 655990
rect 144200 655750 144290 655990
rect 144530 655750 144550 655990
rect 133550 655660 144550 655750
rect 133550 655420 133570 655660
rect 133810 655420 133920 655660
rect 134160 655420 134250 655660
rect 134490 655420 134580 655660
rect 134820 655420 134910 655660
rect 135150 655420 135260 655660
rect 135500 655420 135590 655660
rect 135830 655420 135920 655660
rect 136160 655420 136250 655660
rect 136490 655420 136600 655660
rect 136840 655420 136930 655660
rect 137170 655420 137260 655660
rect 137500 655420 137590 655660
rect 137830 655420 137940 655660
rect 138180 655420 138270 655660
rect 138510 655420 138600 655660
rect 138840 655420 138930 655660
rect 139170 655420 139280 655660
rect 139520 655420 139610 655660
rect 139850 655420 139940 655660
rect 140180 655420 140270 655660
rect 140510 655420 140620 655660
rect 140860 655420 140950 655660
rect 141190 655420 141280 655660
rect 141520 655420 141610 655660
rect 141850 655420 141960 655660
rect 142200 655420 142290 655660
rect 142530 655420 142620 655660
rect 142860 655420 142950 655660
rect 143190 655420 143300 655660
rect 143540 655420 143630 655660
rect 143870 655420 143960 655660
rect 144200 655420 144290 655660
rect 144530 655420 144550 655660
rect 133550 655330 144550 655420
rect 133550 655090 133570 655330
rect 133810 655090 133920 655330
rect 134160 655090 134250 655330
rect 134490 655090 134580 655330
rect 134820 655090 134910 655330
rect 135150 655090 135260 655330
rect 135500 655090 135590 655330
rect 135830 655090 135920 655330
rect 136160 655090 136250 655330
rect 136490 655090 136600 655330
rect 136840 655090 136930 655330
rect 137170 655090 137260 655330
rect 137500 655090 137590 655330
rect 137830 655090 137940 655330
rect 138180 655090 138270 655330
rect 138510 655090 138600 655330
rect 138840 655090 138930 655330
rect 139170 655090 139280 655330
rect 139520 655090 139610 655330
rect 139850 655090 139940 655330
rect 140180 655090 140270 655330
rect 140510 655090 140620 655330
rect 140860 655090 140950 655330
rect 141190 655090 141280 655330
rect 141520 655090 141610 655330
rect 141850 655090 141960 655330
rect 142200 655090 142290 655330
rect 142530 655090 142620 655330
rect 142860 655090 142950 655330
rect 143190 655090 143300 655330
rect 143540 655090 143630 655330
rect 143870 655090 143960 655330
rect 144200 655090 144290 655330
rect 144530 655090 144550 655330
rect 133550 654980 144550 655090
rect 133550 654740 133570 654980
rect 133810 654740 133920 654980
rect 134160 654740 134250 654980
rect 134490 654740 134580 654980
rect 134820 654740 134910 654980
rect 135150 654740 135260 654980
rect 135500 654740 135590 654980
rect 135830 654740 135920 654980
rect 136160 654740 136250 654980
rect 136490 654740 136600 654980
rect 136840 654740 136930 654980
rect 137170 654740 137260 654980
rect 137500 654740 137590 654980
rect 137830 654740 137940 654980
rect 138180 654740 138270 654980
rect 138510 654740 138600 654980
rect 138840 654740 138930 654980
rect 139170 654740 139280 654980
rect 139520 654740 139610 654980
rect 139850 654740 139940 654980
rect 140180 654740 140270 654980
rect 140510 654740 140620 654980
rect 140860 654740 140950 654980
rect 141190 654740 141280 654980
rect 141520 654740 141610 654980
rect 141850 654740 141960 654980
rect 142200 654740 142290 654980
rect 142530 654740 142620 654980
rect 142860 654740 142950 654980
rect 143190 654740 143300 654980
rect 143540 654740 143630 654980
rect 143870 654740 143960 654980
rect 144200 654740 144290 654980
rect 144530 654740 144550 654980
rect 133550 654650 144550 654740
rect 133550 654410 133570 654650
rect 133810 654410 133920 654650
rect 134160 654410 134250 654650
rect 134490 654410 134580 654650
rect 134820 654410 134910 654650
rect 135150 654410 135260 654650
rect 135500 654410 135590 654650
rect 135830 654410 135920 654650
rect 136160 654410 136250 654650
rect 136490 654410 136600 654650
rect 136840 654410 136930 654650
rect 137170 654410 137260 654650
rect 137500 654410 137590 654650
rect 137830 654410 137940 654650
rect 138180 654410 138270 654650
rect 138510 654410 138600 654650
rect 138840 654410 138930 654650
rect 139170 654410 139280 654650
rect 139520 654410 139610 654650
rect 139850 654410 139940 654650
rect 140180 654410 140270 654650
rect 140510 654410 140620 654650
rect 140860 654410 140950 654650
rect 141190 654410 141280 654650
rect 141520 654410 141610 654650
rect 141850 654410 141960 654650
rect 142200 654410 142290 654650
rect 142530 654410 142620 654650
rect 142860 654410 142950 654650
rect 143190 654410 143300 654650
rect 143540 654410 143630 654650
rect 143870 654410 143960 654650
rect 144200 654410 144290 654650
rect 144530 654410 144550 654650
rect 133550 654320 144550 654410
rect 133550 654080 133570 654320
rect 133810 654080 133920 654320
rect 134160 654080 134250 654320
rect 134490 654080 134580 654320
rect 134820 654080 134910 654320
rect 135150 654080 135260 654320
rect 135500 654080 135590 654320
rect 135830 654080 135920 654320
rect 136160 654080 136250 654320
rect 136490 654080 136600 654320
rect 136840 654080 136930 654320
rect 137170 654080 137260 654320
rect 137500 654080 137590 654320
rect 137830 654080 137940 654320
rect 138180 654080 138270 654320
rect 138510 654080 138600 654320
rect 138840 654080 138930 654320
rect 139170 654080 139280 654320
rect 139520 654080 139610 654320
rect 139850 654080 139940 654320
rect 140180 654080 140270 654320
rect 140510 654080 140620 654320
rect 140860 654080 140950 654320
rect 141190 654080 141280 654320
rect 141520 654080 141610 654320
rect 141850 654080 141960 654320
rect 142200 654080 142290 654320
rect 142530 654080 142620 654320
rect 142860 654080 142950 654320
rect 143190 654080 143300 654320
rect 143540 654080 143630 654320
rect 143870 654080 143960 654320
rect 144200 654080 144290 654320
rect 144530 654080 144550 654320
rect 133550 653990 144550 654080
rect 133550 653750 133570 653990
rect 133810 653750 133920 653990
rect 134160 653750 134250 653990
rect 134490 653750 134580 653990
rect 134820 653750 134910 653990
rect 135150 653750 135260 653990
rect 135500 653750 135590 653990
rect 135830 653750 135920 653990
rect 136160 653750 136250 653990
rect 136490 653750 136600 653990
rect 136840 653750 136930 653990
rect 137170 653750 137260 653990
rect 137500 653750 137590 653990
rect 137830 653750 137940 653990
rect 138180 653750 138270 653990
rect 138510 653750 138600 653990
rect 138840 653750 138930 653990
rect 139170 653750 139280 653990
rect 139520 653750 139610 653990
rect 139850 653750 139940 653990
rect 140180 653750 140270 653990
rect 140510 653750 140620 653990
rect 140860 653750 140950 653990
rect 141190 653750 141280 653990
rect 141520 653750 141610 653990
rect 141850 653750 141960 653990
rect 142200 653750 142290 653990
rect 142530 653750 142620 653990
rect 142860 653750 142950 653990
rect 143190 653750 143300 653990
rect 143540 653750 143630 653990
rect 143870 653750 143960 653990
rect 144200 653750 144290 653990
rect 144530 653750 144550 653990
rect 133550 653640 144550 653750
rect 133550 653400 133570 653640
rect 133810 653400 133920 653640
rect 134160 653400 134250 653640
rect 134490 653400 134580 653640
rect 134820 653400 134910 653640
rect 135150 653400 135260 653640
rect 135500 653400 135590 653640
rect 135830 653400 135920 653640
rect 136160 653400 136250 653640
rect 136490 653400 136600 653640
rect 136840 653400 136930 653640
rect 137170 653400 137260 653640
rect 137500 653400 137590 653640
rect 137830 653400 137940 653640
rect 138180 653400 138270 653640
rect 138510 653400 138600 653640
rect 138840 653400 138930 653640
rect 139170 653400 139280 653640
rect 139520 653400 139610 653640
rect 139850 653400 139940 653640
rect 140180 653400 140270 653640
rect 140510 653400 140620 653640
rect 140860 653400 140950 653640
rect 141190 653400 141280 653640
rect 141520 653400 141610 653640
rect 141850 653400 141960 653640
rect 142200 653400 142290 653640
rect 142530 653400 142620 653640
rect 142860 653400 142950 653640
rect 143190 653400 143300 653640
rect 143540 653400 143630 653640
rect 143870 653400 143960 653640
rect 144200 653400 144290 653640
rect 144530 653400 144550 653640
rect 133550 653310 144550 653400
rect 133550 653070 133570 653310
rect 133810 653070 133920 653310
rect 134160 653070 134250 653310
rect 134490 653070 134580 653310
rect 134820 653070 134910 653310
rect 135150 653070 135260 653310
rect 135500 653070 135590 653310
rect 135830 653070 135920 653310
rect 136160 653070 136250 653310
rect 136490 653070 136600 653310
rect 136840 653070 136930 653310
rect 137170 653070 137260 653310
rect 137500 653070 137590 653310
rect 137830 653070 137940 653310
rect 138180 653070 138270 653310
rect 138510 653070 138600 653310
rect 138840 653070 138930 653310
rect 139170 653070 139280 653310
rect 139520 653070 139610 653310
rect 139850 653070 139940 653310
rect 140180 653070 140270 653310
rect 140510 653070 140620 653310
rect 140860 653070 140950 653310
rect 141190 653070 141280 653310
rect 141520 653070 141610 653310
rect 141850 653070 141960 653310
rect 142200 653070 142290 653310
rect 142530 653070 142620 653310
rect 142860 653070 142950 653310
rect 143190 653070 143300 653310
rect 143540 653070 143630 653310
rect 143870 653070 143960 653310
rect 144200 653070 144290 653310
rect 144530 653070 144550 653310
rect 133550 652980 144550 653070
rect 133550 652740 133570 652980
rect 133810 652740 133920 652980
rect 134160 652740 134250 652980
rect 134490 652740 134580 652980
rect 134820 652740 134910 652980
rect 135150 652740 135260 652980
rect 135500 652740 135590 652980
rect 135830 652740 135920 652980
rect 136160 652740 136250 652980
rect 136490 652740 136600 652980
rect 136840 652740 136930 652980
rect 137170 652740 137260 652980
rect 137500 652740 137590 652980
rect 137830 652740 137940 652980
rect 138180 652740 138270 652980
rect 138510 652740 138600 652980
rect 138840 652740 138930 652980
rect 139170 652740 139280 652980
rect 139520 652740 139610 652980
rect 139850 652740 139940 652980
rect 140180 652740 140270 652980
rect 140510 652740 140620 652980
rect 140860 652740 140950 652980
rect 141190 652740 141280 652980
rect 141520 652740 141610 652980
rect 141850 652740 141960 652980
rect 142200 652740 142290 652980
rect 142530 652740 142620 652980
rect 142860 652740 142950 652980
rect 143190 652740 143300 652980
rect 143540 652740 143630 652980
rect 143870 652740 143960 652980
rect 144200 652740 144290 652980
rect 144530 652740 144550 652980
rect 133550 652650 144550 652740
rect 133550 652410 133570 652650
rect 133810 652410 133920 652650
rect 134160 652410 134250 652650
rect 134490 652410 134580 652650
rect 134820 652410 134910 652650
rect 135150 652410 135260 652650
rect 135500 652410 135590 652650
rect 135830 652410 135920 652650
rect 136160 652410 136250 652650
rect 136490 652410 136600 652650
rect 136840 652410 136930 652650
rect 137170 652410 137260 652650
rect 137500 652410 137590 652650
rect 137830 652410 137940 652650
rect 138180 652410 138270 652650
rect 138510 652410 138600 652650
rect 138840 652410 138930 652650
rect 139170 652410 139280 652650
rect 139520 652410 139610 652650
rect 139850 652410 139940 652650
rect 140180 652410 140270 652650
rect 140510 652410 140620 652650
rect 140860 652410 140950 652650
rect 141190 652410 141280 652650
rect 141520 652410 141610 652650
rect 141850 652410 141960 652650
rect 142200 652410 142290 652650
rect 142530 652410 142620 652650
rect 142860 652410 142950 652650
rect 143190 652410 143300 652650
rect 143540 652410 143630 652650
rect 143870 652410 143960 652650
rect 144200 652410 144290 652650
rect 144530 652410 144550 652650
rect 133550 652300 144550 652410
rect 133550 652060 133570 652300
rect 133810 652060 133920 652300
rect 134160 652060 134250 652300
rect 134490 652060 134580 652300
rect 134820 652060 134910 652300
rect 135150 652060 135260 652300
rect 135500 652060 135590 652300
rect 135830 652060 135920 652300
rect 136160 652060 136250 652300
rect 136490 652060 136600 652300
rect 136840 652060 136930 652300
rect 137170 652060 137260 652300
rect 137500 652060 137590 652300
rect 137830 652060 137940 652300
rect 138180 652060 138270 652300
rect 138510 652060 138600 652300
rect 138840 652060 138930 652300
rect 139170 652060 139280 652300
rect 139520 652060 139610 652300
rect 139850 652060 139940 652300
rect 140180 652060 140270 652300
rect 140510 652060 140620 652300
rect 140860 652060 140950 652300
rect 141190 652060 141280 652300
rect 141520 652060 141610 652300
rect 141850 652060 141960 652300
rect 142200 652060 142290 652300
rect 142530 652060 142620 652300
rect 142860 652060 142950 652300
rect 143190 652060 143300 652300
rect 143540 652060 143630 652300
rect 143870 652060 143960 652300
rect 144200 652060 144290 652300
rect 144530 652060 144550 652300
rect 133550 651970 144550 652060
rect 133550 651730 133570 651970
rect 133810 651730 133920 651970
rect 134160 651730 134250 651970
rect 134490 651730 134580 651970
rect 134820 651730 134910 651970
rect 135150 651730 135260 651970
rect 135500 651730 135590 651970
rect 135830 651730 135920 651970
rect 136160 651730 136250 651970
rect 136490 651730 136600 651970
rect 136840 651730 136930 651970
rect 137170 651730 137260 651970
rect 137500 651730 137590 651970
rect 137830 651730 137940 651970
rect 138180 651730 138270 651970
rect 138510 651730 138600 651970
rect 138840 651730 138930 651970
rect 139170 651730 139280 651970
rect 139520 651730 139610 651970
rect 139850 651730 139940 651970
rect 140180 651730 140270 651970
rect 140510 651730 140620 651970
rect 140860 651730 140950 651970
rect 141190 651730 141280 651970
rect 141520 651730 141610 651970
rect 141850 651730 141960 651970
rect 142200 651730 142290 651970
rect 142530 651730 142620 651970
rect 142860 651730 142950 651970
rect 143190 651730 143300 651970
rect 143540 651730 143630 651970
rect 143870 651730 143960 651970
rect 144200 651730 144290 651970
rect 144530 651730 144550 651970
rect 133550 651640 144550 651730
rect 133550 651400 133570 651640
rect 133810 651400 133920 651640
rect 134160 651400 134250 651640
rect 134490 651400 134580 651640
rect 134820 651400 134910 651640
rect 135150 651400 135260 651640
rect 135500 651400 135590 651640
rect 135830 651400 135920 651640
rect 136160 651400 136250 651640
rect 136490 651400 136600 651640
rect 136840 651400 136930 651640
rect 137170 651400 137260 651640
rect 137500 651400 137590 651640
rect 137830 651400 137940 651640
rect 138180 651400 138270 651640
rect 138510 651400 138600 651640
rect 138840 651400 138930 651640
rect 139170 651400 139280 651640
rect 139520 651400 139610 651640
rect 139850 651400 139940 651640
rect 140180 651400 140270 651640
rect 140510 651400 140620 651640
rect 140860 651400 140950 651640
rect 141190 651400 141280 651640
rect 141520 651400 141610 651640
rect 141850 651400 141960 651640
rect 142200 651400 142290 651640
rect 142530 651400 142620 651640
rect 142860 651400 142950 651640
rect 143190 651400 143300 651640
rect 143540 651400 143630 651640
rect 143870 651400 143960 651640
rect 144200 651400 144290 651640
rect 144530 651400 144550 651640
rect 133550 651310 144550 651400
rect 133550 651070 133570 651310
rect 133810 651070 133920 651310
rect 134160 651070 134250 651310
rect 134490 651070 134580 651310
rect 134820 651070 134910 651310
rect 135150 651070 135260 651310
rect 135500 651070 135590 651310
rect 135830 651070 135920 651310
rect 136160 651070 136250 651310
rect 136490 651070 136600 651310
rect 136840 651070 136930 651310
rect 137170 651070 137260 651310
rect 137500 651070 137590 651310
rect 137830 651070 137940 651310
rect 138180 651070 138270 651310
rect 138510 651070 138600 651310
rect 138840 651070 138930 651310
rect 139170 651070 139280 651310
rect 139520 651070 139610 651310
rect 139850 651070 139940 651310
rect 140180 651070 140270 651310
rect 140510 651070 140620 651310
rect 140860 651070 140950 651310
rect 141190 651070 141280 651310
rect 141520 651070 141610 651310
rect 141850 651070 141960 651310
rect 142200 651070 142290 651310
rect 142530 651070 142620 651310
rect 142860 651070 142950 651310
rect 143190 651070 143300 651310
rect 143540 651070 143630 651310
rect 143870 651070 143960 651310
rect 144200 651070 144290 651310
rect 144530 651070 144550 651310
rect 133550 650960 144550 651070
rect 133550 650720 133570 650960
rect 133810 650720 133920 650960
rect 134160 650720 134250 650960
rect 134490 650720 134580 650960
rect 134820 650720 134910 650960
rect 135150 650720 135260 650960
rect 135500 650720 135590 650960
rect 135830 650720 135920 650960
rect 136160 650720 136250 650960
rect 136490 650720 136600 650960
rect 136840 650720 136930 650960
rect 137170 650720 137260 650960
rect 137500 650720 137590 650960
rect 137830 650720 137940 650960
rect 138180 650720 138270 650960
rect 138510 650720 138600 650960
rect 138840 650720 138930 650960
rect 139170 650720 139280 650960
rect 139520 650720 139610 650960
rect 139850 650720 139940 650960
rect 140180 650720 140270 650960
rect 140510 650720 140620 650960
rect 140860 650720 140950 650960
rect 141190 650720 141280 650960
rect 141520 650720 141610 650960
rect 141850 650720 141960 650960
rect 142200 650720 142290 650960
rect 142530 650720 142620 650960
rect 142860 650720 142950 650960
rect 143190 650720 143300 650960
rect 143540 650720 143630 650960
rect 143870 650720 143960 650960
rect 144200 650720 144290 650960
rect 144530 650720 144550 650960
rect 133550 650630 144550 650720
rect 133550 650390 133570 650630
rect 133810 650390 133920 650630
rect 134160 650390 134250 650630
rect 134490 650390 134580 650630
rect 134820 650390 134910 650630
rect 135150 650390 135260 650630
rect 135500 650390 135590 650630
rect 135830 650390 135920 650630
rect 136160 650390 136250 650630
rect 136490 650390 136600 650630
rect 136840 650390 136930 650630
rect 137170 650390 137260 650630
rect 137500 650390 137590 650630
rect 137830 650390 137940 650630
rect 138180 650390 138270 650630
rect 138510 650390 138600 650630
rect 138840 650390 138930 650630
rect 139170 650390 139280 650630
rect 139520 650390 139610 650630
rect 139850 650390 139940 650630
rect 140180 650390 140270 650630
rect 140510 650390 140620 650630
rect 140860 650390 140950 650630
rect 141190 650390 141280 650630
rect 141520 650390 141610 650630
rect 141850 650390 141960 650630
rect 142200 650390 142290 650630
rect 142530 650390 142620 650630
rect 142860 650390 142950 650630
rect 143190 650390 143300 650630
rect 143540 650390 143630 650630
rect 143870 650390 143960 650630
rect 144200 650390 144290 650630
rect 144530 650390 144550 650630
rect 133550 650300 144550 650390
rect 133550 650060 133570 650300
rect 133810 650060 133920 650300
rect 134160 650060 134250 650300
rect 134490 650060 134580 650300
rect 134820 650060 134910 650300
rect 135150 650060 135260 650300
rect 135500 650060 135590 650300
rect 135830 650060 135920 650300
rect 136160 650060 136250 650300
rect 136490 650060 136600 650300
rect 136840 650060 136930 650300
rect 137170 650060 137260 650300
rect 137500 650060 137590 650300
rect 137830 650060 137940 650300
rect 138180 650060 138270 650300
rect 138510 650060 138600 650300
rect 138840 650060 138930 650300
rect 139170 650060 139280 650300
rect 139520 650060 139610 650300
rect 139850 650060 139940 650300
rect 140180 650060 140270 650300
rect 140510 650060 140620 650300
rect 140860 650060 140950 650300
rect 141190 650060 141280 650300
rect 141520 650060 141610 650300
rect 141850 650060 141960 650300
rect 142200 650060 142290 650300
rect 142530 650060 142620 650300
rect 142860 650060 142950 650300
rect 143190 650060 143300 650300
rect 143540 650060 143630 650300
rect 143870 650060 143960 650300
rect 144200 650060 144290 650300
rect 144530 650060 144550 650300
rect 133550 649970 144550 650060
rect 133550 649730 133570 649970
rect 133810 649730 133920 649970
rect 134160 649730 134250 649970
rect 134490 649730 134580 649970
rect 134820 649730 134910 649970
rect 135150 649730 135260 649970
rect 135500 649730 135590 649970
rect 135830 649730 135920 649970
rect 136160 649730 136250 649970
rect 136490 649730 136600 649970
rect 136840 649730 136930 649970
rect 137170 649730 137260 649970
rect 137500 649730 137590 649970
rect 137830 649730 137940 649970
rect 138180 649730 138270 649970
rect 138510 649730 138600 649970
rect 138840 649730 138930 649970
rect 139170 649730 139280 649970
rect 139520 649730 139610 649970
rect 139850 649730 139940 649970
rect 140180 649730 140270 649970
rect 140510 649730 140620 649970
rect 140860 649730 140950 649970
rect 141190 649730 141280 649970
rect 141520 649730 141610 649970
rect 141850 649730 141960 649970
rect 142200 649730 142290 649970
rect 142530 649730 142620 649970
rect 142860 649730 142950 649970
rect 143190 649730 143300 649970
rect 143540 649730 143630 649970
rect 143870 649730 143960 649970
rect 144200 649730 144290 649970
rect 144530 649730 144550 649970
rect 133550 649620 144550 649730
rect 133550 649380 133570 649620
rect 133810 649380 133920 649620
rect 134160 649380 134250 649620
rect 134490 649380 134580 649620
rect 134820 649380 134910 649620
rect 135150 649380 135260 649620
rect 135500 649380 135590 649620
rect 135830 649380 135920 649620
rect 136160 649380 136250 649620
rect 136490 649380 136600 649620
rect 136840 649380 136930 649620
rect 137170 649380 137260 649620
rect 137500 649380 137590 649620
rect 137830 649380 137940 649620
rect 138180 649380 138270 649620
rect 138510 649380 138600 649620
rect 138840 649380 138930 649620
rect 139170 649380 139280 649620
rect 139520 649380 139610 649620
rect 139850 649380 139940 649620
rect 140180 649380 140270 649620
rect 140510 649380 140620 649620
rect 140860 649380 140950 649620
rect 141190 649380 141280 649620
rect 141520 649380 141610 649620
rect 141850 649380 141960 649620
rect 142200 649380 142290 649620
rect 142530 649380 142620 649620
rect 142860 649380 142950 649620
rect 143190 649380 143300 649620
rect 143540 649380 143630 649620
rect 143870 649380 143960 649620
rect 144200 649380 144290 649620
rect 144530 649380 144550 649620
rect 133550 649360 144550 649380
rect 144930 660340 155930 660360
rect 144930 660100 144950 660340
rect 145190 660100 145300 660340
rect 145540 660100 145630 660340
rect 145870 660100 145960 660340
rect 146200 660100 146290 660340
rect 146530 660100 146640 660340
rect 146880 660100 146970 660340
rect 147210 660100 147300 660340
rect 147540 660100 147630 660340
rect 147870 660100 147980 660340
rect 148220 660100 148310 660340
rect 148550 660100 148640 660340
rect 148880 660100 148970 660340
rect 149210 660100 149320 660340
rect 149560 660100 149650 660340
rect 149890 660100 149980 660340
rect 150220 660100 150310 660340
rect 150550 660100 150660 660340
rect 150900 660100 150990 660340
rect 151230 660100 151320 660340
rect 151560 660100 151650 660340
rect 151890 660100 152000 660340
rect 152240 660100 152330 660340
rect 152570 660100 152660 660340
rect 152900 660100 152990 660340
rect 153230 660100 153340 660340
rect 153580 660100 153670 660340
rect 153910 660100 154000 660340
rect 154240 660100 154330 660340
rect 154570 660100 154680 660340
rect 154920 660100 155010 660340
rect 155250 660100 155340 660340
rect 155580 660100 155670 660340
rect 155910 660100 155930 660340
rect 144930 660010 155930 660100
rect 144930 659770 144950 660010
rect 145190 659770 145300 660010
rect 145540 659770 145630 660010
rect 145870 659770 145960 660010
rect 146200 659770 146290 660010
rect 146530 659770 146640 660010
rect 146880 659770 146970 660010
rect 147210 659770 147300 660010
rect 147540 659770 147630 660010
rect 147870 659770 147980 660010
rect 148220 659770 148310 660010
rect 148550 659770 148640 660010
rect 148880 659770 148970 660010
rect 149210 659770 149320 660010
rect 149560 659770 149650 660010
rect 149890 659770 149980 660010
rect 150220 659770 150310 660010
rect 150550 659770 150660 660010
rect 150900 659770 150990 660010
rect 151230 659770 151320 660010
rect 151560 659770 151650 660010
rect 151890 659770 152000 660010
rect 152240 659770 152330 660010
rect 152570 659770 152660 660010
rect 152900 659770 152990 660010
rect 153230 659770 153340 660010
rect 153580 659770 153670 660010
rect 153910 659770 154000 660010
rect 154240 659770 154330 660010
rect 154570 659770 154680 660010
rect 154920 659770 155010 660010
rect 155250 659770 155340 660010
rect 155580 659770 155670 660010
rect 155910 659770 155930 660010
rect 144930 659680 155930 659770
rect 144930 659440 144950 659680
rect 145190 659440 145300 659680
rect 145540 659440 145630 659680
rect 145870 659440 145960 659680
rect 146200 659440 146290 659680
rect 146530 659440 146640 659680
rect 146880 659440 146970 659680
rect 147210 659440 147300 659680
rect 147540 659440 147630 659680
rect 147870 659440 147980 659680
rect 148220 659440 148310 659680
rect 148550 659440 148640 659680
rect 148880 659440 148970 659680
rect 149210 659440 149320 659680
rect 149560 659440 149650 659680
rect 149890 659440 149980 659680
rect 150220 659440 150310 659680
rect 150550 659440 150660 659680
rect 150900 659440 150990 659680
rect 151230 659440 151320 659680
rect 151560 659440 151650 659680
rect 151890 659440 152000 659680
rect 152240 659440 152330 659680
rect 152570 659440 152660 659680
rect 152900 659440 152990 659680
rect 153230 659440 153340 659680
rect 153580 659440 153670 659680
rect 153910 659440 154000 659680
rect 154240 659440 154330 659680
rect 154570 659440 154680 659680
rect 154920 659440 155010 659680
rect 155250 659440 155340 659680
rect 155580 659440 155670 659680
rect 155910 659440 155930 659680
rect 144930 659350 155930 659440
rect 144930 659110 144950 659350
rect 145190 659110 145300 659350
rect 145540 659110 145630 659350
rect 145870 659110 145960 659350
rect 146200 659110 146290 659350
rect 146530 659110 146640 659350
rect 146880 659110 146970 659350
rect 147210 659110 147300 659350
rect 147540 659110 147630 659350
rect 147870 659110 147980 659350
rect 148220 659110 148310 659350
rect 148550 659110 148640 659350
rect 148880 659110 148970 659350
rect 149210 659110 149320 659350
rect 149560 659110 149650 659350
rect 149890 659110 149980 659350
rect 150220 659110 150310 659350
rect 150550 659110 150660 659350
rect 150900 659110 150990 659350
rect 151230 659110 151320 659350
rect 151560 659110 151650 659350
rect 151890 659110 152000 659350
rect 152240 659110 152330 659350
rect 152570 659110 152660 659350
rect 152900 659110 152990 659350
rect 153230 659110 153340 659350
rect 153580 659110 153670 659350
rect 153910 659110 154000 659350
rect 154240 659110 154330 659350
rect 154570 659110 154680 659350
rect 154920 659110 155010 659350
rect 155250 659110 155340 659350
rect 155580 659110 155670 659350
rect 155910 659110 155930 659350
rect 144930 659000 155930 659110
rect 144930 658760 144950 659000
rect 145190 658760 145300 659000
rect 145540 658760 145630 659000
rect 145870 658760 145960 659000
rect 146200 658760 146290 659000
rect 146530 658760 146640 659000
rect 146880 658760 146970 659000
rect 147210 658760 147300 659000
rect 147540 658760 147630 659000
rect 147870 658760 147980 659000
rect 148220 658760 148310 659000
rect 148550 658760 148640 659000
rect 148880 658760 148970 659000
rect 149210 658760 149320 659000
rect 149560 658760 149650 659000
rect 149890 658760 149980 659000
rect 150220 658760 150310 659000
rect 150550 658760 150660 659000
rect 150900 658760 150990 659000
rect 151230 658760 151320 659000
rect 151560 658760 151650 659000
rect 151890 658760 152000 659000
rect 152240 658760 152330 659000
rect 152570 658760 152660 659000
rect 152900 658760 152990 659000
rect 153230 658760 153340 659000
rect 153580 658760 153670 659000
rect 153910 658760 154000 659000
rect 154240 658760 154330 659000
rect 154570 658760 154680 659000
rect 154920 658760 155010 659000
rect 155250 658760 155340 659000
rect 155580 658760 155670 659000
rect 155910 658760 155930 659000
rect 144930 658670 155930 658760
rect 144930 658430 144950 658670
rect 145190 658430 145300 658670
rect 145540 658430 145630 658670
rect 145870 658430 145960 658670
rect 146200 658430 146290 658670
rect 146530 658430 146640 658670
rect 146880 658430 146970 658670
rect 147210 658430 147300 658670
rect 147540 658430 147630 658670
rect 147870 658430 147980 658670
rect 148220 658430 148310 658670
rect 148550 658430 148640 658670
rect 148880 658430 148970 658670
rect 149210 658430 149320 658670
rect 149560 658430 149650 658670
rect 149890 658430 149980 658670
rect 150220 658430 150310 658670
rect 150550 658430 150660 658670
rect 150900 658430 150990 658670
rect 151230 658430 151320 658670
rect 151560 658430 151650 658670
rect 151890 658430 152000 658670
rect 152240 658430 152330 658670
rect 152570 658430 152660 658670
rect 152900 658430 152990 658670
rect 153230 658430 153340 658670
rect 153580 658430 153670 658670
rect 153910 658430 154000 658670
rect 154240 658430 154330 658670
rect 154570 658430 154680 658670
rect 154920 658430 155010 658670
rect 155250 658430 155340 658670
rect 155580 658430 155670 658670
rect 155910 658430 155930 658670
rect 144930 658340 155930 658430
rect 144930 658100 144950 658340
rect 145190 658100 145300 658340
rect 145540 658100 145630 658340
rect 145870 658100 145960 658340
rect 146200 658100 146290 658340
rect 146530 658100 146640 658340
rect 146880 658100 146970 658340
rect 147210 658100 147300 658340
rect 147540 658100 147630 658340
rect 147870 658100 147980 658340
rect 148220 658100 148310 658340
rect 148550 658100 148640 658340
rect 148880 658100 148970 658340
rect 149210 658100 149320 658340
rect 149560 658100 149650 658340
rect 149890 658100 149980 658340
rect 150220 658100 150310 658340
rect 150550 658100 150660 658340
rect 150900 658100 150990 658340
rect 151230 658100 151320 658340
rect 151560 658100 151650 658340
rect 151890 658100 152000 658340
rect 152240 658100 152330 658340
rect 152570 658100 152660 658340
rect 152900 658100 152990 658340
rect 153230 658100 153340 658340
rect 153580 658100 153670 658340
rect 153910 658100 154000 658340
rect 154240 658100 154330 658340
rect 154570 658100 154680 658340
rect 154920 658100 155010 658340
rect 155250 658100 155340 658340
rect 155580 658100 155670 658340
rect 155910 658100 155930 658340
rect 144930 658010 155930 658100
rect 144930 657770 144950 658010
rect 145190 657770 145300 658010
rect 145540 657770 145630 658010
rect 145870 657770 145960 658010
rect 146200 657770 146290 658010
rect 146530 657770 146640 658010
rect 146880 657770 146970 658010
rect 147210 657770 147300 658010
rect 147540 657770 147630 658010
rect 147870 657770 147980 658010
rect 148220 657770 148310 658010
rect 148550 657770 148640 658010
rect 148880 657770 148970 658010
rect 149210 657770 149320 658010
rect 149560 657770 149650 658010
rect 149890 657770 149980 658010
rect 150220 657770 150310 658010
rect 150550 657770 150660 658010
rect 150900 657770 150990 658010
rect 151230 657770 151320 658010
rect 151560 657770 151650 658010
rect 151890 657770 152000 658010
rect 152240 657770 152330 658010
rect 152570 657770 152660 658010
rect 152900 657770 152990 658010
rect 153230 657770 153340 658010
rect 153580 657770 153670 658010
rect 153910 657770 154000 658010
rect 154240 657770 154330 658010
rect 154570 657770 154680 658010
rect 154920 657770 155010 658010
rect 155250 657770 155340 658010
rect 155580 657770 155670 658010
rect 155910 657770 155930 658010
rect 144930 657660 155930 657770
rect 144930 657420 144950 657660
rect 145190 657420 145300 657660
rect 145540 657420 145630 657660
rect 145870 657420 145960 657660
rect 146200 657420 146290 657660
rect 146530 657420 146640 657660
rect 146880 657420 146970 657660
rect 147210 657420 147300 657660
rect 147540 657420 147630 657660
rect 147870 657420 147980 657660
rect 148220 657420 148310 657660
rect 148550 657420 148640 657660
rect 148880 657420 148970 657660
rect 149210 657420 149320 657660
rect 149560 657420 149650 657660
rect 149890 657420 149980 657660
rect 150220 657420 150310 657660
rect 150550 657420 150660 657660
rect 150900 657420 150990 657660
rect 151230 657420 151320 657660
rect 151560 657420 151650 657660
rect 151890 657420 152000 657660
rect 152240 657420 152330 657660
rect 152570 657420 152660 657660
rect 152900 657420 152990 657660
rect 153230 657420 153340 657660
rect 153580 657420 153670 657660
rect 153910 657420 154000 657660
rect 154240 657420 154330 657660
rect 154570 657420 154680 657660
rect 154920 657420 155010 657660
rect 155250 657420 155340 657660
rect 155580 657420 155670 657660
rect 155910 657420 155930 657660
rect 144930 657330 155930 657420
rect 144930 657090 144950 657330
rect 145190 657090 145300 657330
rect 145540 657090 145630 657330
rect 145870 657090 145960 657330
rect 146200 657090 146290 657330
rect 146530 657090 146640 657330
rect 146880 657090 146970 657330
rect 147210 657090 147300 657330
rect 147540 657090 147630 657330
rect 147870 657090 147980 657330
rect 148220 657090 148310 657330
rect 148550 657090 148640 657330
rect 148880 657090 148970 657330
rect 149210 657090 149320 657330
rect 149560 657090 149650 657330
rect 149890 657090 149980 657330
rect 150220 657090 150310 657330
rect 150550 657090 150660 657330
rect 150900 657090 150990 657330
rect 151230 657090 151320 657330
rect 151560 657090 151650 657330
rect 151890 657090 152000 657330
rect 152240 657090 152330 657330
rect 152570 657090 152660 657330
rect 152900 657090 152990 657330
rect 153230 657090 153340 657330
rect 153580 657090 153670 657330
rect 153910 657090 154000 657330
rect 154240 657090 154330 657330
rect 154570 657090 154680 657330
rect 154920 657090 155010 657330
rect 155250 657090 155340 657330
rect 155580 657090 155670 657330
rect 155910 657090 155930 657330
rect 144930 657000 155930 657090
rect 144930 656760 144950 657000
rect 145190 656760 145300 657000
rect 145540 656760 145630 657000
rect 145870 656760 145960 657000
rect 146200 656760 146290 657000
rect 146530 656760 146640 657000
rect 146880 656760 146970 657000
rect 147210 656760 147300 657000
rect 147540 656760 147630 657000
rect 147870 656760 147980 657000
rect 148220 656760 148310 657000
rect 148550 656760 148640 657000
rect 148880 656760 148970 657000
rect 149210 656760 149320 657000
rect 149560 656760 149650 657000
rect 149890 656760 149980 657000
rect 150220 656760 150310 657000
rect 150550 656760 150660 657000
rect 150900 656760 150990 657000
rect 151230 656760 151320 657000
rect 151560 656760 151650 657000
rect 151890 656760 152000 657000
rect 152240 656760 152330 657000
rect 152570 656760 152660 657000
rect 152900 656760 152990 657000
rect 153230 656760 153340 657000
rect 153580 656760 153670 657000
rect 153910 656760 154000 657000
rect 154240 656760 154330 657000
rect 154570 656760 154680 657000
rect 154920 656760 155010 657000
rect 155250 656760 155340 657000
rect 155580 656760 155670 657000
rect 155910 656760 155930 657000
rect 144930 656670 155930 656760
rect 144930 656430 144950 656670
rect 145190 656430 145300 656670
rect 145540 656430 145630 656670
rect 145870 656430 145960 656670
rect 146200 656430 146290 656670
rect 146530 656430 146640 656670
rect 146880 656430 146970 656670
rect 147210 656430 147300 656670
rect 147540 656430 147630 656670
rect 147870 656430 147980 656670
rect 148220 656430 148310 656670
rect 148550 656430 148640 656670
rect 148880 656430 148970 656670
rect 149210 656430 149320 656670
rect 149560 656430 149650 656670
rect 149890 656430 149980 656670
rect 150220 656430 150310 656670
rect 150550 656430 150660 656670
rect 150900 656430 150990 656670
rect 151230 656430 151320 656670
rect 151560 656430 151650 656670
rect 151890 656430 152000 656670
rect 152240 656430 152330 656670
rect 152570 656430 152660 656670
rect 152900 656430 152990 656670
rect 153230 656430 153340 656670
rect 153580 656430 153670 656670
rect 153910 656430 154000 656670
rect 154240 656430 154330 656670
rect 154570 656430 154680 656670
rect 154920 656430 155010 656670
rect 155250 656430 155340 656670
rect 155580 656430 155670 656670
rect 155910 656430 155930 656670
rect 144930 656320 155930 656430
rect 144930 656080 144950 656320
rect 145190 656080 145300 656320
rect 145540 656080 145630 656320
rect 145870 656080 145960 656320
rect 146200 656080 146290 656320
rect 146530 656080 146640 656320
rect 146880 656080 146970 656320
rect 147210 656080 147300 656320
rect 147540 656080 147630 656320
rect 147870 656080 147980 656320
rect 148220 656080 148310 656320
rect 148550 656080 148640 656320
rect 148880 656080 148970 656320
rect 149210 656080 149320 656320
rect 149560 656080 149650 656320
rect 149890 656080 149980 656320
rect 150220 656080 150310 656320
rect 150550 656080 150660 656320
rect 150900 656080 150990 656320
rect 151230 656080 151320 656320
rect 151560 656080 151650 656320
rect 151890 656080 152000 656320
rect 152240 656080 152330 656320
rect 152570 656080 152660 656320
rect 152900 656080 152990 656320
rect 153230 656080 153340 656320
rect 153580 656080 153670 656320
rect 153910 656080 154000 656320
rect 154240 656080 154330 656320
rect 154570 656080 154680 656320
rect 154920 656080 155010 656320
rect 155250 656080 155340 656320
rect 155580 656080 155670 656320
rect 155910 656080 155930 656320
rect 144930 655990 155930 656080
rect 144930 655750 144950 655990
rect 145190 655750 145300 655990
rect 145540 655750 145630 655990
rect 145870 655750 145960 655990
rect 146200 655750 146290 655990
rect 146530 655750 146640 655990
rect 146880 655750 146970 655990
rect 147210 655750 147300 655990
rect 147540 655750 147630 655990
rect 147870 655750 147980 655990
rect 148220 655750 148310 655990
rect 148550 655750 148640 655990
rect 148880 655750 148970 655990
rect 149210 655750 149320 655990
rect 149560 655750 149650 655990
rect 149890 655750 149980 655990
rect 150220 655750 150310 655990
rect 150550 655750 150660 655990
rect 150900 655750 150990 655990
rect 151230 655750 151320 655990
rect 151560 655750 151650 655990
rect 151890 655750 152000 655990
rect 152240 655750 152330 655990
rect 152570 655750 152660 655990
rect 152900 655750 152990 655990
rect 153230 655750 153340 655990
rect 153580 655750 153670 655990
rect 153910 655750 154000 655990
rect 154240 655750 154330 655990
rect 154570 655750 154680 655990
rect 154920 655750 155010 655990
rect 155250 655750 155340 655990
rect 155580 655750 155670 655990
rect 155910 655750 155930 655990
rect 144930 655660 155930 655750
rect 144930 655420 144950 655660
rect 145190 655420 145300 655660
rect 145540 655420 145630 655660
rect 145870 655420 145960 655660
rect 146200 655420 146290 655660
rect 146530 655420 146640 655660
rect 146880 655420 146970 655660
rect 147210 655420 147300 655660
rect 147540 655420 147630 655660
rect 147870 655420 147980 655660
rect 148220 655420 148310 655660
rect 148550 655420 148640 655660
rect 148880 655420 148970 655660
rect 149210 655420 149320 655660
rect 149560 655420 149650 655660
rect 149890 655420 149980 655660
rect 150220 655420 150310 655660
rect 150550 655420 150660 655660
rect 150900 655420 150990 655660
rect 151230 655420 151320 655660
rect 151560 655420 151650 655660
rect 151890 655420 152000 655660
rect 152240 655420 152330 655660
rect 152570 655420 152660 655660
rect 152900 655420 152990 655660
rect 153230 655420 153340 655660
rect 153580 655420 153670 655660
rect 153910 655420 154000 655660
rect 154240 655420 154330 655660
rect 154570 655420 154680 655660
rect 154920 655420 155010 655660
rect 155250 655420 155340 655660
rect 155580 655420 155670 655660
rect 155910 655420 155930 655660
rect 144930 655330 155930 655420
rect 144930 655090 144950 655330
rect 145190 655090 145300 655330
rect 145540 655090 145630 655330
rect 145870 655090 145960 655330
rect 146200 655090 146290 655330
rect 146530 655090 146640 655330
rect 146880 655090 146970 655330
rect 147210 655090 147300 655330
rect 147540 655090 147630 655330
rect 147870 655090 147980 655330
rect 148220 655090 148310 655330
rect 148550 655090 148640 655330
rect 148880 655090 148970 655330
rect 149210 655090 149320 655330
rect 149560 655090 149650 655330
rect 149890 655090 149980 655330
rect 150220 655090 150310 655330
rect 150550 655090 150660 655330
rect 150900 655090 150990 655330
rect 151230 655090 151320 655330
rect 151560 655090 151650 655330
rect 151890 655090 152000 655330
rect 152240 655090 152330 655330
rect 152570 655090 152660 655330
rect 152900 655090 152990 655330
rect 153230 655090 153340 655330
rect 153580 655090 153670 655330
rect 153910 655090 154000 655330
rect 154240 655090 154330 655330
rect 154570 655090 154680 655330
rect 154920 655090 155010 655330
rect 155250 655090 155340 655330
rect 155580 655090 155670 655330
rect 155910 655090 155930 655330
rect 144930 654980 155930 655090
rect 144930 654740 144950 654980
rect 145190 654740 145300 654980
rect 145540 654740 145630 654980
rect 145870 654740 145960 654980
rect 146200 654740 146290 654980
rect 146530 654740 146640 654980
rect 146880 654740 146970 654980
rect 147210 654740 147300 654980
rect 147540 654740 147630 654980
rect 147870 654740 147980 654980
rect 148220 654740 148310 654980
rect 148550 654740 148640 654980
rect 148880 654740 148970 654980
rect 149210 654740 149320 654980
rect 149560 654740 149650 654980
rect 149890 654740 149980 654980
rect 150220 654740 150310 654980
rect 150550 654740 150660 654980
rect 150900 654740 150990 654980
rect 151230 654740 151320 654980
rect 151560 654740 151650 654980
rect 151890 654740 152000 654980
rect 152240 654740 152330 654980
rect 152570 654740 152660 654980
rect 152900 654740 152990 654980
rect 153230 654740 153340 654980
rect 153580 654740 153670 654980
rect 153910 654740 154000 654980
rect 154240 654740 154330 654980
rect 154570 654740 154680 654980
rect 154920 654740 155010 654980
rect 155250 654740 155340 654980
rect 155580 654740 155670 654980
rect 155910 654740 155930 654980
rect 144930 654650 155930 654740
rect 144930 654410 144950 654650
rect 145190 654410 145300 654650
rect 145540 654410 145630 654650
rect 145870 654410 145960 654650
rect 146200 654410 146290 654650
rect 146530 654410 146640 654650
rect 146880 654410 146970 654650
rect 147210 654410 147300 654650
rect 147540 654410 147630 654650
rect 147870 654410 147980 654650
rect 148220 654410 148310 654650
rect 148550 654410 148640 654650
rect 148880 654410 148970 654650
rect 149210 654410 149320 654650
rect 149560 654410 149650 654650
rect 149890 654410 149980 654650
rect 150220 654410 150310 654650
rect 150550 654410 150660 654650
rect 150900 654410 150990 654650
rect 151230 654410 151320 654650
rect 151560 654410 151650 654650
rect 151890 654410 152000 654650
rect 152240 654410 152330 654650
rect 152570 654410 152660 654650
rect 152900 654410 152990 654650
rect 153230 654410 153340 654650
rect 153580 654410 153670 654650
rect 153910 654410 154000 654650
rect 154240 654410 154330 654650
rect 154570 654410 154680 654650
rect 154920 654410 155010 654650
rect 155250 654410 155340 654650
rect 155580 654410 155670 654650
rect 155910 654410 155930 654650
rect 144930 654320 155930 654410
rect 144930 654080 144950 654320
rect 145190 654080 145300 654320
rect 145540 654080 145630 654320
rect 145870 654080 145960 654320
rect 146200 654080 146290 654320
rect 146530 654080 146640 654320
rect 146880 654080 146970 654320
rect 147210 654080 147300 654320
rect 147540 654080 147630 654320
rect 147870 654080 147980 654320
rect 148220 654080 148310 654320
rect 148550 654080 148640 654320
rect 148880 654080 148970 654320
rect 149210 654080 149320 654320
rect 149560 654080 149650 654320
rect 149890 654080 149980 654320
rect 150220 654080 150310 654320
rect 150550 654080 150660 654320
rect 150900 654080 150990 654320
rect 151230 654080 151320 654320
rect 151560 654080 151650 654320
rect 151890 654080 152000 654320
rect 152240 654080 152330 654320
rect 152570 654080 152660 654320
rect 152900 654080 152990 654320
rect 153230 654080 153340 654320
rect 153580 654080 153670 654320
rect 153910 654080 154000 654320
rect 154240 654080 154330 654320
rect 154570 654080 154680 654320
rect 154920 654080 155010 654320
rect 155250 654080 155340 654320
rect 155580 654080 155670 654320
rect 155910 654080 155930 654320
rect 144930 653990 155930 654080
rect 144930 653750 144950 653990
rect 145190 653750 145300 653990
rect 145540 653750 145630 653990
rect 145870 653750 145960 653990
rect 146200 653750 146290 653990
rect 146530 653750 146640 653990
rect 146880 653750 146970 653990
rect 147210 653750 147300 653990
rect 147540 653750 147630 653990
rect 147870 653750 147980 653990
rect 148220 653750 148310 653990
rect 148550 653750 148640 653990
rect 148880 653750 148970 653990
rect 149210 653750 149320 653990
rect 149560 653750 149650 653990
rect 149890 653750 149980 653990
rect 150220 653750 150310 653990
rect 150550 653750 150660 653990
rect 150900 653750 150990 653990
rect 151230 653750 151320 653990
rect 151560 653750 151650 653990
rect 151890 653750 152000 653990
rect 152240 653750 152330 653990
rect 152570 653750 152660 653990
rect 152900 653750 152990 653990
rect 153230 653750 153340 653990
rect 153580 653750 153670 653990
rect 153910 653750 154000 653990
rect 154240 653750 154330 653990
rect 154570 653750 154680 653990
rect 154920 653750 155010 653990
rect 155250 653750 155340 653990
rect 155580 653750 155670 653990
rect 155910 653750 155930 653990
rect 144930 653640 155930 653750
rect 144930 653400 144950 653640
rect 145190 653400 145300 653640
rect 145540 653400 145630 653640
rect 145870 653400 145960 653640
rect 146200 653400 146290 653640
rect 146530 653400 146640 653640
rect 146880 653400 146970 653640
rect 147210 653400 147300 653640
rect 147540 653400 147630 653640
rect 147870 653400 147980 653640
rect 148220 653400 148310 653640
rect 148550 653400 148640 653640
rect 148880 653400 148970 653640
rect 149210 653400 149320 653640
rect 149560 653400 149650 653640
rect 149890 653400 149980 653640
rect 150220 653400 150310 653640
rect 150550 653400 150660 653640
rect 150900 653400 150990 653640
rect 151230 653400 151320 653640
rect 151560 653400 151650 653640
rect 151890 653400 152000 653640
rect 152240 653400 152330 653640
rect 152570 653400 152660 653640
rect 152900 653400 152990 653640
rect 153230 653400 153340 653640
rect 153580 653400 153670 653640
rect 153910 653400 154000 653640
rect 154240 653400 154330 653640
rect 154570 653400 154680 653640
rect 154920 653400 155010 653640
rect 155250 653400 155340 653640
rect 155580 653400 155670 653640
rect 155910 653400 155930 653640
rect 144930 653310 155930 653400
rect 144930 653070 144950 653310
rect 145190 653070 145300 653310
rect 145540 653070 145630 653310
rect 145870 653070 145960 653310
rect 146200 653070 146290 653310
rect 146530 653070 146640 653310
rect 146880 653070 146970 653310
rect 147210 653070 147300 653310
rect 147540 653070 147630 653310
rect 147870 653070 147980 653310
rect 148220 653070 148310 653310
rect 148550 653070 148640 653310
rect 148880 653070 148970 653310
rect 149210 653070 149320 653310
rect 149560 653070 149650 653310
rect 149890 653070 149980 653310
rect 150220 653070 150310 653310
rect 150550 653070 150660 653310
rect 150900 653070 150990 653310
rect 151230 653070 151320 653310
rect 151560 653070 151650 653310
rect 151890 653070 152000 653310
rect 152240 653070 152330 653310
rect 152570 653070 152660 653310
rect 152900 653070 152990 653310
rect 153230 653070 153340 653310
rect 153580 653070 153670 653310
rect 153910 653070 154000 653310
rect 154240 653070 154330 653310
rect 154570 653070 154680 653310
rect 154920 653070 155010 653310
rect 155250 653070 155340 653310
rect 155580 653070 155670 653310
rect 155910 653070 155930 653310
rect 144930 652980 155930 653070
rect 144930 652740 144950 652980
rect 145190 652740 145300 652980
rect 145540 652740 145630 652980
rect 145870 652740 145960 652980
rect 146200 652740 146290 652980
rect 146530 652740 146640 652980
rect 146880 652740 146970 652980
rect 147210 652740 147300 652980
rect 147540 652740 147630 652980
rect 147870 652740 147980 652980
rect 148220 652740 148310 652980
rect 148550 652740 148640 652980
rect 148880 652740 148970 652980
rect 149210 652740 149320 652980
rect 149560 652740 149650 652980
rect 149890 652740 149980 652980
rect 150220 652740 150310 652980
rect 150550 652740 150660 652980
rect 150900 652740 150990 652980
rect 151230 652740 151320 652980
rect 151560 652740 151650 652980
rect 151890 652740 152000 652980
rect 152240 652740 152330 652980
rect 152570 652740 152660 652980
rect 152900 652740 152990 652980
rect 153230 652740 153340 652980
rect 153580 652740 153670 652980
rect 153910 652740 154000 652980
rect 154240 652740 154330 652980
rect 154570 652740 154680 652980
rect 154920 652740 155010 652980
rect 155250 652740 155340 652980
rect 155580 652740 155670 652980
rect 155910 652740 155930 652980
rect 144930 652650 155930 652740
rect 144930 652410 144950 652650
rect 145190 652410 145300 652650
rect 145540 652410 145630 652650
rect 145870 652410 145960 652650
rect 146200 652410 146290 652650
rect 146530 652410 146640 652650
rect 146880 652410 146970 652650
rect 147210 652410 147300 652650
rect 147540 652410 147630 652650
rect 147870 652410 147980 652650
rect 148220 652410 148310 652650
rect 148550 652410 148640 652650
rect 148880 652410 148970 652650
rect 149210 652410 149320 652650
rect 149560 652410 149650 652650
rect 149890 652410 149980 652650
rect 150220 652410 150310 652650
rect 150550 652410 150660 652650
rect 150900 652410 150990 652650
rect 151230 652410 151320 652650
rect 151560 652410 151650 652650
rect 151890 652410 152000 652650
rect 152240 652410 152330 652650
rect 152570 652410 152660 652650
rect 152900 652410 152990 652650
rect 153230 652410 153340 652650
rect 153580 652410 153670 652650
rect 153910 652410 154000 652650
rect 154240 652410 154330 652650
rect 154570 652410 154680 652650
rect 154920 652410 155010 652650
rect 155250 652410 155340 652650
rect 155580 652410 155670 652650
rect 155910 652410 155930 652650
rect 144930 652300 155930 652410
rect 144930 652060 144950 652300
rect 145190 652060 145300 652300
rect 145540 652060 145630 652300
rect 145870 652060 145960 652300
rect 146200 652060 146290 652300
rect 146530 652060 146640 652300
rect 146880 652060 146970 652300
rect 147210 652060 147300 652300
rect 147540 652060 147630 652300
rect 147870 652060 147980 652300
rect 148220 652060 148310 652300
rect 148550 652060 148640 652300
rect 148880 652060 148970 652300
rect 149210 652060 149320 652300
rect 149560 652060 149650 652300
rect 149890 652060 149980 652300
rect 150220 652060 150310 652300
rect 150550 652060 150660 652300
rect 150900 652060 150990 652300
rect 151230 652060 151320 652300
rect 151560 652060 151650 652300
rect 151890 652060 152000 652300
rect 152240 652060 152330 652300
rect 152570 652060 152660 652300
rect 152900 652060 152990 652300
rect 153230 652060 153340 652300
rect 153580 652060 153670 652300
rect 153910 652060 154000 652300
rect 154240 652060 154330 652300
rect 154570 652060 154680 652300
rect 154920 652060 155010 652300
rect 155250 652060 155340 652300
rect 155580 652060 155670 652300
rect 155910 652060 155930 652300
rect 144930 651970 155930 652060
rect 144930 651730 144950 651970
rect 145190 651730 145300 651970
rect 145540 651730 145630 651970
rect 145870 651730 145960 651970
rect 146200 651730 146290 651970
rect 146530 651730 146640 651970
rect 146880 651730 146970 651970
rect 147210 651730 147300 651970
rect 147540 651730 147630 651970
rect 147870 651730 147980 651970
rect 148220 651730 148310 651970
rect 148550 651730 148640 651970
rect 148880 651730 148970 651970
rect 149210 651730 149320 651970
rect 149560 651730 149650 651970
rect 149890 651730 149980 651970
rect 150220 651730 150310 651970
rect 150550 651730 150660 651970
rect 150900 651730 150990 651970
rect 151230 651730 151320 651970
rect 151560 651730 151650 651970
rect 151890 651730 152000 651970
rect 152240 651730 152330 651970
rect 152570 651730 152660 651970
rect 152900 651730 152990 651970
rect 153230 651730 153340 651970
rect 153580 651730 153670 651970
rect 153910 651730 154000 651970
rect 154240 651730 154330 651970
rect 154570 651730 154680 651970
rect 154920 651730 155010 651970
rect 155250 651730 155340 651970
rect 155580 651730 155670 651970
rect 155910 651730 155930 651970
rect 144930 651640 155930 651730
rect 144930 651400 144950 651640
rect 145190 651400 145300 651640
rect 145540 651400 145630 651640
rect 145870 651400 145960 651640
rect 146200 651400 146290 651640
rect 146530 651400 146640 651640
rect 146880 651400 146970 651640
rect 147210 651400 147300 651640
rect 147540 651400 147630 651640
rect 147870 651400 147980 651640
rect 148220 651400 148310 651640
rect 148550 651400 148640 651640
rect 148880 651400 148970 651640
rect 149210 651400 149320 651640
rect 149560 651400 149650 651640
rect 149890 651400 149980 651640
rect 150220 651400 150310 651640
rect 150550 651400 150660 651640
rect 150900 651400 150990 651640
rect 151230 651400 151320 651640
rect 151560 651400 151650 651640
rect 151890 651400 152000 651640
rect 152240 651400 152330 651640
rect 152570 651400 152660 651640
rect 152900 651400 152990 651640
rect 153230 651400 153340 651640
rect 153580 651400 153670 651640
rect 153910 651400 154000 651640
rect 154240 651400 154330 651640
rect 154570 651400 154680 651640
rect 154920 651400 155010 651640
rect 155250 651400 155340 651640
rect 155580 651400 155670 651640
rect 155910 651400 155930 651640
rect 144930 651310 155930 651400
rect 144930 651070 144950 651310
rect 145190 651070 145300 651310
rect 145540 651070 145630 651310
rect 145870 651070 145960 651310
rect 146200 651070 146290 651310
rect 146530 651070 146640 651310
rect 146880 651070 146970 651310
rect 147210 651070 147300 651310
rect 147540 651070 147630 651310
rect 147870 651070 147980 651310
rect 148220 651070 148310 651310
rect 148550 651070 148640 651310
rect 148880 651070 148970 651310
rect 149210 651070 149320 651310
rect 149560 651070 149650 651310
rect 149890 651070 149980 651310
rect 150220 651070 150310 651310
rect 150550 651070 150660 651310
rect 150900 651070 150990 651310
rect 151230 651070 151320 651310
rect 151560 651070 151650 651310
rect 151890 651070 152000 651310
rect 152240 651070 152330 651310
rect 152570 651070 152660 651310
rect 152900 651070 152990 651310
rect 153230 651070 153340 651310
rect 153580 651070 153670 651310
rect 153910 651070 154000 651310
rect 154240 651070 154330 651310
rect 154570 651070 154680 651310
rect 154920 651070 155010 651310
rect 155250 651070 155340 651310
rect 155580 651070 155670 651310
rect 155910 651070 155930 651310
rect 144930 650960 155930 651070
rect 144930 650720 144950 650960
rect 145190 650720 145300 650960
rect 145540 650720 145630 650960
rect 145870 650720 145960 650960
rect 146200 650720 146290 650960
rect 146530 650720 146640 650960
rect 146880 650720 146970 650960
rect 147210 650720 147300 650960
rect 147540 650720 147630 650960
rect 147870 650720 147980 650960
rect 148220 650720 148310 650960
rect 148550 650720 148640 650960
rect 148880 650720 148970 650960
rect 149210 650720 149320 650960
rect 149560 650720 149650 650960
rect 149890 650720 149980 650960
rect 150220 650720 150310 650960
rect 150550 650720 150660 650960
rect 150900 650720 150990 650960
rect 151230 650720 151320 650960
rect 151560 650720 151650 650960
rect 151890 650720 152000 650960
rect 152240 650720 152330 650960
rect 152570 650720 152660 650960
rect 152900 650720 152990 650960
rect 153230 650720 153340 650960
rect 153580 650720 153670 650960
rect 153910 650720 154000 650960
rect 154240 650720 154330 650960
rect 154570 650720 154680 650960
rect 154920 650720 155010 650960
rect 155250 650720 155340 650960
rect 155580 650720 155670 650960
rect 155910 650720 155930 650960
rect 144930 650630 155930 650720
rect 144930 650390 144950 650630
rect 145190 650390 145300 650630
rect 145540 650390 145630 650630
rect 145870 650390 145960 650630
rect 146200 650390 146290 650630
rect 146530 650390 146640 650630
rect 146880 650390 146970 650630
rect 147210 650390 147300 650630
rect 147540 650390 147630 650630
rect 147870 650390 147980 650630
rect 148220 650390 148310 650630
rect 148550 650390 148640 650630
rect 148880 650390 148970 650630
rect 149210 650390 149320 650630
rect 149560 650390 149650 650630
rect 149890 650390 149980 650630
rect 150220 650390 150310 650630
rect 150550 650390 150660 650630
rect 150900 650390 150990 650630
rect 151230 650390 151320 650630
rect 151560 650390 151650 650630
rect 151890 650390 152000 650630
rect 152240 650390 152330 650630
rect 152570 650390 152660 650630
rect 152900 650390 152990 650630
rect 153230 650390 153340 650630
rect 153580 650390 153670 650630
rect 153910 650390 154000 650630
rect 154240 650390 154330 650630
rect 154570 650390 154680 650630
rect 154920 650390 155010 650630
rect 155250 650390 155340 650630
rect 155580 650390 155670 650630
rect 155910 650390 155930 650630
rect 144930 650300 155930 650390
rect 144930 650060 144950 650300
rect 145190 650060 145300 650300
rect 145540 650060 145630 650300
rect 145870 650060 145960 650300
rect 146200 650060 146290 650300
rect 146530 650060 146640 650300
rect 146880 650060 146970 650300
rect 147210 650060 147300 650300
rect 147540 650060 147630 650300
rect 147870 650060 147980 650300
rect 148220 650060 148310 650300
rect 148550 650060 148640 650300
rect 148880 650060 148970 650300
rect 149210 650060 149320 650300
rect 149560 650060 149650 650300
rect 149890 650060 149980 650300
rect 150220 650060 150310 650300
rect 150550 650060 150660 650300
rect 150900 650060 150990 650300
rect 151230 650060 151320 650300
rect 151560 650060 151650 650300
rect 151890 650060 152000 650300
rect 152240 650060 152330 650300
rect 152570 650060 152660 650300
rect 152900 650060 152990 650300
rect 153230 650060 153340 650300
rect 153580 650060 153670 650300
rect 153910 650060 154000 650300
rect 154240 650060 154330 650300
rect 154570 650060 154680 650300
rect 154920 650060 155010 650300
rect 155250 650060 155340 650300
rect 155580 650060 155670 650300
rect 155910 650060 155930 650300
rect 144930 649970 155930 650060
rect 144930 649730 144950 649970
rect 145190 649730 145300 649970
rect 145540 649730 145630 649970
rect 145870 649730 145960 649970
rect 146200 649730 146290 649970
rect 146530 649730 146640 649970
rect 146880 649730 146970 649970
rect 147210 649730 147300 649970
rect 147540 649730 147630 649970
rect 147870 649730 147980 649970
rect 148220 649730 148310 649970
rect 148550 649730 148640 649970
rect 148880 649730 148970 649970
rect 149210 649730 149320 649970
rect 149560 649730 149650 649970
rect 149890 649730 149980 649970
rect 150220 649730 150310 649970
rect 150550 649730 150660 649970
rect 150900 649730 150990 649970
rect 151230 649730 151320 649970
rect 151560 649730 151650 649970
rect 151890 649730 152000 649970
rect 152240 649730 152330 649970
rect 152570 649730 152660 649970
rect 152900 649730 152990 649970
rect 153230 649730 153340 649970
rect 153580 649730 153670 649970
rect 153910 649730 154000 649970
rect 154240 649730 154330 649970
rect 154570 649730 154680 649970
rect 154920 649730 155010 649970
rect 155250 649730 155340 649970
rect 155580 649730 155670 649970
rect 155910 649730 155930 649970
rect 144930 649620 155930 649730
rect 144930 649380 144950 649620
rect 145190 649380 145300 649620
rect 145540 649380 145630 649620
rect 145870 649380 145960 649620
rect 146200 649380 146290 649620
rect 146530 649380 146640 649620
rect 146880 649380 146970 649620
rect 147210 649380 147300 649620
rect 147540 649380 147630 649620
rect 147870 649380 147980 649620
rect 148220 649380 148310 649620
rect 148550 649380 148640 649620
rect 148880 649380 148970 649620
rect 149210 649380 149320 649620
rect 149560 649380 149650 649620
rect 149890 649380 149980 649620
rect 150220 649380 150310 649620
rect 150550 649380 150660 649620
rect 150900 649380 150990 649620
rect 151230 649380 151320 649620
rect 151560 649380 151650 649620
rect 151890 649380 152000 649620
rect 152240 649380 152330 649620
rect 152570 649380 152660 649620
rect 152900 649380 152990 649620
rect 153230 649380 153340 649620
rect 153580 649380 153670 649620
rect 153910 649380 154000 649620
rect 154240 649380 154330 649620
rect 154570 649380 154680 649620
rect 154920 649380 155010 649620
rect 155250 649380 155340 649620
rect 155580 649380 155670 649620
rect 155910 649380 155930 649620
rect 144930 649360 155930 649380
<< mimcapcontact >>
rect 110810 694600 111050 694840
rect 111140 694600 111380 694840
rect 111470 694600 111710 694840
rect 111800 694600 112040 694840
rect 112150 694600 112390 694840
rect 112480 694600 112720 694840
rect 112810 694600 113050 694840
rect 113140 694600 113380 694840
rect 113490 694600 113730 694840
rect 113820 694600 114060 694840
rect 114150 694600 114390 694840
rect 114480 694600 114720 694840
rect 114830 694600 115070 694840
rect 115160 694600 115400 694840
rect 115490 694600 115730 694840
rect 115820 694600 116060 694840
rect 116170 694600 116410 694840
rect 116500 694600 116740 694840
rect 116830 694600 117070 694840
rect 117160 694600 117400 694840
rect 117510 694600 117750 694840
rect 117840 694600 118080 694840
rect 118170 694600 118410 694840
rect 118500 694600 118740 694840
rect 118850 694600 119090 694840
rect 119180 694600 119420 694840
rect 119510 694600 119750 694840
rect 119840 694600 120080 694840
rect 120190 694600 120430 694840
rect 120520 694600 120760 694840
rect 120850 694600 121090 694840
rect 121180 694600 121420 694840
rect 121530 694600 121770 694840
rect 110810 694250 111050 694490
rect 111140 694250 111380 694490
rect 111470 694250 111710 694490
rect 111800 694250 112040 694490
rect 112150 694250 112390 694490
rect 112480 694250 112720 694490
rect 112810 694250 113050 694490
rect 113140 694250 113380 694490
rect 113490 694250 113730 694490
rect 113820 694250 114060 694490
rect 114150 694250 114390 694490
rect 114480 694250 114720 694490
rect 114830 694250 115070 694490
rect 115160 694250 115400 694490
rect 115490 694250 115730 694490
rect 115820 694250 116060 694490
rect 116170 694250 116410 694490
rect 116500 694250 116740 694490
rect 116830 694250 117070 694490
rect 117160 694250 117400 694490
rect 117510 694250 117750 694490
rect 117840 694250 118080 694490
rect 118170 694250 118410 694490
rect 118500 694250 118740 694490
rect 118850 694250 119090 694490
rect 119180 694250 119420 694490
rect 119510 694250 119750 694490
rect 119840 694250 120080 694490
rect 120190 694250 120430 694490
rect 120520 694250 120760 694490
rect 120850 694250 121090 694490
rect 121180 694250 121420 694490
rect 121530 694250 121770 694490
rect 110810 693920 111050 694160
rect 111140 693920 111380 694160
rect 111470 693920 111710 694160
rect 111800 693920 112040 694160
rect 112150 693920 112390 694160
rect 112480 693920 112720 694160
rect 112810 693920 113050 694160
rect 113140 693920 113380 694160
rect 113490 693920 113730 694160
rect 113820 693920 114060 694160
rect 114150 693920 114390 694160
rect 114480 693920 114720 694160
rect 114830 693920 115070 694160
rect 115160 693920 115400 694160
rect 115490 693920 115730 694160
rect 115820 693920 116060 694160
rect 116170 693920 116410 694160
rect 116500 693920 116740 694160
rect 116830 693920 117070 694160
rect 117160 693920 117400 694160
rect 117510 693920 117750 694160
rect 117840 693920 118080 694160
rect 118170 693920 118410 694160
rect 118500 693920 118740 694160
rect 118850 693920 119090 694160
rect 119180 693920 119420 694160
rect 119510 693920 119750 694160
rect 119840 693920 120080 694160
rect 120190 693920 120430 694160
rect 120520 693920 120760 694160
rect 120850 693920 121090 694160
rect 121180 693920 121420 694160
rect 121530 693920 121770 694160
rect 110810 693590 111050 693830
rect 111140 693590 111380 693830
rect 111470 693590 111710 693830
rect 111800 693590 112040 693830
rect 112150 693590 112390 693830
rect 112480 693590 112720 693830
rect 112810 693590 113050 693830
rect 113140 693590 113380 693830
rect 113490 693590 113730 693830
rect 113820 693590 114060 693830
rect 114150 693590 114390 693830
rect 114480 693590 114720 693830
rect 114830 693590 115070 693830
rect 115160 693590 115400 693830
rect 115490 693590 115730 693830
rect 115820 693590 116060 693830
rect 116170 693590 116410 693830
rect 116500 693590 116740 693830
rect 116830 693590 117070 693830
rect 117160 693590 117400 693830
rect 117510 693590 117750 693830
rect 117840 693590 118080 693830
rect 118170 693590 118410 693830
rect 118500 693590 118740 693830
rect 118850 693590 119090 693830
rect 119180 693590 119420 693830
rect 119510 693590 119750 693830
rect 119840 693590 120080 693830
rect 120190 693590 120430 693830
rect 120520 693590 120760 693830
rect 120850 693590 121090 693830
rect 121180 693590 121420 693830
rect 121530 693590 121770 693830
rect 110810 693260 111050 693500
rect 111140 693260 111380 693500
rect 111470 693260 111710 693500
rect 111800 693260 112040 693500
rect 112150 693260 112390 693500
rect 112480 693260 112720 693500
rect 112810 693260 113050 693500
rect 113140 693260 113380 693500
rect 113490 693260 113730 693500
rect 113820 693260 114060 693500
rect 114150 693260 114390 693500
rect 114480 693260 114720 693500
rect 114830 693260 115070 693500
rect 115160 693260 115400 693500
rect 115490 693260 115730 693500
rect 115820 693260 116060 693500
rect 116170 693260 116410 693500
rect 116500 693260 116740 693500
rect 116830 693260 117070 693500
rect 117160 693260 117400 693500
rect 117510 693260 117750 693500
rect 117840 693260 118080 693500
rect 118170 693260 118410 693500
rect 118500 693260 118740 693500
rect 118850 693260 119090 693500
rect 119180 693260 119420 693500
rect 119510 693260 119750 693500
rect 119840 693260 120080 693500
rect 120190 693260 120430 693500
rect 120520 693260 120760 693500
rect 120850 693260 121090 693500
rect 121180 693260 121420 693500
rect 121530 693260 121770 693500
rect 110810 692910 111050 693150
rect 111140 692910 111380 693150
rect 111470 692910 111710 693150
rect 111800 692910 112040 693150
rect 112150 692910 112390 693150
rect 112480 692910 112720 693150
rect 112810 692910 113050 693150
rect 113140 692910 113380 693150
rect 113490 692910 113730 693150
rect 113820 692910 114060 693150
rect 114150 692910 114390 693150
rect 114480 692910 114720 693150
rect 114830 692910 115070 693150
rect 115160 692910 115400 693150
rect 115490 692910 115730 693150
rect 115820 692910 116060 693150
rect 116170 692910 116410 693150
rect 116500 692910 116740 693150
rect 116830 692910 117070 693150
rect 117160 692910 117400 693150
rect 117510 692910 117750 693150
rect 117840 692910 118080 693150
rect 118170 692910 118410 693150
rect 118500 692910 118740 693150
rect 118850 692910 119090 693150
rect 119180 692910 119420 693150
rect 119510 692910 119750 693150
rect 119840 692910 120080 693150
rect 120190 692910 120430 693150
rect 120520 692910 120760 693150
rect 120850 692910 121090 693150
rect 121180 692910 121420 693150
rect 121530 692910 121770 693150
rect 110810 692580 111050 692820
rect 111140 692580 111380 692820
rect 111470 692580 111710 692820
rect 111800 692580 112040 692820
rect 112150 692580 112390 692820
rect 112480 692580 112720 692820
rect 112810 692580 113050 692820
rect 113140 692580 113380 692820
rect 113490 692580 113730 692820
rect 113820 692580 114060 692820
rect 114150 692580 114390 692820
rect 114480 692580 114720 692820
rect 114830 692580 115070 692820
rect 115160 692580 115400 692820
rect 115490 692580 115730 692820
rect 115820 692580 116060 692820
rect 116170 692580 116410 692820
rect 116500 692580 116740 692820
rect 116830 692580 117070 692820
rect 117160 692580 117400 692820
rect 117510 692580 117750 692820
rect 117840 692580 118080 692820
rect 118170 692580 118410 692820
rect 118500 692580 118740 692820
rect 118850 692580 119090 692820
rect 119180 692580 119420 692820
rect 119510 692580 119750 692820
rect 119840 692580 120080 692820
rect 120190 692580 120430 692820
rect 120520 692580 120760 692820
rect 120850 692580 121090 692820
rect 121180 692580 121420 692820
rect 121530 692580 121770 692820
rect 110810 692250 111050 692490
rect 111140 692250 111380 692490
rect 111470 692250 111710 692490
rect 111800 692250 112040 692490
rect 112150 692250 112390 692490
rect 112480 692250 112720 692490
rect 112810 692250 113050 692490
rect 113140 692250 113380 692490
rect 113490 692250 113730 692490
rect 113820 692250 114060 692490
rect 114150 692250 114390 692490
rect 114480 692250 114720 692490
rect 114830 692250 115070 692490
rect 115160 692250 115400 692490
rect 115490 692250 115730 692490
rect 115820 692250 116060 692490
rect 116170 692250 116410 692490
rect 116500 692250 116740 692490
rect 116830 692250 117070 692490
rect 117160 692250 117400 692490
rect 117510 692250 117750 692490
rect 117840 692250 118080 692490
rect 118170 692250 118410 692490
rect 118500 692250 118740 692490
rect 118850 692250 119090 692490
rect 119180 692250 119420 692490
rect 119510 692250 119750 692490
rect 119840 692250 120080 692490
rect 120190 692250 120430 692490
rect 120520 692250 120760 692490
rect 120850 692250 121090 692490
rect 121180 692250 121420 692490
rect 121530 692250 121770 692490
rect 110810 691920 111050 692160
rect 111140 691920 111380 692160
rect 111470 691920 111710 692160
rect 111800 691920 112040 692160
rect 112150 691920 112390 692160
rect 112480 691920 112720 692160
rect 112810 691920 113050 692160
rect 113140 691920 113380 692160
rect 113490 691920 113730 692160
rect 113820 691920 114060 692160
rect 114150 691920 114390 692160
rect 114480 691920 114720 692160
rect 114830 691920 115070 692160
rect 115160 691920 115400 692160
rect 115490 691920 115730 692160
rect 115820 691920 116060 692160
rect 116170 691920 116410 692160
rect 116500 691920 116740 692160
rect 116830 691920 117070 692160
rect 117160 691920 117400 692160
rect 117510 691920 117750 692160
rect 117840 691920 118080 692160
rect 118170 691920 118410 692160
rect 118500 691920 118740 692160
rect 118850 691920 119090 692160
rect 119180 691920 119420 692160
rect 119510 691920 119750 692160
rect 119840 691920 120080 692160
rect 120190 691920 120430 692160
rect 120520 691920 120760 692160
rect 120850 691920 121090 692160
rect 121180 691920 121420 692160
rect 121530 691920 121770 692160
rect 110810 691570 111050 691810
rect 111140 691570 111380 691810
rect 111470 691570 111710 691810
rect 111800 691570 112040 691810
rect 112150 691570 112390 691810
rect 112480 691570 112720 691810
rect 112810 691570 113050 691810
rect 113140 691570 113380 691810
rect 113490 691570 113730 691810
rect 113820 691570 114060 691810
rect 114150 691570 114390 691810
rect 114480 691570 114720 691810
rect 114830 691570 115070 691810
rect 115160 691570 115400 691810
rect 115490 691570 115730 691810
rect 115820 691570 116060 691810
rect 116170 691570 116410 691810
rect 116500 691570 116740 691810
rect 116830 691570 117070 691810
rect 117160 691570 117400 691810
rect 117510 691570 117750 691810
rect 117840 691570 118080 691810
rect 118170 691570 118410 691810
rect 118500 691570 118740 691810
rect 118850 691570 119090 691810
rect 119180 691570 119420 691810
rect 119510 691570 119750 691810
rect 119840 691570 120080 691810
rect 120190 691570 120430 691810
rect 120520 691570 120760 691810
rect 120850 691570 121090 691810
rect 121180 691570 121420 691810
rect 121530 691570 121770 691810
rect 110810 691240 111050 691480
rect 111140 691240 111380 691480
rect 111470 691240 111710 691480
rect 111800 691240 112040 691480
rect 112150 691240 112390 691480
rect 112480 691240 112720 691480
rect 112810 691240 113050 691480
rect 113140 691240 113380 691480
rect 113490 691240 113730 691480
rect 113820 691240 114060 691480
rect 114150 691240 114390 691480
rect 114480 691240 114720 691480
rect 114830 691240 115070 691480
rect 115160 691240 115400 691480
rect 115490 691240 115730 691480
rect 115820 691240 116060 691480
rect 116170 691240 116410 691480
rect 116500 691240 116740 691480
rect 116830 691240 117070 691480
rect 117160 691240 117400 691480
rect 117510 691240 117750 691480
rect 117840 691240 118080 691480
rect 118170 691240 118410 691480
rect 118500 691240 118740 691480
rect 118850 691240 119090 691480
rect 119180 691240 119420 691480
rect 119510 691240 119750 691480
rect 119840 691240 120080 691480
rect 120190 691240 120430 691480
rect 120520 691240 120760 691480
rect 120850 691240 121090 691480
rect 121180 691240 121420 691480
rect 121530 691240 121770 691480
rect 110810 690910 111050 691150
rect 111140 690910 111380 691150
rect 111470 690910 111710 691150
rect 111800 690910 112040 691150
rect 112150 690910 112390 691150
rect 112480 690910 112720 691150
rect 112810 690910 113050 691150
rect 113140 690910 113380 691150
rect 113490 690910 113730 691150
rect 113820 690910 114060 691150
rect 114150 690910 114390 691150
rect 114480 690910 114720 691150
rect 114830 690910 115070 691150
rect 115160 690910 115400 691150
rect 115490 690910 115730 691150
rect 115820 690910 116060 691150
rect 116170 690910 116410 691150
rect 116500 690910 116740 691150
rect 116830 690910 117070 691150
rect 117160 690910 117400 691150
rect 117510 690910 117750 691150
rect 117840 690910 118080 691150
rect 118170 690910 118410 691150
rect 118500 690910 118740 691150
rect 118850 690910 119090 691150
rect 119180 690910 119420 691150
rect 119510 690910 119750 691150
rect 119840 690910 120080 691150
rect 120190 690910 120430 691150
rect 120520 690910 120760 691150
rect 120850 690910 121090 691150
rect 121180 690910 121420 691150
rect 121530 690910 121770 691150
rect 110810 690580 111050 690820
rect 111140 690580 111380 690820
rect 111470 690580 111710 690820
rect 111800 690580 112040 690820
rect 112150 690580 112390 690820
rect 112480 690580 112720 690820
rect 112810 690580 113050 690820
rect 113140 690580 113380 690820
rect 113490 690580 113730 690820
rect 113820 690580 114060 690820
rect 114150 690580 114390 690820
rect 114480 690580 114720 690820
rect 114830 690580 115070 690820
rect 115160 690580 115400 690820
rect 115490 690580 115730 690820
rect 115820 690580 116060 690820
rect 116170 690580 116410 690820
rect 116500 690580 116740 690820
rect 116830 690580 117070 690820
rect 117160 690580 117400 690820
rect 117510 690580 117750 690820
rect 117840 690580 118080 690820
rect 118170 690580 118410 690820
rect 118500 690580 118740 690820
rect 118850 690580 119090 690820
rect 119180 690580 119420 690820
rect 119510 690580 119750 690820
rect 119840 690580 120080 690820
rect 120190 690580 120430 690820
rect 120520 690580 120760 690820
rect 120850 690580 121090 690820
rect 121180 690580 121420 690820
rect 121530 690580 121770 690820
rect 110810 690230 111050 690470
rect 111140 690230 111380 690470
rect 111470 690230 111710 690470
rect 111800 690230 112040 690470
rect 112150 690230 112390 690470
rect 112480 690230 112720 690470
rect 112810 690230 113050 690470
rect 113140 690230 113380 690470
rect 113490 690230 113730 690470
rect 113820 690230 114060 690470
rect 114150 690230 114390 690470
rect 114480 690230 114720 690470
rect 114830 690230 115070 690470
rect 115160 690230 115400 690470
rect 115490 690230 115730 690470
rect 115820 690230 116060 690470
rect 116170 690230 116410 690470
rect 116500 690230 116740 690470
rect 116830 690230 117070 690470
rect 117160 690230 117400 690470
rect 117510 690230 117750 690470
rect 117840 690230 118080 690470
rect 118170 690230 118410 690470
rect 118500 690230 118740 690470
rect 118850 690230 119090 690470
rect 119180 690230 119420 690470
rect 119510 690230 119750 690470
rect 119840 690230 120080 690470
rect 120190 690230 120430 690470
rect 120520 690230 120760 690470
rect 120850 690230 121090 690470
rect 121180 690230 121420 690470
rect 121530 690230 121770 690470
rect 110810 689900 111050 690140
rect 111140 689900 111380 690140
rect 111470 689900 111710 690140
rect 111800 689900 112040 690140
rect 112150 689900 112390 690140
rect 112480 689900 112720 690140
rect 112810 689900 113050 690140
rect 113140 689900 113380 690140
rect 113490 689900 113730 690140
rect 113820 689900 114060 690140
rect 114150 689900 114390 690140
rect 114480 689900 114720 690140
rect 114830 689900 115070 690140
rect 115160 689900 115400 690140
rect 115490 689900 115730 690140
rect 115820 689900 116060 690140
rect 116170 689900 116410 690140
rect 116500 689900 116740 690140
rect 116830 689900 117070 690140
rect 117160 689900 117400 690140
rect 117510 689900 117750 690140
rect 117840 689900 118080 690140
rect 118170 689900 118410 690140
rect 118500 689900 118740 690140
rect 118850 689900 119090 690140
rect 119180 689900 119420 690140
rect 119510 689900 119750 690140
rect 119840 689900 120080 690140
rect 120190 689900 120430 690140
rect 120520 689900 120760 690140
rect 120850 689900 121090 690140
rect 121180 689900 121420 690140
rect 121530 689900 121770 690140
rect 110810 689570 111050 689810
rect 111140 689570 111380 689810
rect 111470 689570 111710 689810
rect 111800 689570 112040 689810
rect 112150 689570 112390 689810
rect 112480 689570 112720 689810
rect 112810 689570 113050 689810
rect 113140 689570 113380 689810
rect 113490 689570 113730 689810
rect 113820 689570 114060 689810
rect 114150 689570 114390 689810
rect 114480 689570 114720 689810
rect 114830 689570 115070 689810
rect 115160 689570 115400 689810
rect 115490 689570 115730 689810
rect 115820 689570 116060 689810
rect 116170 689570 116410 689810
rect 116500 689570 116740 689810
rect 116830 689570 117070 689810
rect 117160 689570 117400 689810
rect 117510 689570 117750 689810
rect 117840 689570 118080 689810
rect 118170 689570 118410 689810
rect 118500 689570 118740 689810
rect 118850 689570 119090 689810
rect 119180 689570 119420 689810
rect 119510 689570 119750 689810
rect 119840 689570 120080 689810
rect 120190 689570 120430 689810
rect 120520 689570 120760 689810
rect 120850 689570 121090 689810
rect 121180 689570 121420 689810
rect 121530 689570 121770 689810
rect 110810 689240 111050 689480
rect 111140 689240 111380 689480
rect 111470 689240 111710 689480
rect 111800 689240 112040 689480
rect 112150 689240 112390 689480
rect 112480 689240 112720 689480
rect 112810 689240 113050 689480
rect 113140 689240 113380 689480
rect 113490 689240 113730 689480
rect 113820 689240 114060 689480
rect 114150 689240 114390 689480
rect 114480 689240 114720 689480
rect 114830 689240 115070 689480
rect 115160 689240 115400 689480
rect 115490 689240 115730 689480
rect 115820 689240 116060 689480
rect 116170 689240 116410 689480
rect 116500 689240 116740 689480
rect 116830 689240 117070 689480
rect 117160 689240 117400 689480
rect 117510 689240 117750 689480
rect 117840 689240 118080 689480
rect 118170 689240 118410 689480
rect 118500 689240 118740 689480
rect 118850 689240 119090 689480
rect 119180 689240 119420 689480
rect 119510 689240 119750 689480
rect 119840 689240 120080 689480
rect 120190 689240 120430 689480
rect 120520 689240 120760 689480
rect 120850 689240 121090 689480
rect 121180 689240 121420 689480
rect 121530 689240 121770 689480
rect 110810 688890 111050 689130
rect 111140 688890 111380 689130
rect 111470 688890 111710 689130
rect 111800 688890 112040 689130
rect 112150 688890 112390 689130
rect 112480 688890 112720 689130
rect 112810 688890 113050 689130
rect 113140 688890 113380 689130
rect 113490 688890 113730 689130
rect 113820 688890 114060 689130
rect 114150 688890 114390 689130
rect 114480 688890 114720 689130
rect 114830 688890 115070 689130
rect 115160 688890 115400 689130
rect 115490 688890 115730 689130
rect 115820 688890 116060 689130
rect 116170 688890 116410 689130
rect 116500 688890 116740 689130
rect 116830 688890 117070 689130
rect 117160 688890 117400 689130
rect 117510 688890 117750 689130
rect 117840 688890 118080 689130
rect 118170 688890 118410 689130
rect 118500 688890 118740 689130
rect 118850 688890 119090 689130
rect 119180 688890 119420 689130
rect 119510 688890 119750 689130
rect 119840 688890 120080 689130
rect 120190 688890 120430 689130
rect 120520 688890 120760 689130
rect 120850 688890 121090 689130
rect 121180 688890 121420 689130
rect 121530 688890 121770 689130
rect 110810 688560 111050 688800
rect 111140 688560 111380 688800
rect 111470 688560 111710 688800
rect 111800 688560 112040 688800
rect 112150 688560 112390 688800
rect 112480 688560 112720 688800
rect 112810 688560 113050 688800
rect 113140 688560 113380 688800
rect 113490 688560 113730 688800
rect 113820 688560 114060 688800
rect 114150 688560 114390 688800
rect 114480 688560 114720 688800
rect 114830 688560 115070 688800
rect 115160 688560 115400 688800
rect 115490 688560 115730 688800
rect 115820 688560 116060 688800
rect 116170 688560 116410 688800
rect 116500 688560 116740 688800
rect 116830 688560 117070 688800
rect 117160 688560 117400 688800
rect 117510 688560 117750 688800
rect 117840 688560 118080 688800
rect 118170 688560 118410 688800
rect 118500 688560 118740 688800
rect 118850 688560 119090 688800
rect 119180 688560 119420 688800
rect 119510 688560 119750 688800
rect 119840 688560 120080 688800
rect 120190 688560 120430 688800
rect 120520 688560 120760 688800
rect 120850 688560 121090 688800
rect 121180 688560 121420 688800
rect 121530 688560 121770 688800
rect 110810 688230 111050 688470
rect 111140 688230 111380 688470
rect 111470 688230 111710 688470
rect 111800 688230 112040 688470
rect 112150 688230 112390 688470
rect 112480 688230 112720 688470
rect 112810 688230 113050 688470
rect 113140 688230 113380 688470
rect 113490 688230 113730 688470
rect 113820 688230 114060 688470
rect 114150 688230 114390 688470
rect 114480 688230 114720 688470
rect 114830 688230 115070 688470
rect 115160 688230 115400 688470
rect 115490 688230 115730 688470
rect 115820 688230 116060 688470
rect 116170 688230 116410 688470
rect 116500 688230 116740 688470
rect 116830 688230 117070 688470
rect 117160 688230 117400 688470
rect 117510 688230 117750 688470
rect 117840 688230 118080 688470
rect 118170 688230 118410 688470
rect 118500 688230 118740 688470
rect 118850 688230 119090 688470
rect 119180 688230 119420 688470
rect 119510 688230 119750 688470
rect 119840 688230 120080 688470
rect 120190 688230 120430 688470
rect 120520 688230 120760 688470
rect 120850 688230 121090 688470
rect 121180 688230 121420 688470
rect 121530 688230 121770 688470
rect 110810 687900 111050 688140
rect 111140 687900 111380 688140
rect 111470 687900 111710 688140
rect 111800 687900 112040 688140
rect 112150 687900 112390 688140
rect 112480 687900 112720 688140
rect 112810 687900 113050 688140
rect 113140 687900 113380 688140
rect 113490 687900 113730 688140
rect 113820 687900 114060 688140
rect 114150 687900 114390 688140
rect 114480 687900 114720 688140
rect 114830 687900 115070 688140
rect 115160 687900 115400 688140
rect 115490 687900 115730 688140
rect 115820 687900 116060 688140
rect 116170 687900 116410 688140
rect 116500 687900 116740 688140
rect 116830 687900 117070 688140
rect 117160 687900 117400 688140
rect 117510 687900 117750 688140
rect 117840 687900 118080 688140
rect 118170 687900 118410 688140
rect 118500 687900 118740 688140
rect 118850 687900 119090 688140
rect 119180 687900 119420 688140
rect 119510 687900 119750 688140
rect 119840 687900 120080 688140
rect 120190 687900 120430 688140
rect 120520 687900 120760 688140
rect 120850 687900 121090 688140
rect 121180 687900 121420 688140
rect 121530 687900 121770 688140
rect 110810 687550 111050 687790
rect 111140 687550 111380 687790
rect 111470 687550 111710 687790
rect 111800 687550 112040 687790
rect 112150 687550 112390 687790
rect 112480 687550 112720 687790
rect 112810 687550 113050 687790
rect 113140 687550 113380 687790
rect 113490 687550 113730 687790
rect 113820 687550 114060 687790
rect 114150 687550 114390 687790
rect 114480 687550 114720 687790
rect 114830 687550 115070 687790
rect 115160 687550 115400 687790
rect 115490 687550 115730 687790
rect 115820 687550 116060 687790
rect 116170 687550 116410 687790
rect 116500 687550 116740 687790
rect 116830 687550 117070 687790
rect 117160 687550 117400 687790
rect 117510 687550 117750 687790
rect 117840 687550 118080 687790
rect 118170 687550 118410 687790
rect 118500 687550 118740 687790
rect 118850 687550 119090 687790
rect 119180 687550 119420 687790
rect 119510 687550 119750 687790
rect 119840 687550 120080 687790
rect 120190 687550 120430 687790
rect 120520 687550 120760 687790
rect 120850 687550 121090 687790
rect 121180 687550 121420 687790
rect 121530 687550 121770 687790
rect 110810 687220 111050 687460
rect 111140 687220 111380 687460
rect 111470 687220 111710 687460
rect 111800 687220 112040 687460
rect 112150 687220 112390 687460
rect 112480 687220 112720 687460
rect 112810 687220 113050 687460
rect 113140 687220 113380 687460
rect 113490 687220 113730 687460
rect 113820 687220 114060 687460
rect 114150 687220 114390 687460
rect 114480 687220 114720 687460
rect 114830 687220 115070 687460
rect 115160 687220 115400 687460
rect 115490 687220 115730 687460
rect 115820 687220 116060 687460
rect 116170 687220 116410 687460
rect 116500 687220 116740 687460
rect 116830 687220 117070 687460
rect 117160 687220 117400 687460
rect 117510 687220 117750 687460
rect 117840 687220 118080 687460
rect 118170 687220 118410 687460
rect 118500 687220 118740 687460
rect 118850 687220 119090 687460
rect 119180 687220 119420 687460
rect 119510 687220 119750 687460
rect 119840 687220 120080 687460
rect 120190 687220 120430 687460
rect 120520 687220 120760 687460
rect 120850 687220 121090 687460
rect 121180 687220 121420 687460
rect 121530 687220 121770 687460
rect 110810 686890 111050 687130
rect 111140 686890 111380 687130
rect 111470 686890 111710 687130
rect 111800 686890 112040 687130
rect 112150 686890 112390 687130
rect 112480 686890 112720 687130
rect 112810 686890 113050 687130
rect 113140 686890 113380 687130
rect 113490 686890 113730 687130
rect 113820 686890 114060 687130
rect 114150 686890 114390 687130
rect 114480 686890 114720 687130
rect 114830 686890 115070 687130
rect 115160 686890 115400 687130
rect 115490 686890 115730 687130
rect 115820 686890 116060 687130
rect 116170 686890 116410 687130
rect 116500 686890 116740 687130
rect 116830 686890 117070 687130
rect 117160 686890 117400 687130
rect 117510 686890 117750 687130
rect 117840 686890 118080 687130
rect 118170 686890 118410 687130
rect 118500 686890 118740 687130
rect 118850 686890 119090 687130
rect 119180 686890 119420 687130
rect 119510 686890 119750 687130
rect 119840 686890 120080 687130
rect 120190 686890 120430 687130
rect 120520 686890 120760 687130
rect 120850 686890 121090 687130
rect 121180 686890 121420 687130
rect 121530 686890 121770 687130
rect 110810 686560 111050 686800
rect 111140 686560 111380 686800
rect 111470 686560 111710 686800
rect 111800 686560 112040 686800
rect 112150 686560 112390 686800
rect 112480 686560 112720 686800
rect 112810 686560 113050 686800
rect 113140 686560 113380 686800
rect 113490 686560 113730 686800
rect 113820 686560 114060 686800
rect 114150 686560 114390 686800
rect 114480 686560 114720 686800
rect 114830 686560 115070 686800
rect 115160 686560 115400 686800
rect 115490 686560 115730 686800
rect 115820 686560 116060 686800
rect 116170 686560 116410 686800
rect 116500 686560 116740 686800
rect 116830 686560 117070 686800
rect 117160 686560 117400 686800
rect 117510 686560 117750 686800
rect 117840 686560 118080 686800
rect 118170 686560 118410 686800
rect 118500 686560 118740 686800
rect 118850 686560 119090 686800
rect 119180 686560 119420 686800
rect 119510 686560 119750 686800
rect 119840 686560 120080 686800
rect 120190 686560 120430 686800
rect 120520 686560 120760 686800
rect 120850 686560 121090 686800
rect 121180 686560 121420 686800
rect 121530 686560 121770 686800
rect 110810 686210 111050 686450
rect 111140 686210 111380 686450
rect 111470 686210 111710 686450
rect 111800 686210 112040 686450
rect 112150 686210 112390 686450
rect 112480 686210 112720 686450
rect 112810 686210 113050 686450
rect 113140 686210 113380 686450
rect 113490 686210 113730 686450
rect 113820 686210 114060 686450
rect 114150 686210 114390 686450
rect 114480 686210 114720 686450
rect 114830 686210 115070 686450
rect 115160 686210 115400 686450
rect 115490 686210 115730 686450
rect 115820 686210 116060 686450
rect 116170 686210 116410 686450
rect 116500 686210 116740 686450
rect 116830 686210 117070 686450
rect 117160 686210 117400 686450
rect 117510 686210 117750 686450
rect 117840 686210 118080 686450
rect 118170 686210 118410 686450
rect 118500 686210 118740 686450
rect 118850 686210 119090 686450
rect 119180 686210 119420 686450
rect 119510 686210 119750 686450
rect 119840 686210 120080 686450
rect 120190 686210 120430 686450
rect 120520 686210 120760 686450
rect 120850 686210 121090 686450
rect 121180 686210 121420 686450
rect 121530 686210 121770 686450
rect 110810 685880 111050 686120
rect 111140 685880 111380 686120
rect 111470 685880 111710 686120
rect 111800 685880 112040 686120
rect 112150 685880 112390 686120
rect 112480 685880 112720 686120
rect 112810 685880 113050 686120
rect 113140 685880 113380 686120
rect 113490 685880 113730 686120
rect 113820 685880 114060 686120
rect 114150 685880 114390 686120
rect 114480 685880 114720 686120
rect 114830 685880 115070 686120
rect 115160 685880 115400 686120
rect 115490 685880 115730 686120
rect 115820 685880 116060 686120
rect 116170 685880 116410 686120
rect 116500 685880 116740 686120
rect 116830 685880 117070 686120
rect 117160 685880 117400 686120
rect 117510 685880 117750 686120
rect 117840 685880 118080 686120
rect 118170 685880 118410 686120
rect 118500 685880 118740 686120
rect 118850 685880 119090 686120
rect 119180 685880 119420 686120
rect 119510 685880 119750 686120
rect 119840 685880 120080 686120
rect 120190 685880 120430 686120
rect 120520 685880 120760 686120
rect 120850 685880 121090 686120
rect 121180 685880 121420 686120
rect 121530 685880 121770 686120
rect 110810 685550 111050 685790
rect 111140 685550 111380 685790
rect 111470 685550 111710 685790
rect 111800 685550 112040 685790
rect 112150 685550 112390 685790
rect 112480 685550 112720 685790
rect 112810 685550 113050 685790
rect 113140 685550 113380 685790
rect 113490 685550 113730 685790
rect 113820 685550 114060 685790
rect 114150 685550 114390 685790
rect 114480 685550 114720 685790
rect 114830 685550 115070 685790
rect 115160 685550 115400 685790
rect 115490 685550 115730 685790
rect 115820 685550 116060 685790
rect 116170 685550 116410 685790
rect 116500 685550 116740 685790
rect 116830 685550 117070 685790
rect 117160 685550 117400 685790
rect 117510 685550 117750 685790
rect 117840 685550 118080 685790
rect 118170 685550 118410 685790
rect 118500 685550 118740 685790
rect 118850 685550 119090 685790
rect 119180 685550 119420 685790
rect 119510 685550 119750 685790
rect 119840 685550 120080 685790
rect 120190 685550 120430 685790
rect 120520 685550 120760 685790
rect 120850 685550 121090 685790
rect 121180 685550 121420 685790
rect 121530 685550 121770 685790
rect 110810 685220 111050 685460
rect 111140 685220 111380 685460
rect 111470 685220 111710 685460
rect 111800 685220 112040 685460
rect 112150 685220 112390 685460
rect 112480 685220 112720 685460
rect 112810 685220 113050 685460
rect 113140 685220 113380 685460
rect 113490 685220 113730 685460
rect 113820 685220 114060 685460
rect 114150 685220 114390 685460
rect 114480 685220 114720 685460
rect 114830 685220 115070 685460
rect 115160 685220 115400 685460
rect 115490 685220 115730 685460
rect 115820 685220 116060 685460
rect 116170 685220 116410 685460
rect 116500 685220 116740 685460
rect 116830 685220 117070 685460
rect 117160 685220 117400 685460
rect 117510 685220 117750 685460
rect 117840 685220 118080 685460
rect 118170 685220 118410 685460
rect 118500 685220 118740 685460
rect 118850 685220 119090 685460
rect 119180 685220 119420 685460
rect 119510 685220 119750 685460
rect 119840 685220 120080 685460
rect 120190 685220 120430 685460
rect 120520 685220 120760 685460
rect 120850 685220 121090 685460
rect 121180 685220 121420 685460
rect 121530 685220 121770 685460
rect 110810 684870 111050 685110
rect 111140 684870 111380 685110
rect 111470 684870 111710 685110
rect 111800 684870 112040 685110
rect 112150 684870 112390 685110
rect 112480 684870 112720 685110
rect 112810 684870 113050 685110
rect 113140 684870 113380 685110
rect 113490 684870 113730 685110
rect 113820 684870 114060 685110
rect 114150 684870 114390 685110
rect 114480 684870 114720 685110
rect 114830 684870 115070 685110
rect 115160 684870 115400 685110
rect 115490 684870 115730 685110
rect 115820 684870 116060 685110
rect 116170 684870 116410 685110
rect 116500 684870 116740 685110
rect 116830 684870 117070 685110
rect 117160 684870 117400 685110
rect 117510 684870 117750 685110
rect 117840 684870 118080 685110
rect 118170 684870 118410 685110
rect 118500 684870 118740 685110
rect 118850 684870 119090 685110
rect 119180 684870 119420 685110
rect 119510 684870 119750 685110
rect 119840 684870 120080 685110
rect 120190 684870 120430 685110
rect 120520 684870 120760 685110
rect 120850 684870 121090 685110
rect 121180 684870 121420 685110
rect 121530 684870 121770 685110
rect 110810 684540 111050 684780
rect 111140 684540 111380 684780
rect 111470 684540 111710 684780
rect 111800 684540 112040 684780
rect 112150 684540 112390 684780
rect 112480 684540 112720 684780
rect 112810 684540 113050 684780
rect 113140 684540 113380 684780
rect 113490 684540 113730 684780
rect 113820 684540 114060 684780
rect 114150 684540 114390 684780
rect 114480 684540 114720 684780
rect 114830 684540 115070 684780
rect 115160 684540 115400 684780
rect 115490 684540 115730 684780
rect 115820 684540 116060 684780
rect 116170 684540 116410 684780
rect 116500 684540 116740 684780
rect 116830 684540 117070 684780
rect 117160 684540 117400 684780
rect 117510 684540 117750 684780
rect 117840 684540 118080 684780
rect 118170 684540 118410 684780
rect 118500 684540 118740 684780
rect 118850 684540 119090 684780
rect 119180 684540 119420 684780
rect 119510 684540 119750 684780
rect 119840 684540 120080 684780
rect 120190 684540 120430 684780
rect 120520 684540 120760 684780
rect 120850 684540 121090 684780
rect 121180 684540 121420 684780
rect 121530 684540 121770 684780
rect 110810 684210 111050 684450
rect 111140 684210 111380 684450
rect 111470 684210 111710 684450
rect 111800 684210 112040 684450
rect 112150 684210 112390 684450
rect 112480 684210 112720 684450
rect 112810 684210 113050 684450
rect 113140 684210 113380 684450
rect 113490 684210 113730 684450
rect 113820 684210 114060 684450
rect 114150 684210 114390 684450
rect 114480 684210 114720 684450
rect 114830 684210 115070 684450
rect 115160 684210 115400 684450
rect 115490 684210 115730 684450
rect 115820 684210 116060 684450
rect 116170 684210 116410 684450
rect 116500 684210 116740 684450
rect 116830 684210 117070 684450
rect 117160 684210 117400 684450
rect 117510 684210 117750 684450
rect 117840 684210 118080 684450
rect 118170 684210 118410 684450
rect 118500 684210 118740 684450
rect 118850 684210 119090 684450
rect 119180 684210 119420 684450
rect 119510 684210 119750 684450
rect 119840 684210 120080 684450
rect 120190 684210 120430 684450
rect 120520 684210 120760 684450
rect 120850 684210 121090 684450
rect 121180 684210 121420 684450
rect 121530 684210 121770 684450
rect 110810 683880 111050 684120
rect 111140 683880 111380 684120
rect 111470 683880 111710 684120
rect 111800 683880 112040 684120
rect 112150 683880 112390 684120
rect 112480 683880 112720 684120
rect 112810 683880 113050 684120
rect 113140 683880 113380 684120
rect 113490 683880 113730 684120
rect 113820 683880 114060 684120
rect 114150 683880 114390 684120
rect 114480 683880 114720 684120
rect 114830 683880 115070 684120
rect 115160 683880 115400 684120
rect 115490 683880 115730 684120
rect 115820 683880 116060 684120
rect 116170 683880 116410 684120
rect 116500 683880 116740 684120
rect 116830 683880 117070 684120
rect 117160 683880 117400 684120
rect 117510 683880 117750 684120
rect 117840 683880 118080 684120
rect 118170 683880 118410 684120
rect 118500 683880 118740 684120
rect 118850 683880 119090 684120
rect 119180 683880 119420 684120
rect 119510 683880 119750 684120
rect 119840 683880 120080 684120
rect 120190 683880 120430 684120
rect 120520 683880 120760 684120
rect 120850 683880 121090 684120
rect 121180 683880 121420 684120
rect 121530 683880 121770 684120
rect 122190 694600 122430 694840
rect 122520 694600 122760 694840
rect 122850 694600 123090 694840
rect 123180 694600 123420 694840
rect 123530 694600 123770 694840
rect 123860 694600 124100 694840
rect 124190 694600 124430 694840
rect 124520 694600 124760 694840
rect 124870 694600 125110 694840
rect 125200 694600 125440 694840
rect 125530 694600 125770 694840
rect 125860 694600 126100 694840
rect 126210 694600 126450 694840
rect 126540 694600 126780 694840
rect 126870 694600 127110 694840
rect 127200 694600 127440 694840
rect 127550 694600 127790 694840
rect 127880 694600 128120 694840
rect 128210 694600 128450 694840
rect 128540 694600 128780 694840
rect 128890 694600 129130 694840
rect 129220 694600 129460 694840
rect 129550 694600 129790 694840
rect 129880 694600 130120 694840
rect 130230 694600 130470 694840
rect 130560 694600 130800 694840
rect 130890 694600 131130 694840
rect 131220 694600 131460 694840
rect 131570 694600 131810 694840
rect 131900 694600 132140 694840
rect 132230 694600 132470 694840
rect 132560 694600 132800 694840
rect 132910 694600 133150 694840
rect 122190 694250 122430 694490
rect 122520 694250 122760 694490
rect 122850 694250 123090 694490
rect 123180 694250 123420 694490
rect 123530 694250 123770 694490
rect 123860 694250 124100 694490
rect 124190 694250 124430 694490
rect 124520 694250 124760 694490
rect 124870 694250 125110 694490
rect 125200 694250 125440 694490
rect 125530 694250 125770 694490
rect 125860 694250 126100 694490
rect 126210 694250 126450 694490
rect 126540 694250 126780 694490
rect 126870 694250 127110 694490
rect 127200 694250 127440 694490
rect 127550 694250 127790 694490
rect 127880 694250 128120 694490
rect 128210 694250 128450 694490
rect 128540 694250 128780 694490
rect 128890 694250 129130 694490
rect 129220 694250 129460 694490
rect 129550 694250 129790 694490
rect 129880 694250 130120 694490
rect 130230 694250 130470 694490
rect 130560 694250 130800 694490
rect 130890 694250 131130 694490
rect 131220 694250 131460 694490
rect 131570 694250 131810 694490
rect 131900 694250 132140 694490
rect 132230 694250 132470 694490
rect 132560 694250 132800 694490
rect 132910 694250 133150 694490
rect 122190 693920 122430 694160
rect 122520 693920 122760 694160
rect 122850 693920 123090 694160
rect 123180 693920 123420 694160
rect 123530 693920 123770 694160
rect 123860 693920 124100 694160
rect 124190 693920 124430 694160
rect 124520 693920 124760 694160
rect 124870 693920 125110 694160
rect 125200 693920 125440 694160
rect 125530 693920 125770 694160
rect 125860 693920 126100 694160
rect 126210 693920 126450 694160
rect 126540 693920 126780 694160
rect 126870 693920 127110 694160
rect 127200 693920 127440 694160
rect 127550 693920 127790 694160
rect 127880 693920 128120 694160
rect 128210 693920 128450 694160
rect 128540 693920 128780 694160
rect 128890 693920 129130 694160
rect 129220 693920 129460 694160
rect 129550 693920 129790 694160
rect 129880 693920 130120 694160
rect 130230 693920 130470 694160
rect 130560 693920 130800 694160
rect 130890 693920 131130 694160
rect 131220 693920 131460 694160
rect 131570 693920 131810 694160
rect 131900 693920 132140 694160
rect 132230 693920 132470 694160
rect 132560 693920 132800 694160
rect 132910 693920 133150 694160
rect 122190 693590 122430 693830
rect 122520 693590 122760 693830
rect 122850 693590 123090 693830
rect 123180 693590 123420 693830
rect 123530 693590 123770 693830
rect 123860 693590 124100 693830
rect 124190 693590 124430 693830
rect 124520 693590 124760 693830
rect 124870 693590 125110 693830
rect 125200 693590 125440 693830
rect 125530 693590 125770 693830
rect 125860 693590 126100 693830
rect 126210 693590 126450 693830
rect 126540 693590 126780 693830
rect 126870 693590 127110 693830
rect 127200 693590 127440 693830
rect 127550 693590 127790 693830
rect 127880 693590 128120 693830
rect 128210 693590 128450 693830
rect 128540 693590 128780 693830
rect 128890 693590 129130 693830
rect 129220 693590 129460 693830
rect 129550 693590 129790 693830
rect 129880 693590 130120 693830
rect 130230 693590 130470 693830
rect 130560 693590 130800 693830
rect 130890 693590 131130 693830
rect 131220 693590 131460 693830
rect 131570 693590 131810 693830
rect 131900 693590 132140 693830
rect 132230 693590 132470 693830
rect 132560 693590 132800 693830
rect 132910 693590 133150 693830
rect 122190 693260 122430 693500
rect 122520 693260 122760 693500
rect 122850 693260 123090 693500
rect 123180 693260 123420 693500
rect 123530 693260 123770 693500
rect 123860 693260 124100 693500
rect 124190 693260 124430 693500
rect 124520 693260 124760 693500
rect 124870 693260 125110 693500
rect 125200 693260 125440 693500
rect 125530 693260 125770 693500
rect 125860 693260 126100 693500
rect 126210 693260 126450 693500
rect 126540 693260 126780 693500
rect 126870 693260 127110 693500
rect 127200 693260 127440 693500
rect 127550 693260 127790 693500
rect 127880 693260 128120 693500
rect 128210 693260 128450 693500
rect 128540 693260 128780 693500
rect 128890 693260 129130 693500
rect 129220 693260 129460 693500
rect 129550 693260 129790 693500
rect 129880 693260 130120 693500
rect 130230 693260 130470 693500
rect 130560 693260 130800 693500
rect 130890 693260 131130 693500
rect 131220 693260 131460 693500
rect 131570 693260 131810 693500
rect 131900 693260 132140 693500
rect 132230 693260 132470 693500
rect 132560 693260 132800 693500
rect 132910 693260 133150 693500
rect 122190 692910 122430 693150
rect 122520 692910 122760 693150
rect 122850 692910 123090 693150
rect 123180 692910 123420 693150
rect 123530 692910 123770 693150
rect 123860 692910 124100 693150
rect 124190 692910 124430 693150
rect 124520 692910 124760 693150
rect 124870 692910 125110 693150
rect 125200 692910 125440 693150
rect 125530 692910 125770 693150
rect 125860 692910 126100 693150
rect 126210 692910 126450 693150
rect 126540 692910 126780 693150
rect 126870 692910 127110 693150
rect 127200 692910 127440 693150
rect 127550 692910 127790 693150
rect 127880 692910 128120 693150
rect 128210 692910 128450 693150
rect 128540 692910 128780 693150
rect 128890 692910 129130 693150
rect 129220 692910 129460 693150
rect 129550 692910 129790 693150
rect 129880 692910 130120 693150
rect 130230 692910 130470 693150
rect 130560 692910 130800 693150
rect 130890 692910 131130 693150
rect 131220 692910 131460 693150
rect 131570 692910 131810 693150
rect 131900 692910 132140 693150
rect 132230 692910 132470 693150
rect 132560 692910 132800 693150
rect 132910 692910 133150 693150
rect 122190 692580 122430 692820
rect 122520 692580 122760 692820
rect 122850 692580 123090 692820
rect 123180 692580 123420 692820
rect 123530 692580 123770 692820
rect 123860 692580 124100 692820
rect 124190 692580 124430 692820
rect 124520 692580 124760 692820
rect 124870 692580 125110 692820
rect 125200 692580 125440 692820
rect 125530 692580 125770 692820
rect 125860 692580 126100 692820
rect 126210 692580 126450 692820
rect 126540 692580 126780 692820
rect 126870 692580 127110 692820
rect 127200 692580 127440 692820
rect 127550 692580 127790 692820
rect 127880 692580 128120 692820
rect 128210 692580 128450 692820
rect 128540 692580 128780 692820
rect 128890 692580 129130 692820
rect 129220 692580 129460 692820
rect 129550 692580 129790 692820
rect 129880 692580 130120 692820
rect 130230 692580 130470 692820
rect 130560 692580 130800 692820
rect 130890 692580 131130 692820
rect 131220 692580 131460 692820
rect 131570 692580 131810 692820
rect 131900 692580 132140 692820
rect 132230 692580 132470 692820
rect 132560 692580 132800 692820
rect 132910 692580 133150 692820
rect 122190 692250 122430 692490
rect 122520 692250 122760 692490
rect 122850 692250 123090 692490
rect 123180 692250 123420 692490
rect 123530 692250 123770 692490
rect 123860 692250 124100 692490
rect 124190 692250 124430 692490
rect 124520 692250 124760 692490
rect 124870 692250 125110 692490
rect 125200 692250 125440 692490
rect 125530 692250 125770 692490
rect 125860 692250 126100 692490
rect 126210 692250 126450 692490
rect 126540 692250 126780 692490
rect 126870 692250 127110 692490
rect 127200 692250 127440 692490
rect 127550 692250 127790 692490
rect 127880 692250 128120 692490
rect 128210 692250 128450 692490
rect 128540 692250 128780 692490
rect 128890 692250 129130 692490
rect 129220 692250 129460 692490
rect 129550 692250 129790 692490
rect 129880 692250 130120 692490
rect 130230 692250 130470 692490
rect 130560 692250 130800 692490
rect 130890 692250 131130 692490
rect 131220 692250 131460 692490
rect 131570 692250 131810 692490
rect 131900 692250 132140 692490
rect 132230 692250 132470 692490
rect 132560 692250 132800 692490
rect 132910 692250 133150 692490
rect 122190 691920 122430 692160
rect 122520 691920 122760 692160
rect 122850 691920 123090 692160
rect 123180 691920 123420 692160
rect 123530 691920 123770 692160
rect 123860 691920 124100 692160
rect 124190 691920 124430 692160
rect 124520 691920 124760 692160
rect 124870 691920 125110 692160
rect 125200 691920 125440 692160
rect 125530 691920 125770 692160
rect 125860 691920 126100 692160
rect 126210 691920 126450 692160
rect 126540 691920 126780 692160
rect 126870 691920 127110 692160
rect 127200 691920 127440 692160
rect 127550 691920 127790 692160
rect 127880 691920 128120 692160
rect 128210 691920 128450 692160
rect 128540 691920 128780 692160
rect 128890 691920 129130 692160
rect 129220 691920 129460 692160
rect 129550 691920 129790 692160
rect 129880 691920 130120 692160
rect 130230 691920 130470 692160
rect 130560 691920 130800 692160
rect 130890 691920 131130 692160
rect 131220 691920 131460 692160
rect 131570 691920 131810 692160
rect 131900 691920 132140 692160
rect 132230 691920 132470 692160
rect 132560 691920 132800 692160
rect 132910 691920 133150 692160
rect 122190 691570 122430 691810
rect 122520 691570 122760 691810
rect 122850 691570 123090 691810
rect 123180 691570 123420 691810
rect 123530 691570 123770 691810
rect 123860 691570 124100 691810
rect 124190 691570 124430 691810
rect 124520 691570 124760 691810
rect 124870 691570 125110 691810
rect 125200 691570 125440 691810
rect 125530 691570 125770 691810
rect 125860 691570 126100 691810
rect 126210 691570 126450 691810
rect 126540 691570 126780 691810
rect 126870 691570 127110 691810
rect 127200 691570 127440 691810
rect 127550 691570 127790 691810
rect 127880 691570 128120 691810
rect 128210 691570 128450 691810
rect 128540 691570 128780 691810
rect 128890 691570 129130 691810
rect 129220 691570 129460 691810
rect 129550 691570 129790 691810
rect 129880 691570 130120 691810
rect 130230 691570 130470 691810
rect 130560 691570 130800 691810
rect 130890 691570 131130 691810
rect 131220 691570 131460 691810
rect 131570 691570 131810 691810
rect 131900 691570 132140 691810
rect 132230 691570 132470 691810
rect 132560 691570 132800 691810
rect 132910 691570 133150 691810
rect 122190 691240 122430 691480
rect 122520 691240 122760 691480
rect 122850 691240 123090 691480
rect 123180 691240 123420 691480
rect 123530 691240 123770 691480
rect 123860 691240 124100 691480
rect 124190 691240 124430 691480
rect 124520 691240 124760 691480
rect 124870 691240 125110 691480
rect 125200 691240 125440 691480
rect 125530 691240 125770 691480
rect 125860 691240 126100 691480
rect 126210 691240 126450 691480
rect 126540 691240 126780 691480
rect 126870 691240 127110 691480
rect 127200 691240 127440 691480
rect 127550 691240 127790 691480
rect 127880 691240 128120 691480
rect 128210 691240 128450 691480
rect 128540 691240 128780 691480
rect 128890 691240 129130 691480
rect 129220 691240 129460 691480
rect 129550 691240 129790 691480
rect 129880 691240 130120 691480
rect 130230 691240 130470 691480
rect 130560 691240 130800 691480
rect 130890 691240 131130 691480
rect 131220 691240 131460 691480
rect 131570 691240 131810 691480
rect 131900 691240 132140 691480
rect 132230 691240 132470 691480
rect 132560 691240 132800 691480
rect 132910 691240 133150 691480
rect 122190 690910 122430 691150
rect 122520 690910 122760 691150
rect 122850 690910 123090 691150
rect 123180 690910 123420 691150
rect 123530 690910 123770 691150
rect 123860 690910 124100 691150
rect 124190 690910 124430 691150
rect 124520 690910 124760 691150
rect 124870 690910 125110 691150
rect 125200 690910 125440 691150
rect 125530 690910 125770 691150
rect 125860 690910 126100 691150
rect 126210 690910 126450 691150
rect 126540 690910 126780 691150
rect 126870 690910 127110 691150
rect 127200 690910 127440 691150
rect 127550 690910 127790 691150
rect 127880 690910 128120 691150
rect 128210 690910 128450 691150
rect 128540 690910 128780 691150
rect 128890 690910 129130 691150
rect 129220 690910 129460 691150
rect 129550 690910 129790 691150
rect 129880 690910 130120 691150
rect 130230 690910 130470 691150
rect 130560 690910 130800 691150
rect 130890 690910 131130 691150
rect 131220 690910 131460 691150
rect 131570 690910 131810 691150
rect 131900 690910 132140 691150
rect 132230 690910 132470 691150
rect 132560 690910 132800 691150
rect 132910 690910 133150 691150
rect 122190 690580 122430 690820
rect 122520 690580 122760 690820
rect 122850 690580 123090 690820
rect 123180 690580 123420 690820
rect 123530 690580 123770 690820
rect 123860 690580 124100 690820
rect 124190 690580 124430 690820
rect 124520 690580 124760 690820
rect 124870 690580 125110 690820
rect 125200 690580 125440 690820
rect 125530 690580 125770 690820
rect 125860 690580 126100 690820
rect 126210 690580 126450 690820
rect 126540 690580 126780 690820
rect 126870 690580 127110 690820
rect 127200 690580 127440 690820
rect 127550 690580 127790 690820
rect 127880 690580 128120 690820
rect 128210 690580 128450 690820
rect 128540 690580 128780 690820
rect 128890 690580 129130 690820
rect 129220 690580 129460 690820
rect 129550 690580 129790 690820
rect 129880 690580 130120 690820
rect 130230 690580 130470 690820
rect 130560 690580 130800 690820
rect 130890 690580 131130 690820
rect 131220 690580 131460 690820
rect 131570 690580 131810 690820
rect 131900 690580 132140 690820
rect 132230 690580 132470 690820
rect 132560 690580 132800 690820
rect 132910 690580 133150 690820
rect 122190 690230 122430 690470
rect 122520 690230 122760 690470
rect 122850 690230 123090 690470
rect 123180 690230 123420 690470
rect 123530 690230 123770 690470
rect 123860 690230 124100 690470
rect 124190 690230 124430 690470
rect 124520 690230 124760 690470
rect 124870 690230 125110 690470
rect 125200 690230 125440 690470
rect 125530 690230 125770 690470
rect 125860 690230 126100 690470
rect 126210 690230 126450 690470
rect 126540 690230 126780 690470
rect 126870 690230 127110 690470
rect 127200 690230 127440 690470
rect 127550 690230 127790 690470
rect 127880 690230 128120 690470
rect 128210 690230 128450 690470
rect 128540 690230 128780 690470
rect 128890 690230 129130 690470
rect 129220 690230 129460 690470
rect 129550 690230 129790 690470
rect 129880 690230 130120 690470
rect 130230 690230 130470 690470
rect 130560 690230 130800 690470
rect 130890 690230 131130 690470
rect 131220 690230 131460 690470
rect 131570 690230 131810 690470
rect 131900 690230 132140 690470
rect 132230 690230 132470 690470
rect 132560 690230 132800 690470
rect 132910 690230 133150 690470
rect 122190 689900 122430 690140
rect 122520 689900 122760 690140
rect 122850 689900 123090 690140
rect 123180 689900 123420 690140
rect 123530 689900 123770 690140
rect 123860 689900 124100 690140
rect 124190 689900 124430 690140
rect 124520 689900 124760 690140
rect 124870 689900 125110 690140
rect 125200 689900 125440 690140
rect 125530 689900 125770 690140
rect 125860 689900 126100 690140
rect 126210 689900 126450 690140
rect 126540 689900 126780 690140
rect 126870 689900 127110 690140
rect 127200 689900 127440 690140
rect 127550 689900 127790 690140
rect 127880 689900 128120 690140
rect 128210 689900 128450 690140
rect 128540 689900 128780 690140
rect 128890 689900 129130 690140
rect 129220 689900 129460 690140
rect 129550 689900 129790 690140
rect 129880 689900 130120 690140
rect 130230 689900 130470 690140
rect 130560 689900 130800 690140
rect 130890 689900 131130 690140
rect 131220 689900 131460 690140
rect 131570 689900 131810 690140
rect 131900 689900 132140 690140
rect 132230 689900 132470 690140
rect 132560 689900 132800 690140
rect 132910 689900 133150 690140
rect 122190 689570 122430 689810
rect 122520 689570 122760 689810
rect 122850 689570 123090 689810
rect 123180 689570 123420 689810
rect 123530 689570 123770 689810
rect 123860 689570 124100 689810
rect 124190 689570 124430 689810
rect 124520 689570 124760 689810
rect 124870 689570 125110 689810
rect 125200 689570 125440 689810
rect 125530 689570 125770 689810
rect 125860 689570 126100 689810
rect 126210 689570 126450 689810
rect 126540 689570 126780 689810
rect 126870 689570 127110 689810
rect 127200 689570 127440 689810
rect 127550 689570 127790 689810
rect 127880 689570 128120 689810
rect 128210 689570 128450 689810
rect 128540 689570 128780 689810
rect 128890 689570 129130 689810
rect 129220 689570 129460 689810
rect 129550 689570 129790 689810
rect 129880 689570 130120 689810
rect 130230 689570 130470 689810
rect 130560 689570 130800 689810
rect 130890 689570 131130 689810
rect 131220 689570 131460 689810
rect 131570 689570 131810 689810
rect 131900 689570 132140 689810
rect 132230 689570 132470 689810
rect 132560 689570 132800 689810
rect 132910 689570 133150 689810
rect 122190 689240 122430 689480
rect 122520 689240 122760 689480
rect 122850 689240 123090 689480
rect 123180 689240 123420 689480
rect 123530 689240 123770 689480
rect 123860 689240 124100 689480
rect 124190 689240 124430 689480
rect 124520 689240 124760 689480
rect 124870 689240 125110 689480
rect 125200 689240 125440 689480
rect 125530 689240 125770 689480
rect 125860 689240 126100 689480
rect 126210 689240 126450 689480
rect 126540 689240 126780 689480
rect 126870 689240 127110 689480
rect 127200 689240 127440 689480
rect 127550 689240 127790 689480
rect 127880 689240 128120 689480
rect 128210 689240 128450 689480
rect 128540 689240 128780 689480
rect 128890 689240 129130 689480
rect 129220 689240 129460 689480
rect 129550 689240 129790 689480
rect 129880 689240 130120 689480
rect 130230 689240 130470 689480
rect 130560 689240 130800 689480
rect 130890 689240 131130 689480
rect 131220 689240 131460 689480
rect 131570 689240 131810 689480
rect 131900 689240 132140 689480
rect 132230 689240 132470 689480
rect 132560 689240 132800 689480
rect 132910 689240 133150 689480
rect 122190 688890 122430 689130
rect 122520 688890 122760 689130
rect 122850 688890 123090 689130
rect 123180 688890 123420 689130
rect 123530 688890 123770 689130
rect 123860 688890 124100 689130
rect 124190 688890 124430 689130
rect 124520 688890 124760 689130
rect 124870 688890 125110 689130
rect 125200 688890 125440 689130
rect 125530 688890 125770 689130
rect 125860 688890 126100 689130
rect 126210 688890 126450 689130
rect 126540 688890 126780 689130
rect 126870 688890 127110 689130
rect 127200 688890 127440 689130
rect 127550 688890 127790 689130
rect 127880 688890 128120 689130
rect 128210 688890 128450 689130
rect 128540 688890 128780 689130
rect 128890 688890 129130 689130
rect 129220 688890 129460 689130
rect 129550 688890 129790 689130
rect 129880 688890 130120 689130
rect 130230 688890 130470 689130
rect 130560 688890 130800 689130
rect 130890 688890 131130 689130
rect 131220 688890 131460 689130
rect 131570 688890 131810 689130
rect 131900 688890 132140 689130
rect 132230 688890 132470 689130
rect 132560 688890 132800 689130
rect 132910 688890 133150 689130
rect 122190 688560 122430 688800
rect 122520 688560 122760 688800
rect 122850 688560 123090 688800
rect 123180 688560 123420 688800
rect 123530 688560 123770 688800
rect 123860 688560 124100 688800
rect 124190 688560 124430 688800
rect 124520 688560 124760 688800
rect 124870 688560 125110 688800
rect 125200 688560 125440 688800
rect 125530 688560 125770 688800
rect 125860 688560 126100 688800
rect 126210 688560 126450 688800
rect 126540 688560 126780 688800
rect 126870 688560 127110 688800
rect 127200 688560 127440 688800
rect 127550 688560 127790 688800
rect 127880 688560 128120 688800
rect 128210 688560 128450 688800
rect 128540 688560 128780 688800
rect 128890 688560 129130 688800
rect 129220 688560 129460 688800
rect 129550 688560 129790 688800
rect 129880 688560 130120 688800
rect 130230 688560 130470 688800
rect 130560 688560 130800 688800
rect 130890 688560 131130 688800
rect 131220 688560 131460 688800
rect 131570 688560 131810 688800
rect 131900 688560 132140 688800
rect 132230 688560 132470 688800
rect 132560 688560 132800 688800
rect 132910 688560 133150 688800
rect 122190 688230 122430 688470
rect 122520 688230 122760 688470
rect 122850 688230 123090 688470
rect 123180 688230 123420 688470
rect 123530 688230 123770 688470
rect 123860 688230 124100 688470
rect 124190 688230 124430 688470
rect 124520 688230 124760 688470
rect 124870 688230 125110 688470
rect 125200 688230 125440 688470
rect 125530 688230 125770 688470
rect 125860 688230 126100 688470
rect 126210 688230 126450 688470
rect 126540 688230 126780 688470
rect 126870 688230 127110 688470
rect 127200 688230 127440 688470
rect 127550 688230 127790 688470
rect 127880 688230 128120 688470
rect 128210 688230 128450 688470
rect 128540 688230 128780 688470
rect 128890 688230 129130 688470
rect 129220 688230 129460 688470
rect 129550 688230 129790 688470
rect 129880 688230 130120 688470
rect 130230 688230 130470 688470
rect 130560 688230 130800 688470
rect 130890 688230 131130 688470
rect 131220 688230 131460 688470
rect 131570 688230 131810 688470
rect 131900 688230 132140 688470
rect 132230 688230 132470 688470
rect 132560 688230 132800 688470
rect 132910 688230 133150 688470
rect 122190 687900 122430 688140
rect 122520 687900 122760 688140
rect 122850 687900 123090 688140
rect 123180 687900 123420 688140
rect 123530 687900 123770 688140
rect 123860 687900 124100 688140
rect 124190 687900 124430 688140
rect 124520 687900 124760 688140
rect 124870 687900 125110 688140
rect 125200 687900 125440 688140
rect 125530 687900 125770 688140
rect 125860 687900 126100 688140
rect 126210 687900 126450 688140
rect 126540 687900 126780 688140
rect 126870 687900 127110 688140
rect 127200 687900 127440 688140
rect 127550 687900 127790 688140
rect 127880 687900 128120 688140
rect 128210 687900 128450 688140
rect 128540 687900 128780 688140
rect 128890 687900 129130 688140
rect 129220 687900 129460 688140
rect 129550 687900 129790 688140
rect 129880 687900 130120 688140
rect 130230 687900 130470 688140
rect 130560 687900 130800 688140
rect 130890 687900 131130 688140
rect 131220 687900 131460 688140
rect 131570 687900 131810 688140
rect 131900 687900 132140 688140
rect 132230 687900 132470 688140
rect 132560 687900 132800 688140
rect 132910 687900 133150 688140
rect 122190 687550 122430 687790
rect 122520 687550 122760 687790
rect 122850 687550 123090 687790
rect 123180 687550 123420 687790
rect 123530 687550 123770 687790
rect 123860 687550 124100 687790
rect 124190 687550 124430 687790
rect 124520 687550 124760 687790
rect 124870 687550 125110 687790
rect 125200 687550 125440 687790
rect 125530 687550 125770 687790
rect 125860 687550 126100 687790
rect 126210 687550 126450 687790
rect 126540 687550 126780 687790
rect 126870 687550 127110 687790
rect 127200 687550 127440 687790
rect 127550 687550 127790 687790
rect 127880 687550 128120 687790
rect 128210 687550 128450 687790
rect 128540 687550 128780 687790
rect 128890 687550 129130 687790
rect 129220 687550 129460 687790
rect 129550 687550 129790 687790
rect 129880 687550 130120 687790
rect 130230 687550 130470 687790
rect 130560 687550 130800 687790
rect 130890 687550 131130 687790
rect 131220 687550 131460 687790
rect 131570 687550 131810 687790
rect 131900 687550 132140 687790
rect 132230 687550 132470 687790
rect 132560 687550 132800 687790
rect 132910 687550 133150 687790
rect 122190 687220 122430 687460
rect 122520 687220 122760 687460
rect 122850 687220 123090 687460
rect 123180 687220 123420 687460
rect 123530 687220 123770 687460
rect 123860 687220 124100 687460
rect 124190 687220 124430 687460
rect 124520 687220 124760 687460
rect 124870 687220 125110 687460
rect 125200 687220 125440 687460
rect 125530 687220 125770 687460
rect 125860 687220 126100 687460
rect 126210 687220 126450 687460
rect 126540 687220 126780 687460
rect 126870 687220 127110 687460
rect 127200 687220 127440 687460
rect 127550 687220 127790 687460
rect 127880 687220 128120 687460
rect 128210 687220 128450 687460
rect 128540 687220 128780 687460
rect 128890 687220 129130 687460
rect 129220 687220 129460 687460
rect 129550 687220 129790 687460
rect 129880 687220 130120 687460
rect 130230 687220 130470 687460
rect 130560 687220 130800 687460
rect 130890 687220 131130 687460
rect 131220 687220 131460 687460
rect 131570 687220 131810 687460
rect 131900 687220 132140 687460
rect 132230 687220 132470 687460
rect 132560 687220 132800 687460
rect 132910 687220 133150 687460
rect 122190 686890 122430 687130
rect 122520 686890 122760 687130
rect 122850 686890 123090 687130
rect 123180 686890 123420 687130
rect 123530 686890 123770 687130
rect 123860 686890 124100 687130
rect 124190 686890 124430 687130
rect 124520 686890 124760 687130
rect 124870 686890 125110 687130
rect 125200 686890 125440 687130
rect 125530 686890 125770 687130
rect 125860 686890 126100 687130
rect 126210 686890 126450 687130
rect 126540 686890 126780 687130
rect 126870 686890 127110 687130
rect 127200 686890 127440 687130
rect 127550 686890 127790 687130
rect 127880 686890 128120 687130
rect 128210 686890 128450 687130
rect 128540 686890 128780 687130
rect 128890 686890 129130 687130
rect 129220 686890 129460 687130
rect 129550 686890 129790 687130
rect 129880 686890 130120 687130
rect 130230 686890 130470 687130
rect 130560 686890 130800 687130
rect 130890 686890 131130 687130
rect 131220 686890 131460 687130
rect 131570 686890 131810 687130
rect 131900 686890 132140 687130
rect 132230 686890 132470 687130
rect 132560 686890 132800 687130
rect 132910 686890 133150 687130
rect 122190 686560 122430 686800
rect 122520 686560 122760 686800
rect 122850 686560 123090 686800
rect 123180 686560 123420 686800
rect 123530 686560 123770 686800
rect 123860 686560 124100 686800
rect 124190 686560 124430 686800
rect 124520 686560 124760 686800
rect 124870 686560 125110 686800
rect 125200 686560 125440 686800
rect 125530 686560 125770 686800
rect 125860 686560 126100 686800
rect 126210 686560 126450 686800
rect 126540 686560 126780 686800
rect 126870 686560 127110 686800
rect 127200 686560 127440 686800
rect 127550 686560 127790 686800
rect 127880 686560 128120 686800
rect 128210 686560 128450 686800
rect 128540 686560 128780 686800
rect 128890 686560 129130 686800
rect 129220 686560 129460 686800
rect 129550 686560 129790 686800
rect 129880 686560 130120 686800
rect 130230 686560 130470 686800
rect 130560 686560 130800 686800
rect 130890 686560 131130 686800
rect 131220 686560 131460 686800
rect 131570 686560 131810 686800
rect 131900 686560 132140 686800
rect 132230 686560 132470 686800
rect 132560 686560 132800 686800
rect 132910 686560 133150 686800
rect 122190 686210 122430 686450
rect 122520 686210 122760 686450
rect 122850 686210 123090 686450
rect 123180 686210 123420 686450
rect 123530 686210 123770 686450
rect 123860 686210 124100 686450
rect 124190 686210 124430 686450
rect 124520 686210 124760 686450
rect 124870 686210 125110 686450
rect 125200 686210 125440 686450
rect 125530 686210 125770 686450
rect 125860 686210 126100 686450
rect 126210 686210 126450 686450
rect 126540 686210 126780 686450
rect 126870 686210 127110 686450
rect 127200 686210 127440 686450
rect 127550 686210 127790 686450
rect 127880 686210 128120 686450
rect 128210 686210 128450 686450
rect 128540 686210 128780 686450
rect 128890 686210 129130 686450
rect 129220 686210 129460 686450
rect 129550 686210 129790 686450
rect 129880 686210 130120 686450
rect 130230 686210 130470 686450
rect 130560 686210 130800 686450
rect 130890 686210 131130 686450
rect 131220 686210 131460 686450
rect 131570 686210 131810 686450
rect 131900 686210 132140 686450
rect 132230 686210 132470 686450
rect 132560 686210 132800 686450
rect 132910 686210 133150 686450
rect 122190 685880 122430 686120
rect 122520 685880 122760 686120
rect 122850 685880 123090 686120
rect 123180 685880 123420 686120
rect 123530 685880 123770 686120
rect 123860 685880 124100 686120
rect 124190 685880 124430 686120
rect 124520 685880 124760 686120
rect 124870 685880 125110 686120
rect 125200 685880 125440 686120
rect 125530 685880 125770 686120
rect 125860 685880 126100 686120
rect 126210 685880 126450 686120
rect 126540 685880 126780 686120
rect 126870 685880 127110 686120
rect 127200 685880 127440 686120
rect 127550 685880 127790 686120
rect 127880 685880 128120 686120
rect 128210 685880 128450 686120
rect 128540 685880 128780 686120
rect 128890 685880 129130 686120
rect 129220 685880 129460 686120
rect 129550 685880 129790 686120
rect 129880 685880 130120 686120
rect 130230 685880 130470 686120
rect 130560 685880 130800 686120
rect 130890 685880 131130 686120
rect 131220 685880 131460 686120
rect 131570 685880 131810 686120
rect 131900 685880 132140 686120
rect 132230 685880 132470 686120
rect 132560 685880 132800 686120
rect 132910 685880 133150 686120
rect 122190 685550 122430 685790
rect 122520 685550 122760 685790
rect 122850 685550 123090 685790
rect 123180 685550 123420 685790
rect 123530 685550 123770 685790
rect 123860 685550 124100 685790
rect 124190 685550 124430 685790
rect 124520 685550 124760 685790
rect 124870 685550 125110 685790
rect 125200 685550 125440 685790
rect 125530 685550 125770 685790
rect 125860 685550 126100 685790
rect 126210 685550 126450 685790
rect 126540 685550 126780 685790
rect 126870 685550 127110 685790
rect 127200 685550 127440 685790
rect 127550 685550 127790 685790
rect 127880 685550 128120 685790
rect 128210 685550 128450 685790
rect 128540 685550 128780 685790
rect 128890 685550 129130 685790
rect 129220 685550 129460 685790
rect 129550 685550 129790 685790
rect 129880 685550 130120 685790
rect 130230 685550 130470 685790
rect 130560 685550 130800 685790
rect 130890 685550 131130 685790
rect 131220 685550 131460 685790
rect 131570 685550 131810 685790
rect 131900 685550 132140 685790
rect 132230 685550 132470 685790
rect 132560 685550 132800 685790
rect 132910 685550 133150 685790
rect 122190 685220 122430 685460
rect 122520 685220 122760 685460
rect 122850 685220 123090 685460
rect 123180 685220 123420 685460
rect 123530 685220 123770 685460
rect 123860 685220 124100 685460
rect 124190 685220 124430 685460
rect 124520 685220 124760 685460
rect 124870 685220 125110 685460
rect 125200 685220 125440 685460
rect 125530 685220 125770 685460
rect 125860 685220 126100 685460
rect 126210 685220 126450 685460
rect 126540 685220 126780 685460
rect 126870 685220 127110 685460
rect 127200 685220 127440 685460
rect 127550 685220 127790 685460
rect 127880 685220 128120 685460
rect 128210 685220 128450 685460
rect 128540 685220 128780 685460
rect 128890 685220 129130 685460
rect 129220 685220 129460 685460
rect 129550 685220 129790 685460
rect 129880 685220 130120 685460
rect 130230 685220 130470 685460
rect 130560 685220 130800 685460
rect 130890 685220 131130 685460
rect 131220 685220 131460 685460
rect 131570 685220 131810 685460
rect 131900 685220 132140 685460
rect 132230 685220 132470 685460
rect 132560 685220 132800 685460
rect 132910 685220 133150 685460
rect 122190 684870 122430 685110
rect 122520 684870 122760 685110
rect 122850 684870 123090 685110
rect 123180 684870 123420 685110
rect 123530 684870 123770 685110
rect 123860 684870 124100 685110
rect 124190 684870 124430 685110
rect 124520 684870 124760 685110
rect 124870 684870 125110 685110
rect 125200 684870 125440 685110
rect 125530 684870 125770 685110
rect 125860 684870 126100 685110
rect 126210 684870 126450 685110
rect 126540 684870 126780 685110
rect 126870 684870 127110 685110
rect 127200 684870 127440 685110
rect 127550 684870 127790 685110
rect 127880 684870 128120 685110
rect 128210 684870 128450 685110
rect 128540 684870 128780 685110
rect 128890 684870 129130 685110
rect 129220 684870 129460 685110
rect 129550 684870 129790 685110
rect 129880 684870 130120 685110
rect 130230 684870 130470 685110
rect 130560 684870 130800 685110
rect 130890 684870 131130 685110
rect 131220 684870 131460 685110
rect 131570 684870 131810 685110
rect 131900 684870 132140 685110
rect 132230 684870 132470 685110
rect 132560 684870 132800 685110
rect 132910 684870 133150 685110
rect 122190 684540 122430 684780
rect 122520 684540 122760 684780
rect 122850 684540 123090 684780
rect 123180 684540 123420 684780
rect 123530 684540 123770 684780
rect 123860 684540 124100 684780
rect 124190 684540 124430 684780
rect 124520 684540 124760 684780
rect 124870 684540 125110 684780
rect 125200 684540 125440 684780
rect 125530 684540 125770 684780
rect 125860 684540 126100 684780
rect 126210 684540 126450 684780
rect 126540 684540 126780 684780
rect 126870 684540 127110 684780
rect 127200 684540 127440 684780
rect 127550 684540 127790 684780
rect 127880 684540 128120 684780
rect 128210 684540 128450 684780
rect 128540 684540 128780 684780
rect 128890 684540 129130 684780
rect 129220 684540 129460 684780
rect 129550 684540 129790 684780
rect 129880 684540 130120 684780
rect 130230 684540 130470 684780
rect 130560 684540 130800 684780
rect 130890 684540 131130 684780
rect 131220 684540 131460 684780
rect 131570 684540 131810 684780
rect 131900 684540 132140 684780
rect 132230 684540 132470 684780
rect 132560 684540 132800 684780
rect 132910 684540 133150 684780
rect 122190 684210 122430 684450
rect 122520 684210 122760 684450
rect 122850 684210 123090 684450
rect 123180 684210 123420 684450
rect 123530 684210 123770 684450
rect 123860 684210 124100 684450
rect 124190 684210 124430 684450
rect 124520 684210 124760 684450
rect 124870 684210 125110 684450
rect 125200 684210 125440 684450
rect 125530 684210 125770 684450
rect 125860 684210 126100 684450
rect 126210 684210 126450 684450
rect 126540 684210 126780 684450
rect 126870 684210 127110 684450
rect 127200 684210 127440 684450
rect 127550 684210 127790 684450
rect 127880 684210 128120 684450
rect 128210 684210 128450 684450
rect 128540 684210 128780 684450
rect 128890 684210 129130 684450
rect 129220 684210 129460 684450
rect 129550 684210 129790 684450
rect 129880 684210 130120 684450
rect 130230 684210 130470 684450
rect 130560 684210 130800 684450
rect 130890 684210 131130 684450
rect 131220 684210 131460 684450
rect 131570 684210 131810 684450
rect 131900 684210 132140 684450
rect 132230 684210 132470 684450
rect 132560 684210 132800 684450
rect 132910 684210 133150 684450
rect 122190 683880 122430 684120
rect 122520 683880 122760 684120
rect 122850 683880 123090 684120
rect 123180 683880 123420 684120
rect 123530 683880 123770 684120
rect 123860 683880 124100 684120
rect 124190 683880 124430 684120
rect 124520 683880 124760 684120
rect 124870 683880 125110 684120
rect 125200 683880 125440 684120
rect 125530 683880 125770 684120
rect 125860 683880 126100 684120
rect 126210 683880 126450 684120
rect 126540 683880 126780 684120
rect 126870 683880 127110 684120
rect 127200 683880 127440 684120
rect 127550 683880 127790 684120
rect 127880 683880 128120 684120
rect 128210 683880 128450 684120
rect 128540 683880 128780 684120
rect 128890 683880 129130 684120
rect 129220 683880 129460 684120
rect 129550 683880 129790 684120
rect 129880 683880 130120 684120
rect 130230 683880 130470 684120
rect 130560 683880 130800 684120
rect 130890 683880 131130 684120
rect 131220 683880 131460 684120
rect 131570 683880 131810 684120
rect 131900 683880 132140 684120
rect 132230 683880 132470 684120
rect 132560 683880 132800 684120
rect 132910 683880 133150 684120
rect 133570 694600 133810 694840
rect 133900 694600 134140 694840
rect 134230 694600 134470 694840
rect 134560 694600 134800 694840
rect 134910 694600 135150 694840
rect 135240 694600 135480 694840
rect 135570 694600 135810 694840
rect 135900 694600 136140 694840
rect 136250 694600 136490 694840
rect 136580 694600 136820 694840
rect 136910 694600 137150 694840
rect 137240 694600 137480 694840
rect 137590 694600 137830 694840
rect 137920 694600 138160 694840
rect 138250 694600 138490 694840
rect 138580 694600 138820 694840
rect 138930 694600 139170 694840
rect 139260 694600 139500 694840
rect 139590 694600 139830 694840
rect 139920 694600 140160 694840
rect 140270 694600 140510 694840
rect 140600 694600 140840 694840
rect 140930 694600 141170 694840
rect 141260 694600 141500 694840
rect 141610 694600 141850 694840
rect 141940 694600 142180 694840
rect 142270 694600 142510 694840
rect 142600 694600 142840 694840
rect 142950 694600 143190 694840
rect 143280 694600 143520 694840
rect 143610 694600 143850 694840
rect 143940 694600 144180 694840
rect 144290 694600 144530 694840
rect 133570 694250 133810 694490
rect 133900 694250 134140 694490
rect 134230 694250 134470 694490
rect 134560 694250 134800 694490
rect 134910 694250 135150 694490
rect 135240 694250 135480 694490
rect 135570 694250 135810 694490
rect 135900 694250 136140 694490
rect 136250 694250 136490 694490
rect 136580 694250 136820 694490
rect 136910 694250 137150 694490
rect 137240 694250 137480 694490
rect 137590 694250 137830 694490
rect 137920 694250 138160 694490
rect 138250 694250 138490 694490
rect 138580 694250 138820 694490
rect 138930 694250 139170 694490
rect 139260 694250 139500 694490
rect 139590 694250 139830 694490
rect 139920 694250 140160 694490
rect 140270 694250 140510 694490
rect 140600 694250 140840 694490
rect 140930 694250 141170 694490
rect 141260 694250 141500 694490
rect 141610 694250 141850 694490
rect 141940 694250 142180 694490
rect 142270 694250 142510 694490
rect 142600 694250 142840 694490
rect 142950 694250 143190 694490
rect 143280 694250 143520 694490
rect 143610 694250 143850 694490
rect 143940 694250 144180 694490
rect 144290 694250 144530 694490
rect 133570 693920 133810 694160
rect 133900 693920 134140 694160
rect 134230 693920 134470 694160
rect 134560 693920 134800 694160
rect 134910 693920 135150 694160
rect 135240 693920 135480 694160
rect 135570 693920 135810 694160
rect 135900 693920 136140 694160
rect 136250 693920 136490 694160
rect 136580 693920 136820 694160
rect 136910 693920 137150 694160
rect 137240 693920 137480 694160
rect 137590 693920 137830 694160
rect 137920 693920 138160 694160
rect 138250 693920 138490 694160
rect 138580 693920 138820 694160
rect 138930 693920 139170 694160
rect 139260 693920 139500 694160
rect 139590 693920 139830 694160
rect 139920 693920 140160 694160
rect 140270 693920 140510 694160
rect 140600 693920 140840 694160
rect 140930 693920 141170 694160
rect 141260 693920 141500 694160
rect 141610 693920 141850 694160
rect 141940 693920 142180 694160
rect 142270 693920 142510 694160
rect 142600 693920 142840 694160
rect 142950 693920 143190 694160
rect 143280 693920 143520 694160
rect 143610 693920 143850 694160
rect 143940 693920 144180 694160
rect 144290 693920 144530 694160
rect 133570 693590 133810 693830
rect 133900 693590 134140 693830
rect 134230 693590 134470 693830
rect 134560 693590 134800 693830
rect 134910 693590 135150 693830
rect 135240 693590 135480 693830
rect 135570 693590 135810 693830
rect 135900 693590 136140 693830
rect 136250 693590 136490 693830
rect 136580 693590 136820 693830
rect 136910 693590 137150 693830
rect 137240 693590 137480 693830
rect 137590 693590 137830 693830
rect 137920 693590 138160 693830
rect 138250 693590 138490 693830
rect 138580 693590 138820 693830
rect 138930 693590 139170 693830
rect 139260 693590 139500 693830
rect 139590 693590 139830 693830
rect 139920 693590 140160 693830
rect 140270 693590 140510 693830
rect 140600 693590 140840 693830
rect 140930 693590 141170 693830
rect 141260 693590 141500 693830
rect 141610 693590 141850 693830
rect 141940 693590 142180 693830
rect 142270 693590 142510 693830
rect 142600 693590 142840 693830
rect 142950 693590 143190 693830
rect 143280 693590 143520 693830
rect 143610 693590 143850 693830
rect 143940 693590 144180 693830
rect 144290 693590 144530 693830
rect 133570 693260 133810 693500
rect 133900 693260 134140 693500
rect 134230 693260 134470 693500
rect 134560 693260 134800 693500
rect 134910 693260 135150 693500
rect 135240 693260 135480 693500
rect 135570 693260 135810 693500
rect 135900 693260 136140 693500
rect 136250 693260 136490 693500
rect 136580 693260 136820 693500
rect 136910 693260 137150 693500
rect 137240 693260 137480 693500
rect 137590 693260 137830 693500
rect 137920 693260 138160 693500
rect 138250 693260 138490 693500
rect 138580 693260 138820 693500
rect 138930 693260 139170 693500
rect 139260 693260 139500 693500
rect 139590 693260 139830 693500
rect 139920 693260 140160 693500
rect 140270 693260 140510 693500
rect 140600 693260 140840 693500
rect 140930 693260 141170 693500
rect 141260 693260 141500 693500
rect 141610 693260 141850 693500
rect 141940 693260 142180 693500
rect 142270 693260 142510 693500
rect 142600 693260 142840 693500
rect 142950 693260 143190 693500
rect 143280 693260 143520 693500
rect 143610 693260 143850 693500
rect 143940 693260 144180 693500
rect 144290 693260 144530 693500
rect 133570 692910 133810 693150
rect 133900 692910 134140 693150
rect 134230 692910 134470 693150
rect 134560 692910 134800 693150
rect 134910 692910 135150 693150
rect 135240 692910 135480 693150
rect 135570 692910 135810 693150
rect 135900 692910 136140 693150
rect 136250 692910 136490 693150
rect 136580 692910 136820 693150
rect 136910 692910 137150 693150
rect 137240 692910 137480 693150
rect 137590 692910 137830 693150
rect 137920 692910 138160 693150
rect 138250 692910 138490 693150
rect 138580 692910 138820 693150
rect 138930 692910 139170 693150
rect 139260 692910 139500 693150
rect 139590 692910 139830 693150
rect 139920 692910 140160 693150
rect 140270 692910 140510 693150
rect 140600 692910 140840 693150
rect 140930 692910 141170 693150
rect 141260 692910 141500 693150
rect 141610 692910 141850 693150
rect 141940 692910 142180 693150
rect 142270 692910 142510 693150
rect 142600 692910 142840 693150
rect 142950 692910 143190 693150
rect 143280 692910 143520 693150
rect 143610 692910 143850 693150
rect 143940 692910 144180 693150
rect 144290 692910 144530 693150
rect 133570 692580 133810 692820
rect 133900 692580 134140 692820
rect 134230 692580 134470 692820
rect 134560 692580 134800 692820
rect 134910 692580 135150 692820
rect 135240 692580 135480 692820
rect 135570 692580 135810 692820
rect 135900 692580 136140 692820
rect 136250 692580 136490 692820
rect 136580 692580 136820 692820
rect 136910 692580 137150 692820
rect 137240 692580 137480 692820
rect 137590 692580 137830 692820
rect 137920 692580 138160 692820
rect 138250 692580 138490 692820
rect 138580 692580 138820 692820
rect 138930 692580 139170 692820
rect 139260 692580 139500 692820
rect 139590 692580 139830 692820
rect 139920 692580 140160 692820
rect 140270 692580 140510 692820
rect 140600 692580 140840 692820
rect 140930 692580 141170 692820
rect 141260 692580 141500 692820
rect 141610 692580 141850 692820
rect 141940 692580 142180 692820
rect 142270 692580 142510 692820
rect 142600 692580 142840 692820
rect 142950 692580 143190 692820
rect 143280 692580 143520 692820
rect 143610 692580 143850 692820
rect 143940 692580 144180 692820
rect 144290 692580 144530 692820
rect 133570 692250 133810 692490
rect 133900 692250 134140 692490
rect 134230 692250 134470 692490
rect 134560 692250 134800 692490
rect 134910 692250 135150 692490
rect 135240 692250 135480 692490
rect 135570 692250 135810 692490
rect 135900 692250 136140 692490
rect 136250 692250 136490 692490
rect 136580 692250 136820 692490
rect 136910 692250 137150 692490
rect 137240 692250 137480 692490
rect 137590 692250 137830 692490
rect 137920 692250 138160 692490
rect 138250 692250 138490 692490
rect 138580 692250 138820 692490
rect 138930 692250 139170 692490
rect 139260 692250 139500 692490
rect 139590 692250 139830 692490
rect 139920 692250 140160 692490
rect 140270 692250 140510 692490
rect 140600 692250 140840 692490
rect 140930 692250 141170 692490
rect 141260 692250 141500 692490
rect 141610 692250 141850 692490
rect 141940 692250 142180 692490
rect 142270 692250 142510 692490
rect 142600 692250 142840 692490
rect 142950 692250 143190 692490
rect 143280 692250 143520 692490
rect 143610 692250 143850 692490
rect 143940 692250 144180 692490
rect 144290 692250 144530 692490
rect 133570 691920 133810 692160
rect 133900 691920 134140 692160
rect 134230 691920 134470 692160
rect 134560 691920 134800 692160
rect 134910 691920 135150 692160
rect 135240 691920 135480 692160
rect 135570 691920 135810 692160
rect 135900 691920 136140 692160
rect 136250 691920 136490 692160
rect 136580 691920 136820 692160
rect 136910 691920 137150 692160
rect 137240 691920 137480 692160
rect 137590 691920 137830 692160
rect 137920 691920 138160 692160
rect 138250 691920 138490 692160
rect 138580 691920 138820 692160
rect 138930 691920 139170 692160
rect 139260 691920 139500 692160
rect 139590 691920 139830 692160
rect 139920 691920 140160 692160
rect 140270 691920 140510 692160
rect 140600 691920 140840 692160
rect 140930 691920 141170 692160
rect 141260 691920 141500 692160
rect 141610 691920 141850 692160
rect 141940 691920 142180 692160
rect 142270 691920 142510 692160
rect 142600 691920 142840 692160
rect 142950 691920 143190 692160
rect 143280 691920 143520 692160
rect 143610 691920 143850 692160
rect 143940 691920 144180 692160
rect 144290 691920 144530 692160
rect 133570 691570 133810 691810
rect 133900 691570 134140 691810
rect 134230 691570 134470 691810
rect 134560 691570 134800 691810
rect 134910 691570 135150 691810
rect 135240 691570 135480 691810
rect 135570 691570 135810 691810
rect 135900 691570 136140 691810
rect 136250 691570 136490 691810
rect 136580 691570 136820 691810
rect 136910 691570 137150 691810
rect 137240 691570 137480 691810
rect 137590 691570 137830 691810
rect 137920 691570 138160 691810
rect 138250 691570 138490 691810
rect 138580 691570 138820 691810
rect 138930 691570 139170 691810
rect 139260 691570 139500 691810
rect 139590 691570 139830 691810
rect 139920 691570 140160 691810
rect 140270 691570 140510 691810
rect 140600 691570 140840 691810
rect 140930 691570 141170 691810
rect 141260 691570 141500 691810
rect 141610 691570 141850 691810
rect 141940 691570 142180 691810
rect 142270 691570 142510 691810
rect 142600 691570 142840 691810
rect 142950 691570 143190 691810
rect 143280 691570 143520 691810
rect 143610 691570 143850 691810
rect 143940 691570 144180 691810
rect 144290 691570 144530 691810
rect 133570 691240 133810 691480
rect 133900 691240 134140 691480
rect 134230 691240 134470 691480
rect 134560 691240 134800 691480
rect 134910 691240 135150 691480
rect 135240 691240 135480 691480
rect 135570 691240 135810 691480
rect 135900 691240 136140 691480
rect 136250 691240 136490 691480
rect 136580 691240 136820 691480
rect 136910 691240 137150 691480
rect 137240 691240 137480 691480
rect 137590 691240 137830 691480
rect 137920 691240 138160 691480
rect 138250 691240 138490 691480
rect 138580 691240 138820 691480
rect 138930 691240 139170 691480
rect 139260 691240 139500 691480
rect 139590 691240 139830 691480
rect 139920 691240 140160 691480
rect 140270 691240 140510 691480
rect 140600 691240 140840 691480
rect 140930 691240 141170 691480
rect 141260 691240 141500 691480
rect 141610 691240 141850 691480
rect 141940 691240 142180 691480
rect 142270 691240 142510 691480
rect 142600 691240 142840 691480
rect 142950 691240 143190 691480
rect 143280 691240 143520 691480
rect 143610 691240 143850 691480
rect 143940 691240 144180 691480
rect 144290 691240 144530 691480
rect 133570 690910 133810 691150
rect 133900 690910 134140 691150
rect 134230 690910 134470 691150
rect 134560 690910 134800 691150
rect 134910 690910 135150 691150
rect 135240 690910 135480 691150
rect 135570 690910 135810 691150
rect 135900 690910 136140 691150
rect 136250 690910 136490 691150
rect 136580 690910 136820 691150
rect 136910 690910 137150 691150
rect 137240 690910 137480 691150
rect 137590 690910 137830 691150
rect 137920 690910 138160 691150
rect 138250 690910 138490 691150
rect 138580 690910 138820 691150
rect 138930 690910 139170 691150
rect 139260 690910 139500 691150
rect 139590 690910 139830 691150
rect 139920 690910 140160 691150
rect 140270 690910 140510 691150
rect 140600 690910 140840 691150
rect 140930 690910 141170 691150
rect 141260 690910 141500 691150
rect 141610 690910 141850 691150
rect 141940 690910 142180 691150
rect 142270 690910 142510 691150
rect 142600 690910 142840 691150
rect 142950 690910 143190 691150
rect 143280 690910 143520 691150
rect 143610 690910 143850 691150
rect 143940 690910 144180 691150
rect 144290 690910 144530 691150
rect 133570 690580 133810 690820
rect 133900 690580 134140 690820
rect 134230 690580 134470 690820
rect 134560 690580 134800 690820
rect 134910 690580 135150 690820
rect 135240 690580 135480 690820
rect 135570 690580 135810 690820
rect 135900 690580 136140 690820
rect 136250 690580 136490 690820
rect 136580 690580 136820 690820
rect 136910 690580 137150 690820
rect 137240 690580 137480 690820
rect 137590 690580 137830 690820
rect 137920 690580 138160 690820
rect 138250 690580 138490 690820
rect 138580 690580 138820 690820
rect 138930 690580 139170 690820
rect 139260 690580 139500 690820
rect 139590 690580 139830 690820
rect 139920 690580 140160 690820
rect 140270 690580 140510 690820
rect 140600 690580 140840 690820
rect 140930 690580 141170 690820
rect 141260 690580 141500 690820
rect 141610 690580 141850 690820
rect 141940 690580 142180 690820
rect 142270 690580 142510 690820
rect 142600 690580 142840 690820
rect 142950 690580 143190 690820
rect 143280 690580 143520 690820
rect 143610 690580 143850 690820
rect 143940 690580 144180 690820
rect 144290 690580 144530 690820
rect 133570 690230 133810 690470
rect 133900 690230 134140 690470
rect 134230 690230 134470 690470
rect 134560 690230 134800 690470
rect 134910 690230 135150 690470
rect 135240 690230 135480 690470
rect 135570 690230 135810 690470
rect 135900 690230 136140 690470
rect 136250 690230 136490 690470
rect 136580 690230 136820 690470
rect 136910 690230 137150 690470
rect 137240 690230 137480 690470
rect 137590 690230 137830 690470
rect 137920 690230 138160 690470
rect 138250 690230 138490 690470
rect 138580 690230 138820 690470
rect 138930 690230 139170 690470
rect 139260 690230 139500 690470
rect 139590 690230 139830 690470
rect 139920 690230 140160 690470
rect 140270 690230 140510 690470
rect 140600 690230 140840 690470
rect 140930 690230 141170 690470
rect 141260 690230 141500 690470
rect 141610 690230 141850 690470
rect 141940 690230 142180 690470
rect 142270 690230 142510 690470
rect 142600 690230 142840 690470
rect 142950 690230 143190 690470
rect 143280 690230 143520 690470
rect 143610 690230 143850 690470
rect 143940 690230 144180 690470
rect 144290 690230 144530 690470
rect 133570 689900 133810 690140
rect 133900 689900 134140 690140
rect 134230 689900 134470 690140
rect 134560 689900 134800 690140
rect 134910 689900 135150 690140
rect 135240 689900 135480 690140
rect 135570 689900 135810 690140
rect 135900 689900 136140 690140
rect 136250 689900 136490 690140
rect 136580 689900 136820 690140
rect 136910 689900 137150 690140
rect 137240 689900 137480 690140
rect 137590 689900 137830 690140
rect 137920 689900 138160 690140
rect 138250 689900 138490 690140
rect 138580 689900 138820 690140
rect 138930 689900 139170 690140
rect 139260 689900 139500 690140
rect 139590 689900 139830 690140
rect 139920 689900 140160 690140
rect 140270 689900 140510 690140
rect 140600 689900 140840 690140
rect 140930 689900 141170 690140
rect 141260 689900 141500 690140
rect 141610 689900 141850 690140
rect 141940 689900 142180 690140
rect 142270 689900 142510 690140
rect 142600 689900 142840 690140
rect 142950 689900 143190 690140
rect 143280 689900 143520 690140
rect 143610 689900 143850 690140
rect 143940 689900 144180 690140
rect 144290 689900 144530 690140
rect 133570 689570 133810 689810
rect 133900 689570 134140 689810
rect 134230 689570 134470 689810
rect 134560 689570 134800 689810
rect 134910 689570 135150 689810
rect 135240 689570 135480 689810
rect 135570 689570 135810 689810
rect 135900 689570 136140 689810
rect 136250 689570 136490 689810
rect 136580 689570 136820 689810
rect 136910 689570 137150 689810
rect 137240 689570 137480 689810
rect 137590 689570 137830 689810
rect 137920 689570 138160 689810
rect 138250 689570 138490 689810
rect 138580 689570 138820 689810
rect 138930 689570 139170 689810
rect 139260 689570 139500 689810
rect 139590 689570 139830 689810
rect 139920 689570 140160 689810
rect 140270 689570 140510 689810
rect 140600 689570 140840 689810
rect 140930 689570 141170 689810
rect 141260 689570 141500 689810
rect 141610 689570 141850 689810
rect 141940 689570 142180 689810
rect 142270 689570 142510 689810
rect 142600 689570 142840 689810
rect 142950 689570 143190 689810
rect 143280 689570 143520 689810
rect 143610 689570 143850 689810
rect 143940 689570 144180 689810
rect 144290 689570 144530 689810
rect 133570 689240 133810 689480
rect 133900 689240 134140 689480
rect 134230 689240 134470 689480
rect 134560 689240 134800 689480
rect 134910 689240 135150 689480
rect 135240 689240 135480 689480
rect 135570 689240 135810 689480
rect 135900 689240 136140 689480
rect 136250 689240 136490 689480
rect 136580 689240 136820 689480
rect 136910 689240 137150 689480
rect 137240 689240 137480 689480
rect 137590 689240 137830 689480
rect 137920 689240 138160 689480
rect 138250 689240 138490 689480
rect 138580 689240 138820 689480
rect 138930 689240 139170 689480
rect 139260 689240 139500 689480
rect 139590 689240 139830 689480
rect 139920 689240 140160 689480
rect 140270 689240 140510 689480
rect 140600 689240 140840 689480
rect 140930 689240 141170 689480
rect 141260 689240 141500 689480
rect 141610 689240 141850 689480
rect 141940 689240 142180 689480
rect 142270 689240 142510 689480
rect 142600 689240 142840 689480
rect 142950 689240 143190 689480
rect 143280 689240 143520 689480
rect 143610 689240 143850 689480
rect 143940 689240 144180 689480
rect 144290 689240 144530 689480
rect 133570 688890 133810 689130
rect 133900 688890 134140 689130
rect 134230 688890 134470 689130
rect 134560 688890 134800 689130
rect 134910 688890 135150 689130
rect 135240 688890 135480 689130
rect 135570 688890 135810 689130
rect 135900 688890 136140 689130
rect 136250 688890 136490 689130
rect 136580 688890 136820 689130
rect 136910 688890 137150 689130
rect 137240 688890 137480 689130
rect 137590 688890 137830 689130
rect 137920 688890 138160 689130
rect 138250 688890 138490 689130
rect 138580 688890 138820 689130
rect 138930 688890 139170 689130
rect 139260 688890 139500 689130
rect 139590 688890 139830 689130
rect 139920 688890 140160 689130
rect 140270 688890 140510 689130
rect 140600 688890 140840 689130
rect 140930 688890 141170 689130
rect 141260 688890 141500 689130
rect 141610 688890 141850 689130
rect 141940 688890 142180 689130
rect 142270 688890 142510 689130
rect 142600 688890 142840 689130
rect 142950 688890 143190 689130
rect 143280 688890 143520 689130
rect 143610 688890 143850 689130
rect 143940 688890 144180 689130
rect 144290 688890 144530 689130
rect 133570 688560 133810 688800
rect 133900 688560 134140 688800
rect 134230 688560 134470 688800
rect 134560 688560 134800 688800
rect 134910 688560 135150 688800
rect 135240 688560 135480 688800
rect 135570 688560 135810 688800
rect 135900 688560 136140 688800
rect 136250 688560 136490 688800
rect 136580 688560 136820 688800
rect 136910 688560 137150 688800
rect 137240 688560 137480 688800
rect 137590 688560 137830 688800
rect 137920 688560 138160 688800
rect 138250 688560 138490 688800
rect 138580 688560 138820 688800
rect 138930 688560 139170 688800
rect 139260 688560 139500 688800
rect 139590 688560 139830 688800
rect 139920 688560 140160 688800
rect 140270 688560 140510 688800
rect 140600 688560 140840 688800
rect 140930 688560 141170 688800
rect 141260 688560 141500 688800
rect 141610 688560 141850 688800
rect 141940 688560 142180 688800
rect 142270 688560 142510 688800
rect 142600 688560 142840 688800
rect 142950 688560 143190 688800
rect 143280 688560 143520 688800
rect 143610 688560 143850 688800
rect 143940 688560 144180 688800
rect 144290 688560 144530 688800
rect 133570 688230 133810 688470
rect 133900 688230 134140 688470
rect 134230 688230 134470 688470
rect 134560 688230 134800 688470
rect 134910 688230 135150 688470
rect 135240 688230 135480 688470
rect 135570 688230 135810 688470
rect 135900 688230 136140 688470
rect 136250 688230 136490 688470
rect 136580 688230 136820 688470
rect 136910 688230 137150 688470
rect 137240 688230 137480 688470
rect 137590 688230 137830 688470
rect 137920 688230 138160 688470
rect 138250 688230 138490 688470
rect 138580 688230 138820 688470
rect 138930 688230 139170 688470
rect 139260 688230 139500 688470
rect 139590 688230 139830 688470
rect 139920 688230 140160 688470
rect 140270 688230 140510 688470
rect 140600 688230 140840 688470
rect 140930 688230 141170 688470
rect 141260 688230 141500 688470
rect 141610 688230 141850 688470
rect 141940 688230 142180 688470
rect 142270 688230 142510 688470
rect 142600 688230 142840 688470
rect 142950 688230 143190 688470
rect 143280 688230 143520 688470
rect 143610 688230 143850 688470
rect 143940 688230 144180 688470
rect 144290 688230 144530 688470
rect 133570 687900 133810 688140
rect 133900 687900 134140 688140
rect 134230 687900 134470 688140
rect 134560 687900 134800 688140
rect 134910 687900 135150 688140
rect 135240 687900 135480 688140
rect 135570 687900 135810 688140
rect 135900 687900 136140 688140
rect 136250 687900 136490 688140
rect 136580 687900 136820 688140
rect 136910 687900 137150 688140
rect 137240 687900 137480 688140
rect 137590 687900 137830 688140
rect 137920 687900 138160 688140
rect 138250 687900 138490 688140
rect 138580 687900 138820 688140
rect 138930 687900 139170 688140
rect 139260 687900 139500 688140
rect 139590 687900 139830 688140
rect 139920 687900 140160 688140
rect 140270 687900 140510 688140
rect 140600 687900 140840 688140
rect 140930 687900 141170 688140
rect 141260 687900 141500 688140
rect 141610 687900 141850 688140
rect 141940 687900 142180 688140
rect 142270 687900 142510 688140
rect 142600 687900 142840 688140
rect 142950 687900 143190 688140
rect 143280 687900 143520 688140
rect 143610 687900 143850 688140
rect 143940 687900 144180 688140
rect 144290 687900 144530 688140
rect 133570 687550 133810 687790
rect 133900 687550 134140 687790
rect 134230 687550 134470 687790
rect 134560 687550 134800 687790
rect 134910 687550 135150 687790
rect 135240 687550 135480 687790
rect 135570 687550 135810 687790
rect 135900 687550 136140 687790
rect 136250 687550 136490 687790
rect 136580 687550 136820 687790
rect 136910 687550 137150 687790
rect 137240 687550 137480 687790
rect 137590 687550 137830 687790
rect 137920 687550 138160 687790
rect 138250 687550 138490 687790
rect 138580 687550 138820 687790
rect 138930 687550 139170 687790
rect 139260 687550 139500 687790
rect 139590 687550 139830 687790
rect 139920 687550 140160 687790
rect 140270 687550 140510 687790
rect 140600 687550 140840 687790
rect 140930 687550 141170 687790
rect 141260 687550 141500 687790
rect 141610 687550 141850 687790
rect 141940 687550 142180 687790
rect 142270 687550 142510 687790
rect 142600 687550 142840 687790
rect 142950 687550 143190 687790
rect 143280 687550 143520 687790
rect 143610 687550 143850 687790
rect 143940 687550 144180 687790
rect 144290 687550 144530 687790
rect 133570 687220 133810 687460
rect 133900 687220 134140 687460
rect 134230 687220 134470 687460
rect 134560 687220 134800 687460
rect 134910 687220 135150 687460
rect 135240 687220 135480 687460
rect 135570 687220 135810 687460
rect 135900 687220 136140 687460
rect 136250 687220 136490 687460
rect 136580 687220 136820 687460
rect 136910 687220 137150 687460
rect 137240 687220 137480 687460
rect 137590 687220 137830 687460
rect 137920 687220 138160 687460
rect 138250 687220 138490 687460
rect 138580 687220 138820 687460
rect 138930 687220 139170 687460
rect 139260 687220 139500 687460
rect 139590 687220 139830 687460
rect 139920 687220 140160 687460
rect 140270 687220 140510 687460
rect 140600 687220 140840 687460
rect 140930 687220 141170 687460
rect 141260 687220 141500 687460
rect 141610 687220 141850 687460
rect 141940 687220 142180 687460
rect 142270 687220 142510 687460
rect 142600 687220 142840 687460
rect 142950 687220 143190 687460
rect 143280 687220 143520 687460
rect 143610 687220 143850 687460
rect 143940 687220 144180 687460
rect 144290 687220 144530 687460
rect 133570 686890 133810 687130
rect 133900 686890 134140 687130
rect 134230 686890 134470 687130
rect 134560 686890 134800 687130
rect 134910 686890 135150 687130
rect 135240 686890 135480 687130
rect 135570 686890 135810 687130
rect 135900 686890 136140 687130
rect 136250 686890 136490 687130
rect 136580 686890 136820 687130
rect 136910 686890 137150 687130
rect 137240 686890 137480 687130
rect 137590 686890 137830 687130
rect 137920 686890 138160 687130
rect 138250 686890 138490 687130
rect 138580 686890 138820 687130
rect 138930 686890 139170 687130
rect 139260 686890 139500 687130
rect 139590 686890 139830 687130
rect 139920 686890 140160 687130
rect 140270 686890 140510 687130
rect 140600 686890 140840 687130
rect 140930 686890 141170 687130
rect 141260 686890 141500 687130
rect 141610 686890 141850 687130
rect 141940 686890 142180 687130
rect 142270 686890 142510 687130
rect 142600 686890 142840 687130
rect 142950 686890 143190 687130
rect 143280 686890 143520 687130
rect 143610 686890 143850 687130
rect 143940 686890 144180 687130
rect 144290 686890 144530 687130
rect 133570 686560 133810 686800
rect 133900 686560 134140 686800
rect 134230 686560 134470 686800
rect 134560 686560 134800 686800
rect 134910 686560 135150 686800
rect 135240 686560 135480 686800
rect 135570 686560 135810 686800
rect 135900 686560 136140 686800
rect 136250 686560 136490 686800
rect 136580 686560 136820 686800
rect 136910 686560 137150 686800
rect 137240 686560 137480 686800
rect 137590 686560 137830 686800
rect 137920 686560 138160 686800
rect 138250 686560 138490 686800
rect 138580 686560 138820 686800
rect 138930 686560 139170 686800
rect 139260 686560 139500 686800
rect 139590 686560 139830 686800
rect 139920 686560 140160 686800
rect 140270 686560 140510 686800
rect 140600 686560 140840 686800
rect 140930 686560 141170 686800
rect 141260 686560 141500 686800
rect 141610 686560 141850 686800
rect 141940 686560 142180 686800
rect 142270 686560 142510 686800
rect 142600 686560 142840 686800
rect 142950 686560 143190 686800
rect 143280 686560 143520 686800
rect 143610 686560 143850 686800
rect 143940 686560 144180 686800
rect 144290 686560 144530 686800
rect 133570 686210 133810 686450
rect 133900 686210 134140 686450
rect 134230 686210 134470 686450
rect 134560 686210 134800 686450
rect 134910 686210 135150 686450
rect 135240 686210 135480 686450
rect 135570 686210 135810 686450
rect 135900 686210 136140 686450
rect 136250 686210 136490 686450
rect 136580 686210 136820 686450
rect 136910 686210 137150 686450
rect 137240 686210 137480 686450
rect 137590 686210 137830 686450
rect 137920 686210 138160 686450
rect 138250 686210 138490 686450
rect 138580 686210 138820 686450
rect 138930 686210 139170 686450
rect 139260 686210 139500 686450
rect 139590 686210 139830 686450
rect 139920 686210 140160 686450
rect 140270 686210 140510 686450
rect 140600 686210 140840 686450
rect 140930 686210 141170 686450
rect 141260 686210 141500 686450
rect 141610 686210 141850 686450
rect 141940 686210 142180 686450
rect 142270 686210 142510 686450
rect 142600 686210 142840 686450
rect 142950 686210 143190 686450
rect 143280 686210 143520 686450
rect 143610 686210 143850 686450
rect 143940 686210 144180 686450
rect 144290 686210 144530 686450
rect 133570 685880 133810 686120
rect 133900 685880 134140 686120
rect 134230 685880 134470 686120
rect 134560 685880 134800 686120
rect 134910 685880 135150 686120
rect 135240 685880 135480 686120
rect 135570 685880 135810 686120
rect 135900 685880 136140 686120
rect 136250 685880 136490 686120
rect 136580 685880 136820 686120
rect 136910 685880 137150 686120
rect 137240 685880 137480 686120
rect 137590 685880 137830 686120
rect 137920 685880 138160 686120
rect 138250 685880 138490 686120
rect 138580 685880 138820 686120
rect 138930 685880 139170 686120
rect 139260 685880 139500 686120
rect 139590 685880 139830 686120
rect 139920 685880 140160 686120
rect 140270 685880 140510 686120
rect 140600 685880 140840 686120
rect 140930 685880 141170 686120
rect 141260 685880 141500 686120
rect 141610 685880 141850 686120
rect 141940 685880 142180 686120
rect 142270 685880 142510 686120
rect 142600 685880 142840 686120
rect 142950 685880 143190 686120
rect 143280 685880 143520 686120
rect 143610 685880 143850 686120
rect 143940 685880 144180 686120
rect 144290 685880 144530 686120
rect 133570 685550 133810 685790
rect 133900 685550 134140 685790
rect 134230 685550 134470 685790
rect 134560 685550 134800 685790
rect 134910 685550 135150 685790
rect 135240 685550 135480 685790
rect 135570 685550 135810 685790
rect 135900 685550 136140 685790
rect 136250 685550 136490 685790
rect 136580 685550 136820 685790
rect 136910 685550 137150 685790
rect 137240 685550 137480 685790
rect 137590 685550 137830 685790
rect 137920 685550 138160 685790
rect 138250 685550 138490 685790
rect 138580 685550 138820 685790
rect 138930 685550 139170 685790
rect 139260 685550 139500 685790
rect 139590 685550 139830 685790
rect 139920 685550 140160 685790
rect 140270 685550 140510 685790
rect 140600 685550 140840 685790
rect 140930 685550 141170 685790
rect 141260 685550 141500 685790
rect 141610 685550 141850 685790
rect 141940 685550 142180 685790
rect 142270 685550 142510 685790
rect 142600 685550 142840 685790
rect 142950 685550 143190 685790
rect 143280 685550 143520 685790
rect 143610 685550 143850 685790
rect 143940 685550 144180 685790
rect 144290 685550 144530 685790
rect 133570 685220 133810 685460
rect 133900 685220 134140 685460
rect 134230 685220 134470 685460
rect 134560 685220 134800 685460
rect 134910 685220 135150 685460
rect 135240 685220 135480 685460
rect 135570 685220 135810 685460
rect 135900 685220 136140 685460
rect 136250 685220 136490 685460
rect 136580 685220 136820 685460
rect 136910 685220 137150 685460
rect 137240 685220 137480 685460
rect 137590 685220 137830 685460
rect 137920 685220 138160 685460
rect 138250 685220 138490 685460
rect 138580 685220 138820 685460
rect 138930 685220 139170 685460
rect 139260 685220 139500 685460
rect 139590 685220 139830 685460
rect 139920 685220 140160 685460
rect 140270 685220 140510 685460
rect 140600 685220 140840 685460
rect 140930 685220 141170 685460
rect 141260 685220 141500 685460
rect 141610 685220 141850 685460
rect 141940 685220 142180 685460
rect 142270 685220 142510 685460
rect 142600 685220 142840 685460
rect 142950 685220 143190 685460
rect 143280 685220 143520 685460
rect 143610 685220 143850 685460
rect 143940 685220 144180 685460
rect 144290 685220 144530 685460
rect 133570 684870 133810 685110
rect 133900 684870 134140 685110
rect 134230 684870 134470 685110
rect 134560 684870 134800 685110
rect 134910 684870 135150 685110
rect 135240 684870 135480 685110
rect 135570 684870 135810 685110
rect 135900 684870 136140 685110
rect 136250 684870 136490 685110
rect 136580 684870 136820 685110
rect 136910 684870 137150 685110
rect 137240 684870 137480 685110
rect 137590 684870 137830 685110
rect 137920 684870 138160 685110
rect 138250 684870 138490 685110
rect 138580 684870 138820 685110
rect 138930 684870 139170 685110
rect 139260 684870 139500 685110
rect 139590 684870 139830 685110
rect 139920 684870 140160 685110
rect 140270 684870 140510 685110
rect 140600 684870 140840 685110
rect 140930 684870 141170 685110
rect 141260 684870 141500 685110
rect 141610 684870 141850 685110
rect 141940 684870 142180 685110
rect 142270 684870 142510 685110
rect 142600 684870 142840 685110
rect 142950 684870 143190 685110
rect 143280 684870 143520 685110
rect 143610 684870 143850 685110
rect 143940 684870 144180 685110
rect 144290 684870 144530 685110
rect 133570 684540 133810 684780
rect 133900 684540 134140 684780
rect 134230 684540 134470 684780
rect 134560 684540 134800 684780
rect 134910 684540 135150 684780
rect 135240 684540 135480 684780
rect 135570 684540 135810 684780
rect 135900 684540 136140 684780
rect 136250 684540 136490 684780
rect 136580 684540 136820 684780
rect 136910 684540 137150 684780
rect 137240 684540 137480 684780
rect 137590 684540 137830 684780
rect 137920 684540 138160 684780
rect 138250 684540 138490 684780
rect 138580 684540 138820 684780
rect 138930 684540 139170 684780
rect 139260 684540 139500 684780
rect 139590 684540 139830 684780
rect 139920 684540 140160 684780
rect 140270 684540 140510 684780
rect 140600 684540 140840 684780
rect 140930 684540 141170 684780
rect 141260 684540 141500 684780
rect 141610 684540 141850 684780
rect 141940 684540 142180 684780
rect 142270 684540 142510 684780
rect 142600 684540 142840 684780
rect 142950 684540 143190 684780
rect 143280 684540 143520 684780
rect 143610 684540 143850 684780
rect 143940 684540 144180 684780
rect 144290 684540 144530 684780
rect 133570 684210 133810 684450
rect 133900 684210 134140 684450
rect 134230 684210 134470 684450
rect 134560 684210 134800 684450
rect 134910 684210 135150 684450
rect 135240 684210 135480 684450
rect 135570 684210 135810 684450
rect 135900 684210 136140 684450
rect 136250 684210 136490 684450
rect 136580 684210 136820 684450
rect 136910 684210 137150 684450
rect 137240 684210 137480 684450
rect 137590 684210 137830 684450
rect 137920 684210 138160 684450
rect 138250 684210 138490 684450
rect 138580 684210 138820 684450
rect 138930 684210 139170 684450
rect 139260 684210 139500 684450
rect 139590 684210 139830 684450
rect 139920 684210 140160 684450
rect 140270 684210 140510 684450
rect 140600 684210 140840 684450
rect 140930 684210 141170 684450
rect 141260 684210 141500 684450
rect 141610 684210 141850 684450
rect 141940 684210 142180 684450
rect 142270 684210 142510 684450
rect 142600 684210 142840 684450
rect 142950 684210 143190 684450
rect 143280 684210 143520 684450
rect 143610 684210 143850 684450
rect 143940 684210 144180 684450
rect 144290 684210 144530 684450
rect 133570 683880 133810 684120
rect 133900 683880 134140 684120
rect 134230 683880 134470 684120
rect 134560 683880 134800 684120
rect 134910 683880 135150 684120
rect 135240 683880 135480 684120
rect 135570 683880 135810 684120
rect 135900 683880 136140 684120
rect 136250 683880 136490 684120
rect 136580 683880 136820 684120
rect 136910 683880 137150 684120
rect 137240 683880 137480 684120
rect 137590 683880 137830 684120
rect 137920 683880 138160 684120
rect 138250 683880 138490 684120
rect 138580 683880 138820 684120
rect 138930 683880 139170 684120
rect 139260 683880 139500 684120
rect 139590 683880 139830 684120
rect 139920 683880 140160 684120
rect 140270 683880 140510 684120
rect 140600 683880 140840 684120
rect 140930 683880 141170 684120
rect 141260 683880 141500 684120
rect 141610 683880 141850 684120
rect 141940 683880 142180 684120
rect 142270 683880 142510 684120
rect 142600 683880 142840 684120
rect 142950 683880 143190 684120
rect 143280 683880 143520 684120
rect 143610 683880 143850 684120
rect 143940 683880 144180 684120
rect 144290 683880 144530 684120
rect 144950 694600 145190 694840
rect 145280 694600 145520 694840
rect 145610 694600 145850 694840
rect 145940 694600 146180 694840
rect 146290 694600 146530 694840
rect 146620 694600 146860 694840
rect 146950 694600 147190 694840
rect 147280 694600 147520 694840
rect 147630 694600 147870 694840
rect 147960 694600 148200 694840
rect 148290 694600 148530 694840
rect 148620 694600 148860 694840
rect 148970 694600 149210 694840
rect 149300 694600 149540 694840
rect 149630 694600 149870 694840
rect 149960 694600 150200 694840
rect 150310 694600 150550 694840
rect 150640 694600 150880 694840
rect 150970 694600 151210 694840
rect 151300 694600 151540 694840
rect 151650 694600 151890 694840
rect 151980 694600 152220 694840
rect 152310 694600 152550 694840
rect 152640 694600 152880 694840
rect 152990 694600 153230 694840
rect 153320 694600 153560 694840
rect 153650 694600 153890 694840
rect 153980 694600 154220 694840
rect 154330 694600 154570 694840
rect 154660 694600 154900 694840
rect 154990 694600 155230 694840
rect 155320 694600 155560 694840
rect 155670 694600 155910 694840
rect 144950 694250 145190 694490
rect 145280 694250 145520 694490
rect 145610 694250 145850 694490
rect 145940 694250 146180 694490
rect 146290 694250 146530 694490
rect 146620 694250 146860 694490
rect 146950 694250 147190 694490
rect 147280 694250 147520 694490
rect 147630 694250 147870 694490
rect 147960 694250 148200 694490
rect 148290 694250 148530 694490
rect 148620 694250 148860 694490
rect 148970 694250 149210 694490
rect 149300 694250 149540 694490
rect 149630 694250 149870 694490
rect 149960 694250 150200 694490
rect 150310 694250 150550 694490
rect 150640 694250 150880 694490
rect 150970 694250 151210 694490
rect 151300 694250 151540 694490
rect 151650 694250 151890 694490
rect 151980 694250 152220 694490
rect 152310 694250 152550 694490
rect 152640 694250 152880 694490
rect 152990 694250 153230 694490
rect 153320 694250 153560 694490
rect 153650 694250 153890 694490
rect 153980 694250 154220 694490
rect 154330 694250 154570 694490
rect 154660 694250 154900 694490
rect 154990 694250 155230 694490
rect 155320 694250 155560 694490
rect 155670 694250 155910 694490
rect 144950 693920 145190 694160
rect 145280 693920 145520 694160
rect 145610 693920 145850 694160
rect 145940 693920 146180 694160
rect 146290 693920 146530 694160
rect 146620 693920 146860 694160
rect 146950 693920 147190 694160
rect 147280 693920 147520 694160
rect 147630 693920 147870 694160
rect 147960 693920 148200 694160
rect 148290 693920 148530 694160
rect 148620 693920 148860 694160
rect 148970 693920 149210 694160
rect 149300 693920 149540 694160
rect 149630 693920 149870 694160
rect 149960 693920 150200 694160
rect 150310 693920 150550 694160
rect 150640 693920 150880 694160
rect 150970 693920 151210 694160
rect 151300 693920 151540 694160
rect 151650 693920 151890 694160
rect 151980 693920 152220 694160
rect 152310 693920 152550 694160
rect 152640 693920 152880 694160
rect 152990 693920 153230 694160
rect 153320 693920 153560 694160
rect 153650 693920 153890 694160
rect 153980 693920 154220 694160
rect 154330 693920 154570 694160
rect 154660 693920 154900 694160
rect 154990 693920 155230 694160
rect 155320 693920 155560 694160
rect 155670 693920 155910 694160
rect 144950 693590 145190 693830
rect 145280 693590 145520 693830
rect 145610 693590 145850 693830
rect 145940 693590 146180 693830
rect 146290 693590 146530 693830
rect 146620 693590 146860 693830
rect 146950 693590 147190 693830
rect 147280 693590 147520 693830
rect 147630 693590 147870 693830
rect 147960 693590 148200 693830
rect 148290 693590 148530 693830
rect 148620 693590 148860 693830
rect 148970 693590 149210 693830
rect 149300 693590 149540 693830
rect 149630 693590 149870 693830
rect 149960 693590 150200 693830
rect 150310 693590 150550 693830
rect 150640 693590 150880 693830
rect 150970 693590 151210 693830
rect 151300 693590 151540 693830
rect 151650 693590 151890 693830
rect 151980 693590 152220 693830
rect 152310 693590 152550 693830
rect 152640 693590 152880 693830
rect 152990 693590 153230 693830
rect 153320 693590 153560 693830
rect 153650 693590 153890 693830
rect 153980 693590 154220 693830
rect 154330 693590 154570 693830
rect 154660 693590 154900 693830
rect 154990 693590 155230 693830
rect 155320 693590 155560 693830
rect 155670 693590 155910 693830
rect 144950 693260 145190 693500
rect 145280 693260 145520 693500
rect 145610 693260 145850 693500
rect 145940 693260 146180 693500
rect 146290 693260 146530 693500
rect 146620 693260 146860 693500
rect 146950 693260 147190 693500
rect 147280 693260 147520 693500
rect 147630 693260 147870 693500
rect 147960 693260 148200 693500
rect 148290 693260 148530 693500
rect 148620 693260 148860 693500
rect 148970 693260 149210 693500
rect 149300 693260 149540 693500
rect 149630 693260 149870 693500
rect 149960 693260 150200 693500
rect 150310 693260 150550 693500
rect 150640 693260 150880 693500
rect 150970 693260 151210 693500
rect 151300 693260 151540 693500
rect 151650 693260 151890 693500
rect 151980 693260 152220 693500
rect 152310 693260 152550 693500
rect 152640 693260 152880 693500
rect 152990 693260 153230 693500
rect 153320 693260 153560 693500
rect 153650 693260 153890 693500
rect 153980 693260 154220 693500
rect 154330 693260 154570 693500
rect 154660 693260 154900 693500
rect 154990 693260 155230 693500
rect 155320 693260 155560 693500
rect 155670 693260 155910 693500
rect 144950 692910 145190 693150
rect 145280 692910 145520 693150
rect 145610 692910 145850 693150
rect 145940 692910 146180 693150
rect 146290 692910 146530 693150
rect 146620 692910 146860 693150
rect 146950 692910 147190 693150
rect 147280 692910 147520 693150
rect 147630 692910 147870 693150
rect 147960 692910 148200 693150
rect 148290 692910 148530 693150
rect 148620 692910 148860 693150
rect 148970 692910 149210 693150
rect 149300 692910 149540 693150
rect 149630 692910 149870 693150
rect 149960 692910 150200 693150
rect 150310 692910 150550 693150
rect 150640 692910 150880 693150
rect 150970 692910 151210 693150
rect 151300 692910 151540 693150
rect 151650 692910 151890 693150
rect 151980 692910 152220 693150
rect 152310 692910 152550 693150
rect 152640 692910 152880 693150
rect 152990 692910 153230 693150
rect 153320 692910 153560 693150
rect 153650 692910 153890 693150
rect 153980 692910 154220 693150
rect 154330 692910 154570 693150
rect 154660 692910 154900 693150
rect 154990 692910 155230 693150
rect 155320 692910 155560 693150
rect 155670 692910 155910 693150
rect 144950 692580 145190 692820
rect 145280 692580 145520 692820
rect 145610 692580 145850 692820
rect 145940 692580 146180 692820
rect 146290 692580 146530 692820
rect 146620 692580 146860 692820
rect 146950 692580 147190 692820
rect 147280 692580 147520 692820
rect 147630 692580 147870 692820
rect 147960 692580 148200 692820
rect 148290 692580 148530 692820
rect 148620 692580 148860 692820
rect 148970 692580 149210 692820
rect 149300 692580 149540 692820
rect 149630 692580 149870 692820
rect 149960 692580 150200 692820
rect 150310 692580 150550 692820
rect 150640 692580 150880 692820
rect 150970 692580 151210 692820
rect 151300 692580 151540 692820
rect 151650 692580 151890 692820
rect 151980 692580 152220 692820
rect 152310 692580 152550 692820
rect 152640 692580 152880 692820
rect 152990 692580 153230 692820
rect 153320 692580 153560 692820
rect 153650 692580 153890 692820
rect 153980 692580 154220 692820
rect 154330 692580 154570 692820
rect 154660 692580 154900 692820
rect 154990 692580 155230 692820
rect 155320 692580 155560 692820
rect 155670 692580 155910 692820
rect 144950 692250 145190 692490
rect 145280 692250 145520 692490
rect 145610 692250 145850 692490
rect 145940 692250 146180 692490
rect 146290 692250 146530 692490
rect 146620 692250 146860 692490
rect 146950 692250 147190 692490
rect 147280 692250 147520 692490
rect 147630 692250 147870 692490
rect 147960 692250 148200 692490
rect 148290 692250 148530 692490
rect 148620 692250 148860 692490
rect 148970 692250 149210 692490
rect 149300 692250 149540 692490
rect 149630 692250 149870 692490
rect 149960 692250 150200 692490
rect 150310 692250 150550 692490
rect 150640 692250 150880 692490
rect 150970 692250 151210 692490
rect 151300 692250 151540 692490
rect 151650 692250 151890 692490
rect 151980 692250 152220 692490
rect 152310 692250 152550 692490
rect 152640 692250 152880 692490
rect 152990 692250 153230 692490
rect 153320 692250 153560 692490
rect 153650 692250 153890 692490
rect 153980 692250 154220 692490
rect 154330 692250 154570 692490
rect 154660 692250 154900 692490
rect 154990 692250 155230 692490
rect 155320 692250 155560 692490
rect 155670 692250 155910 692490
rect 144950 691920 145190 692160
rect 145280 691920 145520 692160
rect 145610 691920 145850 692160
rect 145940 691920 146180 692160
rect 146290 691920 146530 692160
rect 146620 691920 146860 692160
rect 146950 691920 147190 692160
rect 147280 691920 147520 692160
rect 147630 691920 147870 692160
rect 147960 691920 148200 692160
rect 148290 691920 148530 692160
rect 148620 691920 148860 692160
rect 148970 691920 149210 692160
rect 149300 691920 149540 692160
rect 149630 691920 149870 692160
rect 149960 691920 150200 692160
rect 150310 691920 150550 692160
rect 150640 691920 150880 692160
rect 150970 691920 151210 692160
rect 151300 691920 151540 692160
rect 151650 691920 151890 692160
rect 151980 691920 152220 692160
rect 152310 691920 152550 692160
rect 152640 691920 152880 692160
rect 152990 691920 153230 692160
rect 153320 691920 153560 692160
rect 153650 691920 153890 692160
rect 153980 691920 154220 692160
rect 154330 691920 154570 692160
rect 154660 691920 154900 692160
rect 154990 691920 155230 692160
rect 155320 691920 155560 692160
rect 155670 691920 155910 692160
rect 144950 691570 145190 691810
rect 145280 691570 145520 691810
rect 145610 691570 145850 691810
rect 145940 691570 146180 691810
rect 146290 691570 146530 691810
rect 146620 691570 146860 691810
rect 146950 691570 147190 691810
rect 147280 691570 147520 691810
rect 147630 691570 147870 691810
rect 147960 691570 148200 691810
rect 148290 691570 148530 691810
rect 148620 691570 148860 691810
rect 148970 691570 149210 691810
rect 149300 691570 149540 691810
rect 149630 691570 149870 691810
rect 149960 691570 150200 691810
rect 150310 691570 150550 691810
rect 150640 691570 150880 691810
rect 150970 691570 151210 691810
rect 151300 691570 151540 691810
rect 151650 691570 151890 691810
rect 151980 691570 152220 691810
rect 152310 691570 152550 691810
rect 152640 691570 152880 691810
rect 152990 691570 153230 691810
rect 153320 691570 153560 691810
rect 153650 691570 153890 691810
rect 153980 691570 154220 691810
rect 154330 691570 154570 691810
rect 154660 691570 154900 691810
rect 154990 691570 155230 691810
rect 155320 691570 155560 691810
rect 155670 691570 155910 691810
rect 144950 691240 145190 691480
rect 145280 691240 145520 691480
rect 145610 691240 145850 691480
rect 145940 691240 146180 691480
rect 146290 691240 146530 691480
rect 146620 691240 146860 691480
rect 146950 691240 147190 691480
rect 147280 691240 147520 691480
rect 147630 691240 147870 691480
rect 147960 691240 148200 691480
rect 148290 691240 148530 691480
rect 148620 691240 148860 691480
rect 148970 691240 149210 691480
rect 149300 691240 149540 691480
rect 149630 691240 149870 691480
rect 149960 691240 150200 691480
rect 150310 691240 150550 691480
rect 150640 691240 150880 691480
rect 150970 691240 151210 691480
rect 151300 691240 151540 691480
rect 151650 691240 151890 691480
rect 151980 691240 152220 691480
rect 152310 691240 152550 691480
rect 152640 691240 152880 691480
rect 152990 691240 153230 691480
rect 153320 691240 153560 691480
rect 153650 691240 153890 691480
rect 153980 691240 154220 691480
rect 154330 691240 154570 691480
rect 154660 691240 154900 691480
rect 154990 691240 155230 691480
rect 155320 691240 155560 691480
rect 155670 691240 155910 691480
rect 144950 690910 145190 691150
rect 145280 690910 145520 691150
rect 145610 690910 145850 691150
rect 145940 690910 146180 691150
rect 146290 690910 146530 691150
rect 146620 690910 146860 691150
rect 146950 690910 147190 691150
rect 147280 690910 147520 691150
rect 147630 690910 147870 691150
rect 147960 690910 148200 691150
rect 148290 690910 148530 691150
rect 148620 690910 148860 691150
rect 148970 690910 149210 691150
rect 149300 690910 149540 691150
rect 149630 690910 149870 691150
rect 149960 690910 150200 691150
rect 150310 690910 150550 691150
rect 150640 690910 150880 691150
rect 150970 690910 151210 691150
rect 151300 690910 151540 691150
rect 151650 690910 151890 691150
rect 151980 690910 152220 691150
rect 152310 690910 152550 691150
rect 152640 690910 152880 691150
rect 152990 690910 153230 691150
rect 153320 690910 153560 691150
rect 153650 690910 153890 691150
rect 153980 690910 154220 691150
rect 154330 690910 154570 691150
rect 154660 690910 154900 691150
rect 154990 690910 155230 691150
rect 155320 690910 155560 691150
rect 155670 690910 155910 691150
rect 144950 690580 145190 690820
rect 145280 690580 145520 690820
rect 145610 690580 145850 690820
rect 145940 690580 146180 690820
rect 146290 690580 146530 690820
rect 146620 690580 146860 690820
rect 146950 690580 147190 690820
rect 147280 690580 147520 690820
rect 147630 690580 147870 690820
rect 147960 690580 148200 690820
rect 148290 690580 148530 690820
rect 148620 690580 148860 690820
rect 148970 690580 149210 690820
rect 149300 690580 149540 690820
rect 149630 690580 149870 690820
rect 149960 690580 150200 690820
rect 150310 690580 150550 690820
rect 150640 690580 150880 690820
rect 150970 690580 151210 690820
rect 151300 690580 151540 690820
rect 151650 690580 151890 690820
rect 151980 690580 152220 690820
rect 152310 690580 152550 690820
rect 152640 690580 152880 690820
rect 152990 690580 153230 690820
rect 153320 690580 153560 690820
rect 153650 690580 153890 690820
rect 153980 690580 154220 690820
rect 154330 690580 154570 690820
rect 154660 690580 154900 690820
rect 154990 690580 155230 690820
rect 155320 690580 155560 690820
rect 155670 690580 155910 690820
rect 144950 690230 145190 690470
rect 145280 690230 145520 690470
rect 145610 690230 145850 690470
rect 145940 690230 146180 690470
rect 146290 690230 146530 690470
rect 146620 690230 146860 690470
rect 146950 690230 147190 690470
rect 147280 690230 147520 690470
rect 147630 690230 147870 690470
rect 147960 690230 148200 690470
rect 148290 690230 148530 690470
rect 148620 690230 148860 690470
rect 148970 690230 149210 690470
rect 149300 690230 149540 690470
rect 149630 690230 149870 690470
rect 149960 690230 150200 690470
rect 150310 690230 150550 690470
rect 150640 690230 150880 690470
rect 150970 690230 151210 690470
rect 151300 690230 151540 690470
rect 151650 690230 151890 690470
rect 151980 690230 152220 690470
rect 152310 690230 152550 690470
rect 152640 690230 152880 690470
rect 152990 690230 153230 690470
rect 153320 690230 153560 690470
rect 153650 690230 153890 690470
rect 153980 690230 154220 690470
rect 154330 690230 154570 690470
rect 154660 690230 154900 690470
rect 154990 690230 155230 690470
rect 155320 690230 155560 690470
rect 155670 690230 155910 690470
rect 144950 689900 145190 690140
rect 145280 689900 145520 690140
rect 145610 689900 145850 690140
rect 145940 689900 146180 690140
rect 146290 689900 146530 690140
rect 146620 689900 146860 690140
rect 146950 689900 147190 690140
rect 147280 689900 147520 690140
rect 147630 689900 147870 690140
rect 147960 689900 148200 690140
rect 148290 689900 148530 690140
rect 148620 689900 148860 690140
rect 148970 689900 149210 690140
rect 149300 689900 149540 690140
rect 149630 689900 149870 690140
rect 149960 689900 150200 690140
rect 150310 689900 150550 690140
rect 150640 689900 150880 690140
rect 150970 689900 151210 690140
rect 151300 689900 151540 690140
rect 151650 689900 151890 690140
rect 151980 689900 152220 690140
rect 152310 689900 152550 690140
rect 152640 689900 152880 690140
rect 152990 689900 153230 690140
rect 153320 689900 153560 690140
rect 153650 689900 153890 690140
rect 153980 689900 154220 690140
rect 154330 689900 154570 690140
rect 154660 689900 154900 690140
rect 154990 689900 155230 690140
rect 155320 689900 155560 690140
rect 155670 689900 155910 690140
rect 144950 689570 145190 689810
rect 145280 689570 145520 689810
rect 145610 689570 145850 689810
rect 145940 689570 146180 689810
rect 146290 689570 146530 689810
rect 146620 689570 146860 689810
rect 146950 689570 147190 689810
rect 147280 689570 147520 689810
rect 147630 689570 147870 689810
rect 147960 689570 148200 689810
rect 148290 689570 148530 689810
rect 148620 689570 148860 689810
rect 148970 689570 149210 689810
rect 149300 689570 149540 689810
rect 149630 689570 149870 689810
rect 149960 689570 150200 689810
rect 150310 689570 150550 689810
rect 150640 689570 150880 689810
rect 150970 689570 151210 689810
rect 151300 689570 151540 689810
rect 151650 689570 151890 689810
rect 151980 689570 152220 689810
rect 152310 689570 152550 689810
rect 152640 689570 152880 689810
rect 152990 689570 153230 689810
rect 153320 689570 153560 689810
rect 153650 689570 153890 689810
rect 153980 689570 154220 689810
rect 154330 689570 154570 689810
rect 154660 689570 154900 689810
rect 154990 689570 155230 689810
rect 155320 689570 155560 689810
rect 155670 689570 155910 689810
rect 144950 689240 145190 689480
rect 145280 689240 145520 689480
rect 145610 689240 145850 689480
rect 145940 689240 146180 689480
rect 146290 689240 146530 689480
rect 146620 689240 146860 689480
rect 146950 689240 147190 689480
rect 147280 689240 147520 689480
rect 147630 689240 147870 689480
rect 147960 689240 148200 689480
rect 148290 689240 148530 689480
rect 148620 689240 148860 689480
rect 148970 689240 149210 689480
rect 149300 689240 149540 689480
rect 149630 689240 149870 689480
rect 149960 689240 150200 689480
rect 150310 689240 150550 689480
rect 150640 689240 150880 689480
rect 150970 689240 151210 689480
rect 151300 689240 151540 689480
rect 151650 689240 151890 689480
rect 151980 689240 152220 689480
rect 152310 689240 152550 689480
rect 152640 689240 152880 689480
rect 152990 689240 153230 689480
rect 153320 689240 153560 689480
rect 153650 689240 153890 689480
rect 153980 689240 154220 689480
rect 154330 689240 154570 689480
rect 154660 689240 154900 689480
rect 154990 689240 155230 689480
rect 155320 689240 155560 689480
rect 155670 689240 155910 689480
rect 144950 688890 145190 689130
rect 145280 688890 145520 689130
rect 145610 688890 145850 689130
rect 145940 688890 146180 689130
rect 146290 688890 146530 689130
rect 146620 688890 146860 689130
rect 146950 688890 147190 689130
rect 147280 688890 147520 689130
rect 147630 688890 147870 689130
rect 147960 688890 148200 689130
rect 148290 688890 148530 689130
rect 148620 688890 148860 689130
rect 148970 688890 149210 689130
rect 149300 688890 149540 689130
rect 149630 688890 149870 689130
rect 149960 688890 150200 689130
rect 150310 688890 150550 689130
rect 150640 688890 150880 689130
rect 150970 688890 151210 689130
rect 151300 688890 151540 689130
rect 151650 688890 151890 689130
rect 151980 688890 152220 689130
rect 152310 688890 152550 689130
rect 152640 688890 152880 689130
rect 152990 688890 153230 689130
rect 153320 688890 153560 689130
rect 153650 688890 153890 689130
rect 153980 688890 154220 689130
rect 154330 688890 154570 689130
rect 154660 688890 154900 689130
rect 154990 688890 155230 689130
rect 155320 688890 155560 689130
rect 155670 688890 155910 689130
rect 144950 688560 145190 688800
rect 145280 688560 145520 688800
rect 145610 688560 145850 688800
rect 145940 688560 146180 688800
rect 146290 688560 146530 688800
rect 146620 688560 146860 688800
rect 146950 688560 147190 688800
rect 147280 688560 147520 688800
rect 147630 688560 147870 688800
rect 147960 688560 148200 688800
rect 148290 688560 148530 688800
rect 148620 688560 148860 688800
rect 148970 688560 149210 688800
rect 149300 688560 149540 688800
rect 149630 688560 149870 688800
rect 149960 688560 150200 688800
rect 150310 688560 150550 688800
rect 150640 688560 150880 688800
rect 150970 688560 151210 688800
rect 151300 688560 151540 688800
rect 151650 688560 151890 688800
rect 151980 688560 152220 688800
rect 152310 688560 152550 688800
rect 152640 688560 152880 688800
rect 152990 688560 153230 688800
rect 153320 688560 153560 688800
rect 153650 688560 153890 688800
rect 153980 688560 154220 688800
rect 154330 688560 154570 688800
rect 154660 688560 154900 688800
rect 154990 688560 155230 688800
rect 155320 688560 155560 688800
rect 155670 688560 155910 688800
rect 144950 688230 145190 688470
rect 145280 688230 145520 688470
rect 145610 688230 145850 688470
rect 145940 688230 146180 688470
rect 146290 688230 146530 688470
rect 146620 688230 146860 688470
rect 146950 688230 147190 688470
rect 147280 688230 147520 688470
rect 147630 688230 147870 688470
rect 147960 688230 148200 688470
rect 148290 688230 148530 688470
rect 148620 688230 148860 688470
rect 148970 688230 149210 688470
rect 149300 688230 149540 688470
rect 149630 688230 149870 688470
rect 149960 688230 150200 688470
rect 150310 688230 150550 688470
rect 150640 688230 150880 688470
rect 150970 688230 151210 688470
rect 151300 688230 151540 688470
rect 151650 688230 151890 688470
rect 151980 688230 152220 688470
rect 152310 688230 152550 688470
rect 152640 688230 152880 688470
rect 152990 688230 153230 688470
rect 153320 688230 153560 688470
rect 153650 688230 153890 688470
rect 153980 688230 154220 688470
rect 154330 688230 154570 688470
rect 154660 688230 154900 688470
rect 154990 688230 155230 688470
rect 155320 688230 155560 688470
rect 155670 688230 155910 688470
rect 144950 687900 145190 688140
rect 145280 687900 145520 688140
rect 145610 687900 145850 688140
rect 145940 687900 146180 688140
rect 146290 687900 146530 688140
rect 146620 687900 146860 688140
rect 146950 687900 147190 688140
rect 147280 687900 147520 688140
rect 147630 687900 147870 688140
rect 147960 687900 148200 688140
rect 148290 687900 148530 688140
rect 148620 687900 148860 688140
rect 148970 687900 149210 688140
rect 149300 687900 149540 688140
rect 149630 687900 149870 688140
rect 149960 687900 150200 688140
rect 150310 687900 150550 688140
rect 150640 687900 150880 688140
rect 150970 687900 151210 688140
rect 151300 687900 151540 688140
rect 151650 687900 151890 688140
rect 151980 687900 152220 688140
rect 152310 687900 152550 688140
rect 152640 687900 152880 688140
rect 152990 687900 153230 688140
rect 153320 687900 153560 688140
rect 153650 687900 153890 688140
rect 153980 687900 154220 688140
rect 154330 687900 154570 688140
rect 154660 687900 154900 688140
rect 154990 687900 155230 688140
rect 155320 687900 155560 688140
rect 155670 687900 155910 688140
rect 144950 687550 145190 687790
rect 145280 687550 145520 687790
rect 145610 687550 145850 687790
rect 145940 687550 146180 687790
rect 146290 687550 146530 687790
rect 146620 687550 146860 687790
rect 146950 687550 147190 687790
rect 147280 687550 147520 687790
rect 147630 687550 147870 687790
rect 147960 687550 148200 687790
rect 148290 687550 148530 687790
rect 148620 687550 148860 687790
rect 148970 687550 149210 687790
rect 149300 687550 149540 687790
rect 149630 687550 149870 687790
rect 149960 687550 150200 687790
rect 150310 687550 150550 687790
rect 150640 687550 150880 687790
rect 150970 687550 151210 687790
rect 151300 687550 151540 687790
rect 151650 687550 151890 687790
rect 151980 687550 152220 687790
rect 152310 687550 152550 687790
rect 152640 687550 152880 687790
rect 152990 687550 153230 687790
rect 153320 687550 153560 687790
rect 153650 687550 153890 687790
rect 153980 687550 154220 687790
rect 154330 687550 154570 687790
rect 154660 687550 154900 687790
rect 154990 687550 155230 687790
rect 155320 687550 155560 687790
rect 155670 687550 155910 687790
rect 144950 687220 145190 687460
rect 145280 687220 145520 687460
rect 145610 687220 145850 687460
rect 145940 687220 146180 687460
rect 146290 687220 146530 687460
rect 146620 687220 146860 687460
rect 146950 687220 147190 687460
rect 147280 687220 147520 687460
rect 147630 687220 147870 687460
rect 147960 687220 148200 687460
rect 148290 687220 148530 687460
rect 148620 687220 148860 687460
rect 148970 687220 149210 687460
rect 149300 687220 149540 687460
rect 149630 687220 149870 687460
rect 149960 687220 150200 687460
rect 150310 687220 150550 687460
rect 150640 687220 150880 687460
rect 150970 687220 151210 687460
rect 151300 687220 151540 687460
rect 151650 687220 151890 687460
rect 151980 687220 152220 687460
rect 152310 687220 152550 687460
rect 152640 687220 152880 687460
rect 152990 687220 153230 687460
rect 153320 687220 153560 687460
rect 153650 687220 153890 687460
rect 153980 687220 154220 687460
rect 154330 687220 154570 687460
rect 154660 687220 154900 687460
rect 154990 687220 155230 687460
rect 155320 687220 155560 687460
rect 155670 687220 155910 687460
rect 144950 686890 145190 687130
rect 145280 686890 145520 687130
rect 145610 686890 145850 687130
rect 145940 686890 146180 687130
rect 146290 686890 146530 687130
rect 146620 686890 146860 687130
rect 146950 686890 147190 687130
rect 147280 686890 147520 687130
rect 147630 686890 147870 687130
rect 147960 686890 148200 687130
rect 148290 686890 148530 687130
rect 148620 686890 148860 687130
rect 148970 686890 149210 687130
rect 149300 686890 149540 687130
rect 149630 686890 149870 687130
rect 149960 686890 150200 687130
rect 150310 686890 150550 687130
rect 150640 686890 150880 687130
rect 150970 686890 151210 687130
rect 151300 686890 151540 687130
rect 151650 686890 151890 687130
rect 151980 686890 152220 687130
rect 152310 686890 152550 687130
rect 152640 686890 152880 687130
rect 152990 686890 153230 687130
rect 153320 686890 153560 687130
rect 153650 686890 153890 687130
rect 153980 686890 154220 687130
rect 154330 686890 154570 687130
rect 154660 686890 154900 687130
rect 154990 686890 155230 687130
rect 155320 686890 155560 687130
rect 155670 686890 155910 687130
rect 144950 686560 145190 686800
rect 145280 686560 145520 686800
rect 145610 686560 145850 686800
rect 145940 686560 146180 686800
rect 146290 686560 146530 686800
rect 146620 686560 146860 686800
rect 146950 686560 147190 686800
rect 147280 686560 147520 686800
rect 147630 686560 147870 686800
rect 147960 686560 148200 686800
rect 148290 686560 148530 686800
rect 148620 686560 148860 686800
rect 148970 686560 149210 686800
rect 149300 686560 149540 686800
rect 149630 686560 149870 686800
rect 149960 686560 150200 686800
rect 150310 686560 150550 686800
rect 150640 686560 150880 686800
rect 150970 686560 151210 686800
rect 151300 686560 151540 686800
rect 151650 686560 151890 686800
rect 151980 686560 152220 686800
rect 152310 686560 152550 686800
rect 152640 686560 152880 686800
rect 152990 686560 153230 686800
rect 153320 686560 153560 686800
rect 153650 686560 153890 686800
rect 153980 686560 154220 686800
rect 154330 686560 154570 686800
rect 154660 686560 154900 686800
rect 154990 686560 155230 686800
rect 155320 686560 155560 686800
rect 155670 686560 155910 686800
rect 144950 686210 145190 686450
rect 145280 686210 145520 686450
rect 145610 686210 145850 686450
rect 145940 686210 146180 686450
rect 146290 686210 146530 686450
rect 146620 686210 146860 686450
rect 146950 686210 147190 686450
rect 147280 686210 147520 686450
rect 147630 686210 147870 686450
rect 147960 686210 148200 686450
rect 148290 686210 148530 686450
rect 148620 686210 148860 686450
rect 148970 686210 149210 686450
rect 149300 686210 149540 686450
rect 149630 686210 149870 686450
rect 149960 686210 150200 686450
rect 150310 686210 150550 686450
rect 150640 686210 150880 686450
rect 150970 686210 151210 686450
rect 151300 686210 151540 686450
rect 151650 686210 151890 686450
rect 151980 686210 152220 686450
rect 152310 686210 152550 686450
rect 152640 686210 152880 686450
rect 152990 686210 153230 686450
rect 153320 686210 153560 686450
rect 153650 686210 153890 686450
rect 153980 686210 154220 686450
rect 154330 686210 154570 686450
rect 154660 686210 154900 686450
rect 154990 686210 155230 686450
rect 155320 686210 155560 686450
rect 155670 686210 155910 686450
rect 144950 685880 145190 686120
rect 145280 685880 145520 686120
rect 145610 685880 145850 686120
rect 145940 685880 146180 686120
rect 146290 685880 146530 686120
rect 146620 685880 146860 686120
rect 146950 685880 147190 686120
rect 147280 685880 147520 686120
rect 147630 685880 147870 686120
rect 147960 685880 148200 686120
rect 148290 685880 148530 686120
rect 148620 685880 148860 686120
rect 148970 685880 149210 686120
rect 149300 685880 149540 686120
rect 149630 685880 149870 686120
rect 149960 685880 150200 686120
rect 150310 685880 150550 686120
rect 150640 685880 150880 686120
rect 150970 685880 151210 686120
rect 151300 685880 151540 686120
rect 151650 685880 151890 686120
rect 151980 685880 152220 686120
rect 152310 685880 152550 686120
rect 152640 685880 152880 686120
rect 152990 685880 153230 686120
rect 153320 685880 153560 686120
rect 153650 685880 153890 686120
rect 153980 685880 154220 686120
rect 154330 685880 154570 686120
rect 154660 685880 154900 686120
rect 154990 685880 155230 686120
rect 155320 685880 155560 686120
rect 155670 685880 155910 686120
rect 144950 685550 145190 685790
rect 145280 685550 145520 685790
rect 145610 685550 145850 685790
rect 145940 685550 146180 685790
rect 146290 685550 146530 685790
rect 146620 685550 146860 685790
rect 146950 685550 147190 685790
rect 147280 685550 147520 685790
rect 147630 685550 147870 685790
rect 147960 685550 148200 685790
rect 148290 685550 148530 685790
rect 148620 685550 148860 685790
rect 148970 685550 149210 685790
rect 149300 685550 149540 685790
rect 149630 685550 149870 685790
rect 149960 685550 150200 685790
rect 150310 685550 150550 685790
rect 150640 685550 150880 685790
rect 150970 685550 151210 685790
rect 151300 685550 151540 685790
rect 151650 685550 151890 685790
rect 151980 685550 152220 685790
rect 152310 685550 152550 685790
rect 152640 685550 152880 685790
rect 152990 685550 153230 685790
rect 153320 685550 153560 685790
rect 153650 685550 153890 685790
rect 153980 685550 154220 685790
rect 154330 685550 154570 685790
rect 154660 685550 154900 685790
rect 154990 685550 155230 685790
rect 155320 685550 155560 685790
rect 155670 685550 155910 685790
rect 144950 685220 145190 685460
rect 145280 685220 145520 685460
rect 145610 685220 145850 685460
rect 145940 685220 146180 685460
rect 146290 685220 146530 685460
rect 146620 685220 146860 685460
rect 146950 685220 147190 685460
rect 147280 685220 147520 685460
rect 147630 685220 147870 685460
rect 147960 685220 148200 685460
rect 148290 685220 148530 685460
rect 148620 685220 148860 685460
rect 148970 685220 149210 685460
rect 149300 685220 149540 685460
rect 149630 685220 149870 685460
rect 149960 685220 150200 685460
rect 150310 685220 150550 685460
rect 150640 685220 150880 685460
rect 150970 685220 151210 685460
rect 151300 685220 151540 685460
rect 151650 685220 151890 685460
rect 151980 685220 152220 685460
rect 152310 685220 152550 685460
rect 152640 685220 152880 685460
rect 152990 685220 153230 685460
rect 153320 685220 153560 685460
rect 153650 685220 153890 685460
rect 153980 685220 154220 685460
rect 154330 685220 154570 685460
rect 154660 685220 154900 685460
rect 154990 685220 155230 685460
rect 155320 685220 155560 685460
rect 155670 685220 155910 685460
rect 144950 684870 145190 685110
rect 145280 684870 145520 685110
rect 145610 684870 145850 685110
rect 145940 684870 146180 685110
rect 146290 684870 146530 685110
rect 146620 684870 146860 685110
rect 146950 684870 147190 685110
rect 147280 684870 147520 685110
rect 147630 684870 147870 685110
rect 147960 684870 148200 685110
rect 148290 684870 148530 685110
rect 148620 684870 148860 685110
rect 148970 684870 149210 685110
rect 149300 684870 149540 685110
rect 149630 684870 149870 685110
rect 149960 684870 150200 685110
rect 150310 684870 150550 685110
rect 150640 684870 150880 685110
rect 150970 684870 151210 685110
rect 151300 684870 151540 685110
rect 151650 684870 151890 685110
rect 151980 684870 152220 685110
rect 152310 684870 152550 685110
rect 152640 684870 152880 685110
rect 152990 684870 153230 685110
rect 153320 684870 153560 685110
rect 153650 684870 153890 685110
rect 153980 684870 154220 685110
rect 154330 684870 154570 685110
rect 154660 684870 154900 685110
rect 154990 684870 155230 685110
rect 155320 684870 155560 685110
rect 155670 684870 155910 685110
rect 144950 684540 145190 684780
rect 145280 684540 145520 684780
rect 145610 684540 145850 684780
rect 145940 684540 146180 684780
rect 146290 684540 146530 684780
rect 146620 684540 146860 684780
rect 146950 684540 147190 684780
rect 147280 684540 147520 684780
rect 147630 684540 147870 684780
rect 147960 684540 148200 684780
rect 148290 684540 148530 684780
rect 148620 684540 148860 684780
rect 148970 684540 149210 684780
rect 149300 684540 149540 684780
rect 149630 684540 149870 684780
rect 149960 684540 150200 684780
rect 150310 684540 150550 684780
rect 150640 684540 150880 684780
rect 150970 684540 151210 684780
rect 151300 684540 151540 684780
rect 151650 684540 151890 684780
rect 151980 684540 152220 684780
rect 152310 684540 152550 684780
rect 152640 684540 152880 684780
rect 152990 684540 153230 684780
rect 153320 684540 153560 684780
rect 153650 684540 153890 684780
rect 153980 684540 154220 684780
rect 154330 684540 154570 684780
rect 154660 684540 154900 684780
rect 154990 684540 155230 684780
rect 155320 684540 155560 684780
rect 155670 684540 155910 684780
rect 144950 684210 145190 684450
rect 145280 684210 145520 684450
rect 145610 684210 145850 684450
rect 145940 684210 146180 684450
rect 146290 684210 146530 684450
rect 146620 684210 146860 684450
rect 146950 684210 147190 684450
rect 147280 684210 147520 684450
rect 147630 684210 147870 684450
rect 147960 684210 148200 684450
rect 148290 684210 148530 684450
rect 148620 684210 148860 684450
rect 148970 684210 149210 684450
rect 149300 684210 149540 684450
rect 149630 684210 149870 684450
rect 149960 684210 150200 684450
rect 150310 684210 150550 684450
rect 150640 684210 150880 684450
rect 150970 684210 151210 684450
rect 151300 684210 151540 684450
rect 151650 684210 151890 684450
rect 151980 684210 152220 684450
rect 152310 684210 152550 684450
rect 152640 684210 152880 684450
rect 152990 684210 153230 684450
rect 153320 684210 153560 684450
rect 153650 684210 153890 684450
rect 153980 684210 154220 684450
rect 154330 684210 154570 684450
rect 154660 684210 154900 684450
rect 154990 684210 155230 684450
rect 155320 684210 155560 684450
rect 155670 684210 155910 684450
rect 144950 683880 145190 684120
rect 145280 683880 145520 684120
rect 145610 683880 145850 684120
rect 145940 683880 146180 684120
rect 146290 683880 146530 684120
rect 146620 683880 146860 684120
rect 146950 683880 147190 684120
rect 147280 683880 147520 684120
rect 147630 683880 147870 684120
rect 147960 683880 148200 684120
rect 148290 683880 148530 684120
rect 148620 683880 148860 684120
rect 148970 683880 149210 684120
rect 149300 683880 149540 684120
rect 149630 683880 149870 684120
rect 149960 683880 150200 684120
rect 150310 683880 150550 684120
rect 150640 683880 150880 684120
rect 150970 683880 151210 684120
rect 151300 683880 151540 684120
rect 151650 683880 151890 684120
rect 151980 683880 152220 684120
rect 152310 683880 152550 684120
rect 152640 683880 152880 684120
rect 152990 683880 153230 684120
rect 153320 683880 153560 684120
rect 153650 683880 153890 684120
rect 153980 683880 154220 684120
rect 154330 683880 154570 684120
rect 154660 683880 154900 684120
rect 154990 683880 155230 684120
rect 155320 683880 155560 684120
rect 155670 683880 155910 684120
rect 110810 683040 111050 683280
rect 111160 683040 111400 683280
rect 111490 683040 111730 683280
rect 111820 683040 112060 683280
rect 112150 683040 112390 683280
rect 112500 683040 112740 683280
rect 112830 683040 113070 683280
rect 113160 683040 113400 683280
rect 113490 683040 113730 683280
rect 113840 683040 114080 683280
rect 114170 683040 114410 683280
rect 114500 683040 114740 683280
rect 114830 683040 115070 683280
rect 115180 683040 115420 683280
rect 115510 683040 115750 683280
rect 115840 683040 116080 683280
rect 116170 683040 116410 683280
rect 116520 683040 116760 683280
rect 116850 683040 117090 683280
rect 117180 683040 117420 683280
rect 117510 683040 117750 683280
rect 117860 683040 118100 683280
rect 118190 683040 118430 683280
rect 118520 683040 118760 683280
rect 118850 683040 119090 683280
rect 119200 683040 119440 683280
rect 119530 683040 119770 683280
rect 119860 683040 120100 683280
rect 120190 683040 120430 683280
rect 120540 683040 120780 683280
rect 120870 683040 121110 683280
rect 121200 683040 121440 683280
rect 121530 683040 121770 683280
rect 110810 682710 111050 682950
rect 111160 682710 111400 682950
rect 111490 682710 111730 682950
rect 111820 682710 112060 682950
rect 112150 682710 112390 682950
rect 112500 682710 112740 682950
rect 112830 682710 113070 682950
rect 113160 682710 113400 682950
rect 113490 682710 113730 682950
rect 113840 682710 114080 682950
rect 114170 682710 114410 682950
rect 114500 682710 114740 682950
rect 114830 682710 115070 682950
rect 115180 682710 115420 682950
rect 115510 682710 115750 682950
rect 115840 682710 116080 682950
rect 116170 682710 116410 682950
rect 116520 682710 116760 682950
rect 116850 682710 117090 682950
rect 117180 682710 117420 682950
rect 117510 682710 117750 682950
rect 117860 682710 118100 682950
rect 118190 682710 118430 682950
rect 118520 682710 118760 682950
rect 118850 682710 119090 682950
rect 119200 682710 119440 682950
rect 119530 682710 119770 682950
rect 119860 682710 120100 682950
rect 120190 682710 120430 682950
rect 120540 682710 120780 682950
rect 120870 682710 121110 682950
rect 121200 682710 121440 682950
rect 121530 682710 121770 682950
rect 110810 682380 111050 682620
rect 111160 682380 111400 682620
rect 111490 682380 111730 682620
rect 111820 682380 112060 682620
rect 112150 682380 112390 682620
rect 112500 682380 112740 682620
rect 112830 682380 113070 682620
rect 113160 682380 113400 682620
rect 113490 682380 113730 682620
rect 113840 682380 114080 682620
rect 114170 682380 114410 682620
rect 114500 682380 114740 682620
rect 114830 682380 115070 682620
rect 115180 682380 115420 682620
rect 115510 682380 115750 682620
rect 115840 682380 116080 682620
rect 116170 682380 116410 682620
rect 116520 682380 116760 682620
rect 116850 682380 117090 682620
rect 117180 682380 117420 682620
rect 117510 682380 117750 682620
rect 117860 682380 118100 682620
rect 118190 682380 118430 682620
rect 118520 682380 118760 682620
rect 118850 682380 119090 682620
rect 119200 682380 119440 682620
rect 119530 682380 119770 682620
rect 119860 682380 120100 682620
rect 120190 682380 120430 682620
rect 120540 682380 120780 682620
rect 120870 682380 121110 682620
rect 121200 682380 121440 682620
rect 121530 682380 121770 682620
rect 110810 682050 111050 682290
rect 111160 682050 111400 682290
rect 111490 682050 111730 682290
rect 111820 682050 112060 682290
rect 112150 682050 112390 682290
rect 112500 682050 112740 682290
rect 112830 682050 113070 682290
rect 113160 682050 113400 682290
rect 113490 682050 113730 682290
rect 113840 682050 114080 682290
rect 114170 682050 114410 682290
rect 114500 682050 114740 682290
rect 114830 682050 115070 682290
rect 115180 682050 115420 682290
rect 115510 682050 115750 682290
rect 115840 682050 116080 682290
rect 116170 682050 116410 682290
rect 116520 682050 116760 682290
rect 116850 682050 117090 682290
rect 117180 682050 117420 682290
rect 117510 682050 117750 682290
rect 117860 682050 118100 682290
rect 118190 682050 118430 682290
rect 118520 682050 118760 682290
rect 118850 682050 119090 682290
rect 119200 682050 119440 682290
rect 119530 682050 119770 682290
rect 119860 682050 120100 682290
rect 120190 682050 120430 682290
rect 120540 682050 120780 682290
rect 120870 682050 121110 682290
rect 121200 682050 121440 682290
rect 121530 682050 121770 682290
rect 110810 681700 111050 681940
rect 111160 681700 111400 681940
rect 111490 681700 111730 681940
rect 111820 681700 112060 681940
rect 112150 681700 112390 681940
rect 112500 681700 112740 681940
rect 112830 681700 113070 681940
rect 113160 681700 113400 681940
rect 113490 681700 113730 681940
rect 113840 681700 114080 681940
rect 114170 681700 114410 681940
rect 114500 681700 114740 681940
rect 114830 681700 115070 681940
rect 115180 681700 115420 681940
rect 115510 681700 115750 681940
rect 115840 681700 116080 681940
rect 116170 681700 116410 681940
rect 116520 681700 116760 681940
rect 116850 681700 117090 681940
rect 117180 681700 117420 681940
rect 117510 681700 117750 681940
rect 117860 681700 118100 681940
rect 118190 681700 118430 681940
rect 118520 681700 118760 681940
rect 118850 681700 119090 681940
rect 119200 681700 119440 681940
rect 119530 681700 119770 681940
rect 119860 681700 120100 681940
rect 120190 681700 120430 681940
rect 120540 681700 120780 681940
rect 120870 681700 121110 681940
rect 121200 681700 121440 681940
rect 121530 681700 121770 681940
rect 110810 681370 111050 681610
rect 111160 681370 111400 681610
rect 111490 681370 111730 681610
rect 111820 681370 112060 681610
rect 112150 681370 112390 681610
rect 112500 681370 112740 681610
rect 112830 681370 113070 681610
rect 113160 681370 113400 681610
rect 113490 681370 113730 681610
rect 113840 681370 114080 681610
rect 114170 681370 114410 681610
rect 114500 681370 114740 681610
rect 114830 681370 115070 681610
rect 115180 681370 115420 681610
rect 115510 681370 115750 681610
rect 115840 681370 116080 681610
rect 116170 681370 116410 681610
rect 116520 681370 116760 681610
rect 116850 681370 117090 681610
rect 117180 681370 117420 681610
rect 117510 681370 117750 681610
rect 117860 681370 118100 681610
rect 118190 681370 118430 681610
rect 118520 681370 118760 681610
rect 118850 681370 119090 681610
rect 119200 681370 119440 681610
rect 119530 681370 119770 681610
rect 119860 681370 120100 681610
rect 120190 681370 120430 681610
rect 120540 681370 120780 681610
rect 120870 681370 121110 681610
rect 121200 681370 121440 681610
rect 121530 681370 121770 681610
rect 110810 681040 111050 681280
rect 111160 681040 111400 681280
rect 111490 681040 111730 681280
rect 111820 681040 112060 681280
rect 112150 681040 112390 681280
rect 112500 681040 112740 681280
rect 112830 681040 113070 681280
rect 113160 681040 113400 681280
rect 113490 681040 113730 681280
rect 113840 681040 114080 681280
rect 114170 681040 114410 681280
rect 114500 681040 114740 681280
rect 114830 681040 115070 681280
rect 115180 681040 115420 681280
rect 115510 681040 115750 681280
rect 115840 681040 116080 681280
rect 116170 681040 116410 681280
rect 116520 681040 116760 681280
rect 116850 681040 117090 681280
rect 117180 681040 117420 681280
rect 117510 681040 117750 681280
rect 117860 681040 118100 681280
rect 118190 681040 118430 681280
rect 118520 681040 118760 681280
rect 118850 681040 119090 681280
rect 119200 681040 119440 681280
rect 119530 681040 119770 681280
rect 119860 681040 120100 681280
rect 120190 681040 120430 681280
rect 120540 681040 120780 681280
rect 120870 681040 121110 681280
rect 121200 681040 121440 681280
rect 121530 681040 121770 681280
rect 110810 680710 111050 680950
rect 111160 680710 111400 680950
rect 111490 680710 111730 680950
rect 111820 680710 112060 680950
rect 112150 680710 112390 680950
rect 112500 680710 112740 680950
rect 112830 680710 113070 680950
rect 113160 680710 113400 680950
rect 113490 680710 113730 680950
rect 113840 680710 114080 680950
rect 114170 680710 114410 680950
rect 114500 680710 114740 680950
rect 114830 680710 115070 680950
rect 115180 680710 115420 680950
rect 115510 680710 115750 680950
rect 115840 680710 116080 680950
rect 116170 680710 116410 680950
rect 116520 680710 116760 680950
rect 116850 680710 117090 680950
rect 117180 680710 117420 680950
rect 117510 680710 117750 680950
rect 117860 680710 118100 680950
rect 118190 680710 118430 680950
rect 118520 680710 118760 680950
rect 118850 680710 119090 680950
rect 119200 680710 119440 680950
rect 119530 680710 119770 680950
rect 119860 680710 120100 680950
rect 120190 680710 120430 680950
rect 120540 680710 120780 680950
rect 120870 680710 121110 680950
rect 121200 680710 121440 680950
rect 121530 680710 121770 680950
rect 110810 680360 111050 680600
rect 111160 680360 111400 680600
rect 111490 680360 111730 680600
rect 111820 680360 112060 680600
rect 112150 680360 112390 680600
rect 112500 680360 112740 680600
rect 112830 680360 113070 680600
rect 113160 680360 113400 680600
rect 113490 680360 113730 680600
rect 113840 680360 114080 680600
rect 114170 680360 114410 680600
rect 114500 680360 114740 680600
rect 114830 680360 115070 680600
rect 115180 680360 115420 680600
rect 115510 680360 115750 680600
rect 115840 680360 116080 680600
rect 116170 680360 116410 680600
rect 116520 680360 116760 680600
rect 116850 680360 117090 680600
rect 117180 680360 117420 680600
rect 117510 680360 117750 680600
rect 117860 680360 118100 680600
rect 118190 680360 118430 680600
rect 118520 680360 118760 680600
rect 118850 680360 119090 680600
rect 119200 680360 119440 680600
rect 119530 680360 119770 680600
rect 119860 680360 120100 680600
rect 120190 680360 120430 680600
rect 120540 680360 120780 680600
rect 120870 680360 121110 680600
rect 121200 680360 121440 680600
rect 121530 680360 121770 680600
rect 110810 680030 111050 680270
rect 111160 680030 111400 680270
rect 111490 680030 111730 680270
rect 111820 680030 112060 680270
rect 112150 680030 112390 680270
rect 112500 680030 112740 680270
rect 112830 680030 113070 680270
rect 113160 680030 113400 680270
rect 113490 680030 113730 680270
rect 113840 680030 114080 680270
rect 114170 680030 114410 680270
rect 114500 680030 114740 680270
rect 114830 680030 115070 680270
rect 115180 680030 115420 680270
rect 115510 680030 115750 680270
rect 115840 680030 116080 680270
rect 116170 680030 116410 680270
rect 116520 680030 116760 680270
rect 116850 680030 117090 680270
rect 117180 680030 117420 680270
rect 117510 680030 117750 680270
rect 117860 680030 118100 680270
rect 118190 680030 118430 680270
rect 118520 680030 118760 680270
rect 118850 680030 119090 680270
rect 119200 680030 119440 680270
rect 119530 680030 119770 680270
rect 119860 680030 120100 680270
rect 120190 680030 120430 680270
rect 120540 680030 120780 680270
rect 120870 680030 121110 680270
rect 121200 680030 121440 680270
rect 121530 680030 121770 680270
rect 110810 679700 111050 679940
rect 111160 679700 111400 679940
rect 111490 679700 111730 679940
rect 111820 679700 112060 679940
rect 112150 679700 112390 679940
rect 112500 679700 112740 679940
rect 112830 679700 113070 679940
rect 113160 679700 113400 679940
rect 113490 679700 113730 679940
rect 113840 679700 114080 679940
rect 114170 679700 114410 679940
rect 114500 679700 114740 679940
rect 114830 679700 115070 679940
rect 115180 679700 115420 679940
rect 115510 679700 115750 679940
rect 115840 679700 116080 679940
rect 116170 679700 116410 679940
rect 116520 679700 116760 679940
rect 116850 679700 117090 679940
rect 117180 679700 117420 679940
rect 117510 679700 117750 679940
rect 117860 679700 118100 679940
rect 118190 679700 118430 679940
rect 118520 679700 118760 679940
rect 118850 679700 119090 679940
rect 119200 679700 119440 679940
rect 119530 679700 119770 679940
rect 119860 679700 120100 679940
rect 120190 679700 120430 679940
rect 120540 679700 120780 679940
rect 120870 679700 121110 679940
rect 121200 679700 121440 679940
rect 121530 679700 121770 679940
rect 110810 679370 111050 679610
rect 111160 679370 111400 679610
rect 111490 679370 111730 679610
rect 111820 679370 112060 679610
rect 112150 679370 112390 679610
rect 112500 679370 112740 679610
rect 112830 679370 113070 679610
rect 113160 679370 113400 679610
rect 113490 679370 113730 679610
rect 113840 679370 114080 679610
rect 114170 679370 114410 679610
rect 114500 679370 114740 679610
rect 114830 679370 115070 679610
rect 115180 679370 115420 679610
rect 115510 679370 115750 679610
rect 115840 679370 116080 679610
rect 116170 679370 116410 679610
rect 116520 679370 116760 679610
rect 116850 679370 117090 679610
rect 117180 679370 117420 679610
rect 117510 679370 117750 679610
rect 117860 679370 118100 679610
rect 118190 679370 118430 679610
rect 118520 679370 118760 679610
rect 118850 679370 119090 679610
rect 119200 679370 119440 679610
rect 119530 679370 119770 679610
rect 119860 679370 120100 679610
rect 120190 679370 120430 679610
rect 120540 679370 120780 679610
rect 120870 679370 121110 679610
rect 121200 679370 121440 679610
rect 121530 679370 121770 679610
rect 110810 679020 111050 679260
rect 111160 679020 111400 679260
rect 111490 679020 111730 679260
rect 111820 679020 112060 679260
rect 112150 679020 112390 679260
rect 112500 679020 112740 679260
rect 112830 679020 113070 679260
rect 113160 679020 113400 679260
rect 113490 679020 113730 679260
rect 113840 679020 114080 679260
rect 114170 679020 114410 679260
rect 114500 679020 114740 679260
rect 114830 679020 115070 679260
rect 115180 679020 115420 679260
rect 115510 679020 115750 679260
rect 115840 679020 116080 679260
rect 116170 679020 116410 679260
rect 116520 679020 116760 679260
rect 116850 679020 117090 679260
rect 117180 679020 117420 679260
rect 117510 679020 117750 679260
rect 117860 679020 118100 679260
rect 118190 679020 118430 679260
rect 118520 679020 118760 679260
rect 118850 679020 119090 679260
rect 119200 679020 119440 679260
rect 119530 679020 119770 679260
rect 119860 679020 120100 679260
rect 120190 679020 120430 679260
rect 120540 679020 120780 679260
rect 120870 679020 121110 679260
rect 121200 679020 121440 679260
rect 121530 679020 121770 679260
rect 110810 678690 111050 678930
rect 111160 678690 111400 678930
rect 111490 678690 111730 678930
rect 111820 678690 112060 678930
rect 112150 678690 112390 678930
rect 112500 678690 112740 678930
rect 112830 678690 113070 678930
rect 113160 678690 113400 678930
rect 113490 678690 113730 678930
rect 113840 678690 114080 678930
rect 114170 678690 114410 678930
rect 114500 678690 114740 678930
rect 114830 678690 115070 678930
rect 115180 678690 115420 678930
rect 115510 678690 115750 678930
rect 115840 678690 116080 678930
rect 116170 678690 116410 678930
rect 116520 678690 116760 678930
rect 116850 678690 117090 678930
rect 117180 678690 117420 678930
rect 117510 678690 117750 678930
rect 117860 678690 118100 678930
rect 118190 678690 118430 678930
rect 118520 678690 118760 678930
rect 118850 678690 119090 678930
rect 119200 678690 119440 678930
rect 119530 678690 119770 678930
rect 119860 678690 120100 678930
rect 120190 678690 120430 678930
rect 120540 678690 120780 678930
rect 120870 678690 121110 678930
rect 121200 678690 121440 678930
rect 121530 678690 121770 678930
rect 110810 678360 111050 678600
rect 111160 678360 111400 678600
rect 111490 678360 111730 678600
rect 111820 678360 112060 678600
rect 112150 678360 112390 678600
rect 112500 678360 112740 678600
rect 112830 678360 113070 678600
rect 113160 678360 113400 678600
rect 113490 678360 113730 678600
rect 113840 678360 114080 678600
rect 114170 678360 114410 678600
rect 114500 678360 114740 678600
rect 114830 678360 115070 678600
rect 115180 678360 115420 678600
rect 115510 678360 115750 678600
rect 115840 678360 116080 678600
rect 116170 678360 116410 678600
rect 116520 678360 116760 678600
rect 116850 678360 117090 678600
rect 117180 678360 117420 678600
rect 117510 678360 117750 678600
rect 117860 678360 118100 678600
rect 118190 678360 118430 678600
rect 118520 678360 118760 678600
rect 118850 678360 119090 678600
rect 119200 678360 119440 678600
rect 119530 678360 119770 678600
rect 119860 678360 120100 678600
rect 120190 678360 120430 678600
rect 120540 678360 120780 678600
rect 120870 678360 121110 678600
rect 121200 678360 121440 678600
rect 121530 678360 121770 678600
rect 110810 678030 111050 678270
rect 111160 678030 111400 678270
rect 111490 678030 111730 678270
rect 111820 678030 112060 678270
rect 112150 678030 112390 678270
rect 112500 678030 112740 678270
rect 112830 678030 113070 678270
rect 113160 678030 113400 678270
rect 113490 678030 113730 678270
rect 113840 678030 114080 678270
rect 114170 678030 114410 678270
rect 114500 678030 114740 678270
rect 114830 678030 115070 678270
rect 115180 678030 115420 678270
rect 115510 678030 115750 678270
rect 115840 678030 116080 678270
rect 116170 678030 116410 678270
rect 116520 678030 116760 678270
rect 116850 678030 117090 678270
rect 117180 678030 117420 678270
rect 117510 678030 117750 678270
rect 117860 678030 118100 678270
rect 118190 678030 118430 678270
rect 118520 678030 118760 678270
rect 118850 678030 119090 678270
rect 119200 678030 119440 678270
rect 119530 678030 119770 678270
rect 119860 678030 120100 678270
rect 120190 678030 120430 678270
rect 120540 678030 120780 678270
rect 120870 678030 121110 678270
rect 121200 678030 121440 678270
rect 121530 678030 121770 678270
rect 110810 677680 111050 677920
rect 111160 677680 111400 677920
rect 111490 677680 111730 677920
rect 111820 677680 112060 677920
rect 112150 677680 112390 677920
rect 112500 677680 112740 677920
rect 112830 677680 113070 677920
rect 113160 677680 113400 677920
rect 113490 677680 113730 677920
rect 113840 677680 114080 677920
rect 114170 677680 114410 677920
rect 114500 677680 114740 677920
rect 114830 677680 115070 677920
rect 115180 677680 115420 677920
rect 115510 677680 115750 677920
rect 115840 677680 116080 677920
rect 116170 677680 116410 677920
rect 116520 677680 116760 677920
rect 116850 677680 117090 677920
rect 117180 677680 117420 677920
rect 117510 677680 117750 677920
rect 117860 677680 118100 677920
rect 118190 677680 118430 677920
rect 118520 677680 118760 677920
rect 118850 677680 119090 677920
rect 119200 677680 119440 677920
rect 119530 677680 119770 677920
rect 119860 677680 120100 677920
rect 120190 677680 120430 677920
rect 120540 677680 120780 677920
rect 120870 677680 121110 677920
rect 121200 677680 121440 677920
rect 121530 677680 121770 677920
rect 110810 677350 111050 677590
rect 111160 677350 111400 677590
rect 111490 677350 111730 677590
rect 111820 677350 112060 677590
rect 112150 677350 112390 677590
rect 112500 677350 112740 677590
rect 112830 677350 113070 677590
rect 113160 677350 113400 677590
rect 113490 677350 113730 677590
rect 113840 677350 114080 677590
rect 114170 677350 114410 677590
rect 114500 677350 114740 677590
rect 114830 677350 115070 677590
rect 115180 677350 115420 677590
rect 115510 677350 115750 677590
rect 115840 677350 116080 677590
rect 116170 677350 116410 677590
rect 116520 677350 116760 677590
rect 116850 677350 117090 677590
rect 117180 677350 117420 677590
rect 117510 677350 117750 677590
rect 117860 677350 118100 677590
rect 118190 677350 118430 677590
rect 118520 677350 118760 677590
rect 118850 677350 119090 677590
rect 119200 677350 119440 677590
rect 119530 677350 119770 677590
rect 119860 677350 120100 677590
rect 120190 677350 120430 677590
rect 120540 677350 120780 677590
rect 120870 677350 121110 677590
rect 121200 677350 121440 677590
rect 121530 677350 121770 677590
rect 110810 677020 111050 677260
rect 111160 677020 111400 677260
rect 111490 677020 111730 677260
rect 111820 677020 112060 677260
rect 112150 677020 112390 677260
rect 112500 677020 112740 677260
rect 112830 677020 113070 677260
rect 113160 677020 113400 677260
rect 113490 677020 113730 677260
rect 113840 677020 114080 677260
rect 114170 677020 114410 677260
rect 114500 677020 114740 677260
rect 114830 677020 115070 677260
rect 115180 677020 115420 677260
rect 115510 677020 115750 677260
rect 115840 677020 116080 677260
rect 116170 677020 116410 677260
rect 116520 677020 116760 677260
rect 116850 677020 117090 677260
rect 117180 677020 117420 677260
rect 117510 677020 117750 677260
rect 117860 677020 118100 677260
rect 118190 677020 118430 677260
rect 118520 677020 118760 677260
rect 118850 677020 119090 677260
rect 119200 677020 119440 677260
rect 119530 677020 119770 677260
rect 119860 677020 120100 677260
rect 120190 677020 120430 677260
rect 120540 677020 120780 677260
rect 120870 677020 121110 677260
rect 121200 677020 121440 677260
rect 121530 677020 121770 677260
rect 110810 676690 111050 676930
rect 111160 676690 111400 676930
rect 111490 676690 111730 676930
rect 111820 676690 112060 676930
rect 112150 676690 112390 676930
rect 112500 676690 112740 676930
rect 112830 676690 113070 676930
rect 113160 676690 113400 676930
rect 113490 676690 113730 676930
rect 113840 676690 114080 676930
rect 114170 676690 114410 676930
rect 114500 676690 114740 676930
rect 114830 676690 115070 676930
rect 115180 676690 115420 676930
rect 115510 676690 115750 676930
rect 115840 676690 116080 676930
rect 116170 676690 116410 676930
rect 116520 676690 116760 676930
rect 116850 676690 117090 676930
rect 117180 676690 117420 676930
rect 117510 676690 117750 676930
rect 117860 676690 118100 676930
rect 118190 676690 118430 676930
rect 118520 676690 118760 676930
rect 118850 676690 119090 676930
rect 119200 676690 119440 676930
rect 119530 676690 119770 676930
rect 119860 676690 120100 676930
rect 120190 676690 120430 676930
rect 120540 676690 120780 676930
rect 120870 676690 121110 676930
rect 121200 676690 121440 676930
rect 121530 676690 121770 676930
rect 110810 676340 111050 676580
rect 111160 676340 111400 676580
rect 111490 676340 111730 676580
rect 111820 676340 112060 676580
rect 112150 676340 112390 676580
rect 112500 676340 112740 676580
rect 112830 676340 113070 676580
rect 113160 676340 113400 676580
rect 113490 676340 113730 676580
rect 113840 676340 114080 676580
rect 114170 676340 114410 676580
rect 114500 676340 114740 676580
rect 114830 676340 115070 676580
rect 115180 676340 115420 676580
rect 115510 676340 115750 676580
rect 115840 676340 116080 676580
rect 116170 676340 116410 676580
rect 116520 676340 116760 676580
rect 116850 676340 117090 676580
rect 117180 676340 117420 676580
rect 117510 676340 117750 676580
rect 117860 676340 118100 676580
rect 118190 676340 118430 676580
rect 118520 676340 118760 676580
rect 118850 676340 119090 676580
rect 119200 676340 119440 676580
rect 119530 676340 119770 676580
rect 119860 676340 120100 676580
rect 120190 676340 120430 676580
rect 120540 676340 120780 676580
rect 120870 676340 121110 676580
rect 121200 676340 121440 676580
rect 121530 676340 121770 676580
rect 110810 676010 111050 676250
rect 111160 676010 111400 676250
rect 111490 676010 111730 676250
rect 111820 676010 112060 676250
rect 112150 676010 112390 676250
rect 112500 676010 112740 676250
rect 112830 676010 113070 676250
rect 113160 676010 113400 676250
rect 113490 676010 113730 676250
rect 113840 676010 114080 676250
rect 114170 676010 114410 676250
rect 114500 676010 114740 676250
rect 114830 676010 115070 676250
rect 115180 676010 115420 676250
rect 115510 676010 115750 676250
rect 115840 676010 116080 676250
rect 116170 676010 116410 676250
rect 116520 676010 116760 676250
rect 116850 676010 117090 676250
rect 117180 676010 117420 676250
rect 117510 676010 117750 676250
rect 117860 676010 118100 676250
rect 118190 676010 118430 676250
rect 118520 676010 118760 676250
rect 118850 676010 119090 676250
rect 119200 676010 119440 676250
rect 119530 676010 119770 676250
rect 119860 676010 120100 676250
rect 120190 676010 120430 676250
rect 120540 676010 120780 676250
rect 120870 676010 121110 676250
rect 121200 676010 121440 676250
rect 121530 676010 121770 676250
rect 110810 675680 111050 675920
rect 111160 675680 111400 675920
rect 111490 675680 111730 675920
rect 111820 675680 112060 675920
rect 112150 675680 112390 675920
rect 112500 675680 112740 675920
rect 112830 675680 113070 675920
rect 113160 675680 113400 675920
rect 113490 675680 113730 675920
rect 113840 675680 114080 675920
rect 114170 675680 114410 675920
rect 114500 675680 114740 675920
rect 114830 675680 115070 675920
rect 115180 675680 115420 675920
rect 115510 675680 115750 675920
rect 115840 675680 116080 675920
rect 116170 675680 116410 675920
rect 116520 675680 116760 675920
rect 116850 675680 117090 675920
rect 117180 675680 117420 675920
rect 117510 675680 117750 675920
rect 117860 675680 118100 675920
rect 118190 675680 118430 675920
rect 118520 675680 118760 675920
rect 118850 675680 119090 675920
rect 119200 675680 119440 675920
rect 119530 675680 119770 675920
rect 119860 675680 120100 675920
rect 120190 675680 120430 675920
rect 120540 675680 120780 675920
rect 120870 675680 121110 675920
rect 121200 675680 121440 675920
rect 121530 675680 121770 675920
rect 110810 675350 111050 675590
rect 111160 675350 111400 675590
rect 111490 675350 111730 675590
rect 111820 675350 112060 675590
rect 112150 675350 112390 675590
rect 112500 675350 112740 675590
rect 112830 675350 113070 675590
rect 113160 675350 113400 675590
rect 113490 675350 113730 675590
rect 113840 675350 114080 675590
rect 114170 675350 114410 675590
rect 114500 675350 114740 675590
rect 114830 675350 115070 675590
rect 115180 675350 115420 675590
rect 115510 675350 115750 675590
rect 115840 675350 116080 675590
rect 116170 675350 116410 675590
rect 116520 675350 116760 675590
rect 116850 675350 117090 675590
rect 117180 675350 117420 675590
rect 117510 675350 117750 675590
rect 117860 675350 118100 675590
rect 118190 675350 118430 675590
rect 118520 675350 118760 675590
rect 118850 675350 119090 675590
rect 119200 675350 119440 675590
rect 119530 675350 119770 675590
rect 119860 675350 120100 675590
rect 120190 675350 120430 675590
rect 120540 675350 120780 675590
rect 120870 675350 121110 675590
rect 121200 675350 121440 675590
rect 121530 675350 121770 675590
rect 110810 675000 111050 675240
rect 111160 675000 111400 675240
rect 111490 675000 111730 675240
rect 111820 675000 112060 675240
rect 112150 675000 112390 675240
rect 112500 675000 112740 675240
rect 112830 675000 113070 675240
rect 113160 675000 113400 675240
rect 113490 675000 113730 675240
rect 113840 675000 114080 675240
rect 114170 675000 114410 675240
rect 114500 675000 114740 675240
rect 114830 675000 115070 675240
rect 115180 675000 115420 675240
rect 115510 675000 115750 675240
rect 115840 675000 116080 675240
rect 116170 675000 116410 675240
rect 116520 675000 116760 675240
rect 116850 675000 117090 675240
rect 117180 675000 117420 675240
rect 117510 675000 117750 675240
rect 117860 675000 118100 675240
rect 118190 675000 118430 675240
rect 118520 675000 118760 675240
rect 118850 675000 119090 675240
rect 119200 675000 119440 675240
rect 119530 675000 119770 675240
rect 119860 675000 120100 675240
rect 120190 675000 120430 675240
rect 120540 675000 120780 675240
rect 120870 675000 121110 675240
rect 121200 675000 121440 675240
rect 121530 675000 121770 675240
rect 110810 674670 111050 674910
rect 111160 674670 111400 674910
rect 111490 674670 111730 674910
rect 111820 674670 112060 674910
rect 112150 674670 112390 674910
rect 112500 674670 112740 674910
rect 112830 674670 113070 674910
rect 113160 674670 113400 674910
rect 113490 674670 113730 674910
rect 113840 674670 114080 674910
rect 114170 674670 114410 674910
rect 114500 674670 114740 674910
rect 114830 674670 115070 674910
rect 115180 674670 115420 674910
rect 115510 674670 115750 674910
rect 115840 674670 116080 674910
rect 116170 674670 116410 674910
rect 116520 674670 116760 674910
rect 116850 674670 117090 674910
rect 117180 674670 117420 674910
rect 117510 674670 117750 674910
rect 117860 674670 118100 674910
rect 118190 674670 118430 674910
rect 118520 674670 118760 674910
rect 118850 674670 119090 674910
rect 119200 674670 119440 674910
rect 119530 674670 119770 674910
rect 119860 674670 120100 674910
rect 120190 674670 120430 674910
rect 120540 674670 120780 674910
rect 120870 674670 121110 674910
rect 121200 674670 121440 674910
rect 121530 674670 121770 674910
rect 110810 674340 111050 674580
rect 111160 674340 111400 674580
rect 111490 674340 111730 674580
rect 111820 674340 112060 674580
rect 112150 674340 112390 674580
rect 112500 674340 112740 674580
rect 112830 674340 113070 674580
rect 113160 674340 113400 674580
rect 113490 674340 113730 674580
rect 113840 674340 114080 674580
rect 114170 674340 114410 674580
rect 114500 674340 114740 674580
rect 114830 674340 115070 674580
rect 115180 674340 115420 674580
rect 115510 674340 115750 674580
rect 115840 674340 116080 674580
rect 116170 674340 116410 674580
rect 116520 674340 116760 674580
rect 116850 674340 117090 674580
rect 117180 674340 117420 674580
rect 117510 674340 117750 674580
rect 117860 674340 118100 674580
rect 118190 674340 118430 674580
rect 118520 674340 118760 674580
rect 118850 674340 119090 674580
rect 119200 674340 119440 674580
rect 119530 674340 119770 674580
rect 119860 674340 120100 674580
rect 120190 674340 120430 674580
rect 120540 674340 120780 674580
rect 120870 674340 121110 674580
rect 121200 674340 121440 674580
rect 121530 674340 121770 674580
rect 110810 674010 111050 674250
rect 111160 674010 111400 674250
rect 111490 674010 111730 674250
rect 111820 674010 112060 674250
rect 112150 674010 112390 674250
rect 112500 674010 112740 674250
rect 112830 674010 113070 674250
rect 113160 674010 113400 674250
rect 113490 674010 113730 674250
rect 113840 674010 114080 674250
rect 114170 674010 114410 674250
rect 114500 674010 114740 674250
rect 114830 674010 115070 674250
rect 115180 674010 115420 674250
rect 115510 674010 115750 674250
rect 115840 674010 116080 674250
rect 116170 674010 116410 674250
rect 116520 674010 116760 674250
rect 116850 674010 117090 674250
rect 117180 674010 117420 674250
rect 117510 674010 117750 674250
rect 117860 674010 118100 674250
rect 118190 674010 118430 674250
rect 118520 674010 118760 674250
rect 118850 674010 119090 674250
rect 119200 674010 119440 674250
rect 119530 674010 119770 674250
rect 119860 674010 120100 674250
rect 120190 674010 120430 674250
rect 120540 674010 120780 674250
rect 120870 674010 121110 674250
rect 121200 674010 121440 674250
rect 121530 674010 121770 674250
rect 110810 673660 111050 673900
rect 111160 673660 111400 673900
rect 111490 673660 111730 673900
rect 111820 673660 112060 673900
rect 112150 673660 112390 673900
rect 112500 673660 112740 673900
rect 112830 673660 113070 673900
rect 113160 673660 113400 673900
rect 113490 673660 113730 673900
rect 113840 673660 114080 673900
rect 114170 673660 114410 673900
rect 114500 673660 114740 673900
rect 114830 673660 115070 673900
rect 115180 673660 115420 673900
rect 115510 673660 115750 673900
rect 115840 673660 116080 673900
rect 116170 673660 116410 673900
rect 116520 673660 116760 673900
rect 116850 673660 117090 673900
rect 117180 673660 117420 673900
rect 117510 673660 117750 673900
rect 117860 673660 118100 673900
rect 118190 673660 118430 673900
rect 118520 673660 118760 673900
rect 118850 673660 119090 673900
rect 119200 673660 119440 673900
rect 119530 673660 119770 673900
rect 119860 673660 120100 673900
rect 120190 673660 120430 673900
rect 120540 673660 120780 673900
rect 120870 673660 121110 673900
rect 121200 673660 121440 673900
rect 121530 673660 121770 673900
rect 110810 673330 111050 673570
rect 111160 673330 111400 673570
rect 111490 673330 111730 673570
rect 111820 673330 112060 673570
rect 112150 673330 112390 673570
rect 112500 673330 112740 673570
rect 112830 673330 113070 673570
rect 113160 673330 113400 673570
rect 113490 673330 113730 673570
rect 113840 673330 114080 673570
rect 114170 673330 114410 673570
rect 114500 673330 114740 673570
rect 114830 673330 115070 673570
rect 115180 673330 115420 673570
rect 115510 673330 115750 673570
rect 115840 673330 116080 673570
rect 116170 673330 116410 673570
rect 116520 673330 116760 673570
rect 116850 673330 117090 673570
rect 117180 673330 117420 673570
rect 117510 673330 117750 673570
rect 117860 673330 118100 673570
rect 118190 673330 118430 673570
rect 118520 673330 118760 673570
rect 118850 673330 119090 673570
rect 119200 673330 119440 673570
rect 119530 673330 119770 673570
rect 119860 673330 120100 673570
rect 120190 673330 120430 673570
rect 120540 673330 120780 673570
rect 120870 673330 121110 673570
rect 121200 673330 121440 673570
rect 121530 673330 121770 673570
rect 110810 673000 111050 673240
rect 111160 673000 111400 673240
rect 111490 673000 111730 673240
rect 111820 673000 112060 673240
rect 112150 673000 112390 673240
rect 112500 673000 112740 673240
rect 112830 673000 113070 673240
rect 113160 673000 113400 673240
rect 113490 673000 113730 673240
rect 113840 673000 114080 673240
rect 114170 673000 114410 673240
rect 114500 673000 114740 673240
rect 114830 673000 115070 673240
rect 115180 673000 115420 673240
rect 115510 673000 115750 673240
rect 115840 673000 116080 673240
rect 116170 673000 116410 673240
rect 116520 673000 116760 673240
rect 116850 673000 117090 673240
rect 117180 673000 117420 673240
rect 117510 673000 117750 673240
rect 117860 673000 118100 673240
rect 118190 673000 118430 673240
rect 118520 673000 118760 673240
rect 118850 673000 119090 673240
rect 119200 673000 119440 673240
rect 119530 673000 119770 673240
rect 119860 673000 120100 673240
rect 120190 673000 120430 673240
rect 120540 673000 120780 673240
rect 120870 673000 121110 673240
rect 121200 673000 121440 673240
rect 121530 673000 121770 673240
rect 110810 672670 111050 672910
rect 111160 672670 111400 672910
rect 111490 672670 111730 672910
rect 111820 672670 112060 672910
rect 112150 672670 112390 672910
rect 112500 672670 112740 672910
rect 112830 672670 113070 672910
rect 113160 672670 113400 672910
rect 113490 672670 113730 672910
rect 113840 672670 114080 672910
rect 114170 672670 114410 672910
rect 114500 672670 114740 672910
rect 114830 672670 115070 672910
rect 115180 672670 115420 672910
rect 115510 672670 115750 672910
rect 115840 672670 116080 672910
rect 116170 672670 116410 672910
rect 116520 672670 116760 672910
rect 116850 672670 117090 672910
rect 117180 672670 117420 672910
rect 117510 672670 117750 672910
rect 117860 672670 118100 672910
rect 118190 672670 118430 672910
rect 118520 672670 118760 672910
rect 118850 672670 119090 672910
rect 119200 672670 119440 672910
rect 119530 672670 119770 672910
rect 119860 672670 120100 672910
rect 120190 672670 120430 672910
rect 120540 672670 120780 672910
rect 120870 672670 121110 672910
rect 121200 672670 121440 672910
rect 121530 672670 121770 672910
rect 110810 672320 111050 672560
rect 111160 672320 111400 672560
rect 111490 672320 111730 672560
rect 111820 672320 112060 672560
rect 112150 672320 112390 672560
rect 112500 672320 112740 672560
rect 112830 672320 113070 672560
rect 113160 672320 113400 672560
rect 113490 672320 113730 672560
rect 113840 672320 114080 672560
rect 114170 672320 114410 672560
rect 114500 672320 114740 672560
rect 114830 672320 115070 672560
rect 115180 672320 115420 672560
rect 115510 672320 115750 672560
rect 115840 672320 116080 672560
rect 116170 672320 116410 672560
rect 116520 672320 116760 672560
rect 116850 672320 117090 672560
rect 117180 672320 117420 672560
rect 117510 672320 117750 672560
rect 117860 672320 118100 672560
rect 118190 672320 118430 672560
rect 118520 672320 118760 672560
rect 118850 672320 119090 672560
rect 119200 672320 119440 672560
rect 119530 672320 119770 672560
rect 119860 672320 120100 672560
rect 120190 672320 120430 672560
rect 120540 672320 120780 672560
rect 120870 672320 121110 672560
rect 121200 672320 121440 672560
rect 121530 672320 121770 672560
rect 122190 683040 122430 683280
rect 122540 683040 122780 683280
rect 122870 683040 123110 683280
rect 123200 683040 123440 683280
rect 123530 683040 123770 683280
rect 123880 683040 124120 683280
rect 124210 683040 124450 683280
rect 124540 683040 124780 683280
rect 124870 683040 125110 683280
rect 125220 683040 125460 683280
rect 125550 683040 125790 683280
rect 125880 683040 126120 683280
rect 126210 683040 126450 683280
rect 126560 683040 126800 683280
rect 126890 683040 127130 683280
rect 127220 683040 127460 683280
rect 127550 683040 127790 683280
rect 127900 683040 128140 683280
rect 128230 683040 128470 683280
rect 128560 683040 128800 683280
rect 128890 683040 129130 683280
rect 129240 683040 129480 683280
rect 129570 683040 129810 683280
rect 129900 683040 130140 683280
rect 130230 683040 130470 683280
rect 130580 683040 130820 683280
rect 130910 683040 131150 683280
rect 131240 683040 131480 683280
rect 131570 683040 131810 683280
rect 131920 683040 132160 683280
rect 132250 683040 132490 683280
rect 132580 683040 132820 683280
rect 132910 683040 133150 683280
rect 122190 682710 122430 682950
rect 122540 682710 122780 682950
rect 122870 682710 123110 682950
rect 123200 682710 123440 682950
rect 123530 682710 123770 682950
rect 123880 682710 124120 682950
rect 124210 682710 124450 682950
rect 124540 682710 124780 682950
rect 124870 682710 125110 682950
rect 125220 682710 125460 682950
rect 125550 682710 125790 682950
rect 125880 682710 126120 682950
rect 126210 682710 126450 682950
rect 126560 682710 126800 682950
rect 126890 682710 127130 682950
rect 127220 682710 127460 682950
rect 127550 682710 127790 682950
rect 127900 682710 128140 682950
rect 128230 682710 128470 682950
rect 128560 682710 128800 682950
rect 128890 682710 129130 682950
rect 129240 682710 129480 682950
rect 129570 682710 129810 682950
rect 129900 682710 130140 682950
rect 130230 682710 130470 682950
rect 130580 682710 130820 682950
rect 130910 682710 131150 682950
rect 131240 682710 131480 682950
rect 131570 682710 131810 682950
rect 131920 682710 132160 682950
rect 132250 682710 132490 682950
rect 132580 682710 132820 682950
rect 132910 682710 133150 682950
rect 122190 682380 122430 682620
rect 122540 682380 122780 682620
rect 122870 682380 123110 682620
rect 123200 682380 123440 682620
rect 123530 682380 123770 682620
rect 123880 682380 124120 682620
rect 124210 682380 124450 682620
rect 124540 682380 124780 682620
rect 124870 682380 125110 682620
rect 125220 682380 125460 682620
rect 125550 682380 125790 682620
rect 125880 682380 126120 682620
rect 126210 682380 126450 682620
rect 126560 682380 126800 682620
rect 126890 682380 127130 682620
rect 127220 682380 127460 682620
rect 127550 682380 127790 682620
rect 127900 682380 128140 682620
rect 128230 682380 128470 682620
rect 128560 682380 128800 682620
rect 128890 682380 129130 682620
rect 129240 682380 129480 682620
rect 129570 682380 129810 682620
rect 129900 682380 130140 682620
rect 130230 682380 130470 682620
rect 130580 682380 130820 682620
rect 130910 682380 131150 682620
rect 131240 682380 131480 682620
rect 131570 682380 131810 682620
rect 131920 682380 132160 682620
rect 132250 682380 132490 682620
rect 132580 682380 132820 682620
rect 132910 682380 133150 682620
rect 122190 682050 122430 682290
rect 122540 682050 122780 682290
rect 122870 682050 123110 682290
rect 123200 682050 123440 682290
rect 123530 682050 123770 682290
rect 123880 682050 124120 682290
rect 124210 682050 124450 682290
rect 124540 682050 124780 682290
rect 124870 682050 125110 682290
rect 125220 682050 125460 682290
rect 125550 682050 125790 682290
rect 125880 682050 126120 682290
rect 126210 682050 126450 682290
rect 126560 682050 126800 682290
rect 126890 682050 127130 682290
rect 127220 682050 127460 682290
rect 127550 682050 127790 682290
rect 127900 682050 128140 682290
rect 128230 682050 128470 682290
rect 128560 682050 128800 682290
rect 128890 682050 129130 682290
rect 129240 682050 129480 682290
rect 129570 682050 129810 682290
rect 129900 682050 130140 682290
rect 130230 682050 130470 682290
rect 130580 682050 130820 682290
rect 130910 682050 131150 682290
rect 131240 682050 131480 682290
rect 131570 682050 131810 682290
rect 131920 682050 132160 682290
rect 132250 682050 132490 682290
rect 132580 682050 132820 682290
rect 132910 682050 133150 682290
rect 122190 681700 122430 681940
rect 122540 681700 122780 681940
rect 122870 681700 123110 681940
rect 123200 681700 123440 681940
rect 123530 681700 123770 681940
rect 123880 681700 124120 681940
rect 124210 681700 124450 681940
rect 124540 681700 124780 681940
rect 124870 681700 125110 681940
rect 125220 681700 125460 681940
rect 125550 681700 125790 681940
rect 125880 681700 126120 681940
rect 126210 681700 126450 681940
rect 126560 681700 126800 681940
rect 126890 681700 127130 681940
rect 127220 681700 127460 681940
rect 127550 681700 127790 681940
rect 127900 681700 128140 681940
rect 128230 681700 128470 681940
rect 128560 681700 128800 681940
rect 128890 681700 129130 681940
rect 129240 681700 129480 681940
rect 129570 681700 129810 681940
rect 129900 681700 130140 681940
rect 130230 681700 130470 681940
rect 130580 681700 130820 681940
rect 130910 681700 131150 681940
rect 131240 681700 131480 681940
rect 131570 681700 131810 681940
rect 131920 681700 132160 681940
rect 132250 681700 132490 681940
rect 132580 681700 132820 681940
rect 132910 681700 133150 681940
rect 122190 681370 122430 681610
rect 122540 681370 122780 681610
rect 122870 681370 123110 681610
rect 123200 681370 123440 681610
rect 123530 681370 123770 681610
rect 123880 681370 124120 681610
rect 124210 681370 124450 681610
rect 124540 681370 124780 681610
rect 124870 681370 125110 681610
rect 125220 681370 125460 681610
rect 125550 681370 125790 681610
rect 125880 681370 126120 681610
rect 126210 681370 126450 681610
rect 126560 681370 126800 681610
rect 126890 681370 127130 681610
rect 127220 681370 127460 681610
rect 127550 681370 127790 681610
rect 127900 681370 128140 681610
rect 128230 681370 128470 681610
rect 128560 681370 128800 681610
rect 128890 681370 129130 681610
rect 129240 681370 129480 681610
rect 129570 681370 129810 681610
rect 129900 681370 130140 681610
rect 130230 681370 130470 681610
rect 130580 681370 130820 681610
rect 130910 681370 131150 681610
rect 131240 681370 131480 681610
rect 131570 681370 131810 681610
rect 131920 681370 132160 681610
rect 132250 681370 132490 681610
rect 132580 681370 132820 681610
rect 132910 681370 133150 681610
rect 122190 681040 122430 681280
rect 122540 681040 122780 681280
rect 122870 681040 123110 681280
rect 123200 681040 123440 681280
rect 123530 681040 123770 681280
rect 123880 681040 124120 681280
rect 124210 681040 124450 681280
rect 124540 681040 124780 681280
rect 124870 681040 125110 681280
rect 125220 681040 125460 681280
rect 125550 681040 125790 681280
rect 125880 681040 126120 681280
rect 126210 681040 126450 681280
rect 126560 681040 126800 681280
rect 126890 681040 127130 681280
rect 127220 681040 127460 681280
rect 127550 681040 127790 681280
rect 127900 681040 128140 681280
rect 128230 681040 128470 681280
rect 128560 681040 128800 681280
rect 128890 681040 129130 681280
rect 129240 681040 129480 681280
rect 129570 681040 129810 681280
rect 129900 681040 130140 681280
rect 130230 681040 130470 681280
rect 130580 681040 130820 681280
rect 130910 681040 131150 681280
rect 131240 681040 131480 681280
rect 131570 681040 131810 681280
rect 131920 681040 132160 681280
rect 132250 681040 132490 681280
rect 132580 681040 132820 681280
rect 132910 681040 133150 681280
rect 122190 680710 122430 680950
rect 122540 680710 122780 680950
rect 122870 680710 123110 680950
rect 123200 680710 123440 680950
rect 123530 680710 123770 680950
rect 123880 680710 124120 680950
rect 124210 680710 124450 680950
rect 124540 680710 124780 680950
rect 124870 680710 125110 680950
rect 125220 680710 125460 680950
rect 125550 680710 125790 680950
rect 125880 680710 126120 680950
rect 126210 680710 126450 680950
rect 126560 680710 126800 680950
rect 126890 680710 127130 680950
rect 127220 680710 127460 680950
rect 127550 680710 127790 680950
rect 127900 680710 128140 680950
rect 128230 680710 128470 680950
rect 128560 680710 128800 680950
rect 128890 680710 129130 680950
rect 129240 680710 129480 680950
rect 129570 680710 129810 680950
rect 129900 680710 130140 680950
rect 130230 680710 130470 680950
rect 130580 680710 130820 680950
rect 130910 680710 131150 680950
rect 131240 680710 131480 680950
rect 131570 680710 131810 680950
rect 131920 680710 132160 680950
rect 132250 680710 132490 680950
rect 132580 680710 132820 680950
rect 132910 680710 133150 680950
rect 122190 680360 122430 680600
rect 122540 680360 122780 680600
rect 122870 680360 123110 680600
rect 123200 680360 123440 680600
rect 123530 680360 123770 680600
rect 123880 680360 124120 680600
rect 124210 680360 124450 680600
rect 124540 680360 124780 680600
rect 124870 680360 125110 680600
rect 125220 680360 125460 680600
rect 125550 680360 125790 680600
rect 125880 680360 126120 680600
rect 126210 680360 126450 680600
rect 126560 680360 126800 680600
rect 126890 680360 127130 680600
rect 127220 680360 127460 680600
rect 127550 680360 127790 680600
rect 127900 680360 128140 680600
rect 128230 680360 128470 680600
rect 128560 680360 128800 680600
rect 128890 680360 129130 680600
rect 129240 680360 129480 680600
rect 129570 680360 129810 680600
rect 129900 680360 130140 680600
rect 130230 680360 130470 680600
rect 130580 680360 130820 680600
rect 130910 680360 131150 680600
rect 131240 680360 131480 680600
rect 131570 680360 131810 680600
rect 131920 680360 132160 680600
rect 132250 680360 132490 680600
rect 132580 680360 132820 680600
rect 132910 680360 133150 680600
rect 122190 680030 122430 680270
rect 122540 680030 122780 680270
rect 122870 680030 123110 680270
rect 123200 680030 123440 680270
rect 123530 680030 123770 680270
rect 123880 680030 124120 680270
rect 124210 680030 124450 680270
rect 124540 680030 124780 680270
rect 124870 680030 125110 680270
rect 125220 680030 125460 680270
rect 125550 680030 125790 680270
rect 125880 680030 126120 680270
rect 126210 680030 126450 680270
rect 126560 680030 126800 680270
rect 126890 680030 127130 680270
rect 127220 680030 127460 680270
rect 127550 680030 127790 680270
rect 127900 680030 128140 680270
rect 128230 680030 128470 680270
rect 128560 680030 128800 680270
rect 128890 680030 129130 680270
rect 129240 680030 129480 680270
rect 129570 680030 129810 680270
rect 129900 680030 130140 680270
rect 130230 680030 130470 680270
rect 130580 680030 130820 680270
rect 130910 680030 131150 680270
rect 131240 680030 131480 680270
rect 131570 680030 131810 680270
rect 131920 680030 132160 680270
rect 132250 680030 132490 680270
rect 132580 680030 132820 680270
rect 132910 680030 133150 680270
rect 122190 679700 122430 679940
rect 122540 679700 122780 679940
rect 122870 679700 123110 679940
rect 123200 679700 123440 679940
rect 123530 679700 123770 679940
rect 123880 679700 124120 679940
rect 124210 679700 124450 679940
rect 124540 679700 124780 679940
rect 124870 679700 125110 679940
rect 125220 679700 125460 679940
rect 125550 679700 125790 679940
rect 125880 679700 126120 679940
rect 126210 679700 126450 679940
rect 126560 679700 126800 679940
rect 126890 679700 127130 679940
rect 127220 679700 127460 679940
rect 127550 679700 127790 679940
rect 127900 679700 128140 679940
rect 128230 679700 128470 679940
rect 128560 679700 128800 679940
rect 128890 679700 129130 679940
rect 129240 679700 129480 679940
rect 129570 679700 129810 679940
rect 129900 679700 130140 679940
rect 130230 679700 130470 679940
rect 130580 679700 130820 679940
rect 130910 679700 131150 679940
rect 131240 679700 131480 679940
rect 131570 679700 131810 679940
rect 131920 679700 132160 679940
rect 132250 679700 132490 679940
rect 132580 679700 132820 679940
rect 132910 679700 133150 679940
rect 122190 679370 122430 679610
rect 122540 679370 122780 679610
rect 122870 679370 123110 679610
rect 123200 679370 123440 679610
rect 123530 679370 123770 679610
rect 123880 679370 124120 679610
rect 124210 679370 124450 679610
rect 124540 679370 124780 679610
rect 124870 679370 125110 679610
rect 125220 679370 125460 679610
rect 125550 679370 125790 679610
rect 125880 679370 126120 679610
rect 126210 679370 126450 679610
rect 126560 679370 126800 679610
rect 126890 679370 127130 679610
rect 127220 679370 127460 679610
rect 127550 679370 127790 679610
rect 127900 679370 128140 679610
rect 128230 679370 128470 679610
rect 128560 679370 128800 679610
rect 128890 679370 129130 679610
rect 129240 679370 129480 679610
rect 129570 679370 129810 679610
rect 129900 679370 130140 679610
rect 130230 679370 130470 679610
rect 130580 679370 130820 679610
rect 130910 679370 131150 679610
rect 131240 679370 131480 679610
rect 131570 679370 131810 679610
rect 131920 679370 132160 679610
rect 132250 679370 132490 679610
rect 132580 679370 132820 679610
rect 132910 679370 133150 679610
rect 122190 679020 122430 679260
rect 122540 679020 122780 679260
rect 122870 679020 123110 679260
rect 123200 679020 123440 679260
rect 123530 679020 123770 679260
rect 123880 679020 124120 679260
rect 124210 679020 124450 679260
rect 124540 679020 124780 679260
rect 124870 679020 125110 679260
rect 125220 679020 125460 679260
rect 125550 679020 125790 679260
rect 125880 679020 126120 679260
rect 126210 679020 126450 679260
rect 126560 679020 126800 679260
rect 126890 679020 127130 679260
rect 127220 679020 127460 679260
rect 127550 679020 127790 679260
rect 127900 679020 128140 679260
rect 128230 679020 128470 679260
rect 128560 679020 128800 679260
rect 128890 679020 129130 679260
rect 129240 679020 129480 679260
rect 129570 679020 129810 679260
rect 129900 679020 130140 679260
rect 130230 679020 130470 679260
rect 130580 679020 130820 679260
rect 130910 679020 131150 679260
rect 131240 679020 131480 679260
rect 131570 679020 131810 679260
rect 131920 679020 132160 679260
rect 132250 679020 132490 679260
rect 132580 679020 132820 679260
rect 132910 679020 133150 679260
rect 122190 678690 122430 678930
rect 122540 678690 122780 678930
rect 122870 678690 123110 678930
rect 123200 678690 123440 678930
rect 123530 678690 123770 678930
rect 123880 678690 124120 678930
rect 124210 678690 124450 678930
rect 124540 678690 124780 678930
rect 124870 678690 125110 678930
rect 125220 678690 125460 678930
rect 125550 678690 125790 678930
rect 125880 678690 126120 678930
rect 126210 678690 126450 678930
rect 126560 678690 126800 678930
rect 126890 678690 127130 678930
rect 127220 678690 127460 678930
rect 127550 678690 127790 678930
rect 127900 678690 128140 678930
rect 128230 678690 128470 678930
rect 128560 678690 128800 678930
rect 128890 678690 129130 678930
rect 129240 678690 129480 678930
rect 129570 678690 129810 678930
rect 129900 678690 130140 678930
rect 130230 678690 130470 678930
rect 130580 678690 130820 678930
rect 130910 678690 131150 678930
rect 131240 678690 131480 678930
rect 131570 678690 131810 678930
rect 131920 678690 132160 678930
rect 132250 678690 132490 678930
rect 132580 678690 132820 678930
rect 132910 678690 133150 678930
rect 122190 678360 122430 678600
rect 122540 678360 122780 678600
rect 122870 678360 123110 678600
rect 123200 678360 123440 678600
rect 123530 678360 123770 678600
rect 123880 678360 124120 678600
rect 124210 678360 124450 678600
rect 124540 678360 124780 678600
rect 124870 678360 125110 678600
rect 125220 678360 125460 678600
rect 125550 678360 125790 678600
rect 125880 678360 126120 678600
rect 126210 678360 126450 678600
rect 126560 678360 126800 678600
rect 126890 678360 127130 678600
rect 127220 678360 127460 678600
rect 127550 678360 127790 678600
rect 127900 678360 128140 678600
rect 128230 678360 128470 678600
rect 128560 678360 128800 678600
rect 128890 678360 129130 678600
rect 129240 678360 129480 678600
rect 129570 678360 129810 678600
rect 129900 678360 130140 678600
rect 130230 678360 130470 678600
rect 130580 678360 130820 678600
rect 130910 678360 131150 678600
rect 131240 678360 131480 678600
rect 131570 678360 131810 678600
rect 131920 678360 132160 678600
rect 132250 678360 132490 678600
rect 132580 678360 132820 678600
rect 132910 678360 133150 678600
rect 122190 678030 122430 678270
rect 122540 678030 122780 678270
rect 122870 678030 123110 678270
rect 123200 678030 123440 678270
rect 123530 678030 123770 678270
rect 123880 678030 124120 678270
rect 124210 678030 124450 678270
rect 124540 678030 124780 678270
rect 124870 678030 125110 678270
rect 125220 678030 125460 678270
rect 125550 678030 125790 678270
rect 125880 678030 126120 678270
rect 126210 678030 126450 678270
rect 126560 678030 126800 678270
rect 126890 678030 127130 678270
rect 127220 678030 127460 678270
rect 127550 678030 127790 678270
rect 127900 678030 128140 678270
rect 128230 678030 128470 678270
rect 128560 678030 128800 678270
rect 128890 678030 129130 678270
rect 129240 678030 129480 678270
rect 129570 678030 129810 678270
rect 129900 678030 130140 678270
rect 130230 678030 130470 678270
rect 130580 678030 130820 678270
rect 130910 678030 131150 678270
rect 131240 678030 131480 678270
rect 131570 678030 131810 678270
rect 131920 678030 132160 678270
rect 132250 678030 132490 678270
rect 132580 678030 132820 678270
rect 132910 678030 133150 678270
rect 122190 677680 122430 677920
rect 122540 677680 122780 677920
rect 122870 677680 123110 677920
rect 123200 677680 123440 677920
rect 123530 677680 123770 677920
rect 123880 677680 124120 677920
rect 124210 677680 124450 677920
rect 124540 677680 124780 677920
rect 124870 677680 125110 677920
rect 125220 677680 125460 677920
rect 125550 677680 125790 677920
rect 125880 677680 126120 677920
rect 126210 677680 126450 677920
rect 126560 677680 126800 677920
rect 126890 677680 127130 677920
rect 127220 677680 127460 677920
rect 127550 677680 127790 677920
rect 127900 677680 128140 677920
rect 128230 677680 128470 677920
rect 128560 677680 128800 677920
rect 128890 677680 129130 677920
rect 129240 677680 129480 677920
rect 129570 677680 129810 677920
rect 129900 677680 130140 677920
rect 130230 677680 130470 677920
rect 130580 677680 130820 677920
rect 130910 677680 131150 677920
rect 131240 677680 131480 677920
rect 131570 677680 131810 677920
rect 131920 677680 132160 677920
rect 132250 677680 132490 677920
rect 132580 677680 132820 677920
rect 132910 677680 133150 677920
rect 122190 677350 122430 677590
rect 122540 677350 122780 677590
rect 122870 677350 123110 677590
rect 123200 677350 123440 677590
rect 123530 677350 123770 677590
rect 123880 677350 124120 677590
rect 124210 677350 124450 677590
rect 124540 677350 124780 677590
rect 124870 677350 125110 677590
rect 125220 677350 125460 677590
rect 125550 677350 125790 677590
rect 125880 677350 126120 677590
rect 126210 677350 126450 677590
rect 126560 677350 126800 677590
rect 126890 677350 127130 677590
rect 127220 677350 127460 677590
rect 127550 677350 127790 677590
rect 127900 677350 128140 677590
rect 128230 677350 128470 677590
rect 128560 677350 128800 677590
rect 128890 677350 129130 677590
rect 129240 677350 129480 677590
rect 129570 677350 129810 677590
rect 129900 677350 130140 677590
rect 130230 677350 130470 677590
rect 130580 677350 130820 677590
rect 130910 677350 131150 677590
rect 131240 677350 131480 677590
rect 131570 677350 131810 677590
rect 131920 677350 132160 677590
rect 132250 677350 132490 677590
rect 132580 677350 132820 677590
rect 132910 677350 133150 677590
rect 122190 677020 122430 677260
rect 122540 677020 122780 677260
rect 122870 677020 123110 677260
rect 123200 677020 123440 677260
rect 123530 677020 123770 677260
rect 123880 677020 124120 677260
rect 124210 677020 124450 677260
rect 124540 677020 124780 677260
rect 124870 677020 125110 677260
rect 125220 677020 125460 677260
rect 125550 677020 125790 677260
rect 125880 677020 126120 677260
rect 126210 677020 126450 677260
rect 126560 677020 126800 677260
rect 126890 677020 127130 677260
rect 127220 677020 127460 677260
rect 127550 677020 127790 677260
rect 127900 677020 128140 677260
rect 128230 677020 128470 677260
rect 128560 677020 128800 677260
rect 128890 677020 129130 677260
rect 129240 677020 129480 677260
rect 129570 677020 129810 677260
rect 129900 677020 130140 677260
rect 130230 677020 130470 677260
rect 130580 677020 130820 677260
rect 130910 677020 131150 677260
rect 131240 677020 131480 677260
rect 131570 677020 131810 677260
rect 131920 677020 132160 677260
rect 132250 677020 132490 677260
rect 132580 677020 132820 677260
rect 132910 677020 133150 677260
rect 122190 676690 122430 676930
rect 122540 676690 122780 676930
rect 122870 676690 123110 676930
rect 123200 676690 123440 676930
rect 123530 676690 123770 676930
rect 123880 676690 124120 676930
rect 124210 676690 124450 676930
rect 124540 676690 124780 676930
rect 124870 676690 125110 676930
rect 125220 676690 125460 676930
rect 125550 676690 125790 676930
rect 125880 676690 126120 676930
rect 126210 676690 126450 676930
rect 126560 676690 126800 676930
rect 126890 676690 127130 676930
rect 127220 676690 127460 676930
rect 127550 676690 127790 676930
rect 127900 676690 128140 676930
rect 128230 676690 128470 676930
rect 128560 676690 128800 676930
rect 128890 676690 129130 676930
rect 129240 676690 129480 676930
rect 129570 676690 129810 676930
rect 129900 676690 130140 676930
rect 130230 676690 130470 676930
rect 130580 676690 130820 676930
rect 130910 676690 131150 676930
rect 131240 676690 131480 676930
rect 131570 676690 131810 676930
rect 131920 676690 132160 676930
rect 132250 676690 132490 676930
rect 132580 676690 132820 676930
rect 132910 676690 133150 676930
rect 122190 676340 122430 676580
rect 122540 676340 122780 676580
rect 122870 676340 123110 676580
rect 123200 676340 123440 676580
rect 123530 676340 123770 676580
rect 123880 676340 124120 676580
rect 124210 676340 124450 676580
rect 124540 676340 124780 676580
rect 124870 676340 125110 676580
rect 125220 676340 125460 676580
rect 125550 676340 125790 676580
rect 125880 676340 126120 676580
rect 126210 676340 126450 676580
rect 126560 676340 126800 676580
rect 126890 676340 127130 676580
rect 127220 676340 127460 676580
rect 127550 676340 127790 676580
rect 127900 676340 128140 676580
rect 128230 676340 128470 676580
rect 128560 676340 128800 676580
rect 128890 676340 129130 676580
rect 129240 676340 129480 676580
rect 129570 676340 129810 676580
rect 129900 676340 130140 676580
rect 130230 676340 130470 676580
rect 130580 676340 130820 676580
rect 130910 676340 131150 676580
rect 131240 676340 131480 676580
rect 131570 676340 131810 676580
rect 131920 676340 132160 676580
rect 132250 676340 132490 676580
rect 132580 676340 132820 676580
rect 132910 676340 133150 676580
rect 122190 676010 122430 676250
rect 122540 676010 122780 676250
rect 122870 676010 123110 676250
rect 123200 676010 123440 676250
rect 123530 676010 123770 676250
rect 123880 676010 124120 676250
rect 124210 676010 124450 676250
rect 124540 676010 124780 676250
rect 124870 676010 125110 676250
rect 125220 676010 125460 676250
rect 125550 676010 125790 676250
rect 125880 676010 126120 676250
rect 126210 676010 126450 676250
rect 126560 676010 126800 676250
rect 126890 676010 127130 676250
rect 127220 676010 127460 676250
rect 127550 676010 127790 676250
rect 127900 676010 128140 676250
rect 128230 676010 128470 676250
rect 128560 676010 128800 676250
rect 128890 676010 129130 676250
rect 129240 676010 129480 676250
rect 129570 676010 129810 676250
rect 129900 676010 130140 676250
rect 130230 676010 130470 676250
rect 130580 676010 130820 676250
rect 130910 676010 131150 676250
rect 131240 676010 131480 676250
rect 131570 676010 131810 676250
rect 131920 676010 132160 676250
rect 132250 676010 132490 676250
rect 132580 676010 132820 676250
rect 132910 676010 133150 676250
rect 122190 675680 122430 675920
rect 122540 675680 122780 675920
rect 122870 675680 123110 675920
rect 123200 675680 123440 675920
rect 123530 675680 123770 675920
rect 123880 675680 124120 675920
rect 124210 675680 124450 675920
rect 124540 675680 124780 675920
rect 124870 675680 125110 675920
rect 125220 675680 125460 675920
rect 125550 675680 125790 675920
rect 125880 675680 126120 675920
rect 126210 675680 126450 675920
rect 126560 675680 126800 675920
rect 126890 675680 127130 675920
rect 127220 675680 127460 675920
rect 127550 675680 127790 675920
rect 127900 675680 128140 675920
rect 128230 675680 128470 675920
rect 128560 675680 128800 675920
rect 128890 675680 129130 675920
rect 129240 675680 129480 675920
rect 129570 675680 129810 675920
rect 129900 675680 130140 675920
rect 130230 675680 130470 675920
rect 130580 675680 130820 675920
rect 130910 675680 131150 675920
rect 131240 675680 131480 675920
rect 131570 675680 131810 675920
rect 131920 675680 132160 675920
rect 132250 675680 132490 675920
rect 132580 675680 132820 675920
rect 132910 675680 133150 675920
rect 122190 675350 122430 675590
rect 122540 675350 122780 675590
rect 122870 675350 123110 675590
rect 123200 675350 123440 675590
rect 123530 675350 123770 675590
rect 123880 675350 124120 675590
rect 124210 675350 124450 675590
rect 124540 675350 124780 675590
rect 124870 675350 125110 675590
rect 125220 675350 125460 675590
rect 125550 675350 125790 675590
rect 125880 675350 126120 675590
rect 126210 675350 126450 675590
rect 126560 675350 126800 675590
rect 126890 675350 127130 675590
rect 127220 675350 127460 675590
rect 127550 675350 127790 675590
rect 127900 675350 128140 675590
rect 128230 675350 128470 675590
rect 128560 675350 128800 675590
rect 128890 675350 129130 675590
rect 129240 675350 129480 675590
rect 129570 675350 129810 675590
rect 129900 675350 130140 675590
rect 130230 675350 130470 675590
rect 130580 675350 130820 675590
rect 130910 675350 131150 675590
rect 131240 675350 131480 675590
rect 131570 675350 131810 675590
rect 131920 675350 132160 675590
rect 132250 675350 132490 675590
rect 132580 675350 132820 675590
rect 132910 675350 133150 675590
rect 122190 675000 122430 675240
rect 122540 675000 122780 675240
rect 122870 675000 123110 675240
rect 123200 675000 123440 675240
rect 123530 675000 123770 675240
rect 123880 675000 124120 675240
rect 124210 675000 124450 675240
rect 124540 675000 124780 675240
rect 124870 675000 125110 675240
rect 125220 675000 125460 675240
rect 125550 675000 125790 675240
rect 125880 675000 126120 675240
rect 126210 675000 126450 675240
rect 126560 675000 126800 675240
rect 126890 675000 127130 675240
rect 127220 675000 127460 675240
rect 127550 675000 127790 675240
rect 127900 675000 128140 675240
rect 128230 675000 128470 675240
rect 128560 675000 128800 675240
rect 128890 675000 129130 675240
rect 129240 675000 129480 675240
rect 129570 675000 129810 675240
rect 129900 675000 130140 675240
rect 130230 675000 130470 675240
rect 130580 675000 130820 675240
rect 130910 675000 131150 675240
rect 131240 675000 131480 675240
rect 131570 675000 131810 675240
rect 131920 675000 132160 675240
rect 132250 675000 132490 675240
rect 132580 675000 132820 675240
rect 132910 675000 133150 675240
rect 122190 674670 122430 674910
rect 122540 674670 122780 674910
rect 122870 674670 123110 674910
rect 123200 674670 123440 674910
rect 123530 674670 123770 674910
rect 123880 674670 124120 674910
rect 124210 674670 124450 674910
rect 124540 674670 124780 674910
rect 124870 674670 125110 674910
rect 125220 674670 125460 674910
rect 125550 674670 125790 674910
rect 125880 674670 126120 674910
rect 126210 674670 126450 674910
rect 126560 674670 126800 674910
rect 126890 674670 127130 674910
rect 127220 674670 127460 674910
rect 127550 674670 127790 674910
rect 127900 674670 128140 674910
rect 128230 674670 128470 674910
rect 128560 674670 128800 674910
rect 128890 674670 129130 674910
rect 129240 674670 129480 674910
rect 129570 674670 129810 674910
rect 129900 674670 130140 674910
rect 130230 674670 130470 674910
rect 130580 674670 130820 674910
rect 130910 674670 131150 674910
rect 131240 674670 131480 674910
rect 131570 674670 131810 674910
rect 131920 674670 132160 674910
rect 132250 674670 132490 674910
rect 132580 674670 132820 674910
rect 132910 674670 133150 674910
rect 122190 674340 122430 674580
rect 122540 674340 122780 674580
rect 122870 674340 123110 674580
rect 123200 674340 123440 674580
rect 123530 674340 123770 674580
rect 123880 674340 124120 674580
rect 124210 674340 124450 674580
rect 124540 674340 124780 674580
rect 124870 674340 125110 674580
rect 125220 674340 125460 674580
rect 125550 674340 125790 674580
rect 125880 674340 126120 674580
rect 126210 674340 126450 674580
rect 126560 674340 126800 674580
rect 126890 674340 127130 674580
rect 127220 674340 127460 674580
rect 127550 674340 127790 674580
rect 127900 674340 128140 674580
rect 128230 674340 128470 674580
rect 128560 674340 128800 674580
rect 128890 674340 129130 674580
rect 129240 674340 129480 674580
rect 129570 674340 129810 674580
rect 129900 674340 130140 674580
rect 130230 674340 130470 674580
rect 130580 674340 130820 674580
rect 130910 674340 131150 674580
rect 131240 674340 131480 674580
rect 131570 674340 131810 674580
rect 131920 674340 132160 674580
rect 132250 674340 132490 674580
rect 132580 674340 132820 674580
rect 132910 674340 133150 674580
rect 122190 674010 122430 674250
rect 122540 674010 122780 674250
rect 122870 674010 123110 674250
rect 123200 674010 123440 674250
rect 123530 674010 123770 674250
rect 123880 674010 124120 674250
rect 124210 674010 124450 674250
rect 124540 674010 124780 674250
rect 124870 674010 125110 674250
rect 125220 674010 125460 674250
rect 125550 674010 125790 674250
rect 125880 674010 126120 674250
rect 126210 674010 126450 674250
rect 126560 674010 126800 674250
rect 126890 674010 127130 674250
rect 127220 674010 127460 674250
rect 127550 674010 127790 674250
rect 127900 674010 128140 674250
rect 128230 674010 128470 674250
rect 128560 674010 128800 674250
rect 128890 674010 129130 674250
rect 129240 674010 129480 674250
rect 129570 674010 129810 674250
rect 129900 674010 130140 674250
rect 130230 674010 130470 674250
rect 130580 674010 130820 674250
rect 130910 674010 131150 674250
rect 131240 674010 131480 674250
rect 131570 674010 131810 674250
rect 131920 674010 132160 674250
rect 132250 674010 132490 674250
rect 132580 674010 132820 674250
rect 132910 674010 133150 674250
rect 122190 673660 122430 673900
rect 122540 673660 122780 673900
rect 122870 673660 123110 673900
rect 123200 673660 123440 673900
rect 123530 673660 123770 673900
rect 123880 673660 124120 673900
rect 124210 673660 124450 673900
rect 124540 673660 124780 673900
rect 124870 673660 125110 673900
rect 125220 673660 125460 673900
rect 125550 673660 125790 673900
rect 125880 673660 126120 673900
rect 126210 673660 126450 673900
rect 126560 673660 126800 673900
rect 126890 673660 127130 673900
rect 127220 673660 127460 673900
rect 127550 673660 127790 673900
rect 127900 673660 128140 673900
rect 128230 673660 128470 673900
rect 128560 673660 128800 673900
rect 128890 673660 129130 673900
rect 129240 673660 129480 673900
rect 129570 673660 129810 673900
rect 129900 673660 130140 673900
rect 130230 673660 130470 673900
rect 130580 673660 130820 673900
rect 130910 673660 131150 673900
rect 131240 673660 131480 673900
rect 131570 673660 131810 673900
rect 131920 673660 132160 673900
rect 132250 673660 132490 673900
rect 132580 673660 132820 673900
rect 132910 673660 133150 673900
rect 122190 673330 122430 673570
rect 122540 673330 122780 673570
rect 122870 673330 123110 673570
rect 123200 673330 123440 673570
rect 123530 673330 123770 673570
rect 123880 673330 124120 673570
rect 124210 673330 124450 673570
rect 124540 673330 124780 673570
rect 124870 673330 125110 673570
rect 125220 673330 125460 673570
rect 125550 673330 125790 673570
rect 125880 673330 126120 673570
rect 126210 673330 126450 673570
rect 126560 673330 126800 673570
rect 126890 673330 127130 673570
rect 127220 673330 127460 673570
rect 127550 673330 127790 673570
rect 127900 673330 128140 673570
rect 128230 673330 128470 673570
rect 128560 673330 128800 673570
rect 128890 673330 129130 673570
rect 129240 673330 129480 673570
rect 129570 673330 129810 673570
rect 129900 673330 130140 673570
rect 130230 673330 130470 673570
rect 130580 673330 130820 673570
rect 130910 673330 131150 673570
rect 131240 673330 131480 673570
rect 131570 673330 131810 673570
rect 131920 673330 132160 673570
rect 132250 673330 132490 673570
rect 132580 673330 132820 673570
rect 132910 673330 133150 673570
rect 122190 673000 122430 673240
rect 122540 673000 122780 673240
rect 122870 673000 123110 673240
rect 123200 673000 123440 673240
rect 123530 673000 123770 673240
rect 123880 673000 124120 673240
rect 124210 673000 124450 673240
rect 124540 673000 124780 673240
rect 124870 673000 125110 673240
rect 125220 673000 125460 673240
rect 125550 673000 125790 673240
rect 125880 673000 126120 673240
rect 126210 673000 126450 673240
rect 126560 673000 126800 673240
rect 126890 673000 127130 673240
rect 127220 673000 127460 673240
rect 127550 673000 127790 673240
rect 127900 673000 128140 673240
rect 128230 673000 128470 673240
rect 128560 673000 128800 673240
rect 128890 673000 129130 673240
rect 129240 673000 129480 673240
rect 129570 673000 129810 673240
rect 129900 673000 130140 673240
rect 130230 673000 130470 673240
rect 130580 673000 130820 673240
rect 130910 673000 131150 673240
rect 131240 673000 131480 673240
rect 131570 673000 131810 673240
rect 131920 673000 132160 673240
rect 132250 673000 132490 673240
rect 132580 673000 132820 673240
rect 132910 673000 133150 673240
rect 122190 672670 122430 672910
rect 122540 672670 122780 672910
rect 122870 672670 123110 672910
rect 123200 672670 123440 672910
rect 123530 672670 123770 672910
rect 123880 672670 124120 672910
rect 124210 672670 124450 672910
rect 124540 672670 124780 672910
rect 124870 672670 125110 672910
rect 125220 672670 125460 672910
rect 125550 672670 125790 672910
rect 125880 672670 126120 672910
rect 126210 672670 126450 672910
rect 126560 672670 126800 672910
rect 126890 672670 127130 672910
rect 127220 672670 127460 672910
rect 127550 672670 127790 672910
rect 127900 672670 128140 672910
rect 128230 672670 128470 672910
rect 128560 672670 128800 672910
rect 128890 672670 129130 672910
rect 129240 672670 129480 672910
rect 129570 672670 129810 672910
rect 129900 672670 130140 672910
rect 130230 672670 130470 672910
rect 130580 672670 130820 672910
rect 130910 672670 131150 672910
rect 131240 672670 131480 672910
rect 131570 672670 131810 672910
rect 131920 672670 132160 672910
rect 132250 672670 132490 672910
rect 132580 672670 132820 672910
rect 132910 672670 133150 672910
rect 122190 672320 122430 672560
rect 122540 672320 122780 672560
rect 122870 672320 123110 672560
rect 123200 672320 123440 672560
rect 123530 672320 123770 672560
rect 123880 672320 124120 672560
rect 124210 672320 124450 672560
rect 124540 672320 124780 672560
rect 124870 672320 125110 672560
rect 125220 672320 125460 672560
rect 125550 672320 125790 672560
rect 125880 672320 126120 672560
rect 126210 672320 126450 672560
rect 126560 672320 126800 672560
rect 126890 672320 127130 672560
rect 127220 672320 127460 672560
rect 127550 672320 127790 672560
rect 127900 672320 128140 672560
rect 128230 672320 128470 672560
rect 128560 672320 128800 672560
rect 128890 672320 129130 672560
rect 129240 672320 129480 672560
rect 129570 672320 129810 672560
rect 129900 672320 130140 672560
rect 130230 672320 130470 672560
rect 130580 672320 130820 672560
rect 130910 672320 131150 672560
rect 131240 672320 131480 672560
rect 131570 672320 131810 672560
rect 131920 672320 132160 672560
rect 132250 672320 132490 672560
rect 132580 672320 132820 672560
rect 132910 672320 133150 672560
rect 133570 683040 133810 683280
rect 133920 683040 134160 683280
rect 134250 683040 134490 683280
rect 134580 683040 134820 683280
rect 134910 683040 135150 683280
rect 135260 683040 135500 683280
rect 135590 683040 135830 683280
rect 135920 683040 136160 683280
rect 136250 683040 136490 683280
rect 136600 683040 136840 683280
rect 136930 683040 137170 683280
rect 137260 683040 137500 683280
rect 137590 683040 137830 683280
rect 137940 683040 138180 683280
rect 138270 683040 138510 683280
rect 138600 683040 138840 683280
rect 138930 683040 139170 683280
rect 139280 683040 139520 683280
rect 139610 683040 139850 683280
rect 139940 683040 140180 683280
rect 140270 683040 140510 683280
rect 140620 683040 140860 683280
rect 140950 683040 141190 683280
rect 141280 683040 141520 683280
rect 141610 683040 141850 683280
rect 141960 683040 142200 683280
rect 142290 683040 142530 683280
rect 142620 683040 142860 683280
rect 142950 683040 143190 683280
rect 143300 683040 143540 683280
rect 143630 683040 143870 683280
rect 143960 683040 144200 683280
rect 144290 683040 144530 683280
rect 133570 682710 133810 682950
rect 133920 682710 134160 682950
rect 134250 682710 134490 682950
rect 134580 682710 134820 682950
rect 134910 682710 135150 682950
rect 135260 682710 135500 682950
rect 135590 682710 135830 682950
rect 135920 682710 136160 682950
rect 136250 682710 136490 682950
rect 136600 682710 136840 682950
rect 136930 682710 137170 682950
rect 137260 682710 137500 682950
rect 137590 682710 137830 682950
rect 137940 682710 138180 682950
rect 138270 682710 138510 682950
rect 138600 682710 138840 682950
rect 138930 682710 139170 682950
rect 139280 682710 139520 682950
rect 139610 682710 139850 682950
rect 139940 682710 140180 682950
rect 140270 682710 140510 682950
rect 140620 682710 140860 682950
rect 140950 682710 141190 682950
rect 141280 682710 141520 682950
rect 141610 682710 141850 682950
rect 141960 682710 142200 682950
rect 142290 682710 142530 682950
rect 142620 682710 142860 682950
rect 142950 682710 143190 682950
rect 143300 682710 143540 682950
rect 143630 682710 143870 682950
rect 143960 682710 144200 682950
rect 144290 682710 144530 682950
rect 133570 682380 133810 682620
rect 133920 682380 134160 682620
rect 134250 682380 134490 682620
rect 134580 682380 134820 682620
rect 134910 682380 135150 682620
rect 135260 682380 135500 682620
rect 135590 682380 135830 682620
rect 135920 682380 136160 682620
rect 136250 682380 136490 682620
rect 136600 682380 136840 682620
rect 136930 682380 137170 682620
rect 137260 682380 137500 682620
rect 137590 682380 137830 682620
rect 137940 682380 138180 682620
rect 138270 682380 138510 682620
rect 138600 682380 138840 682620
rect 138930 682380 139170 682620
rect 139280 682380 139520 682620
rect 139610 682380 139850 682620
rect 139940 682380 140180 682620
rect 140270 682380 140510 682620
rect 140620 682380 140860 682620
rect 140950 682380 141190 682620
rect 141280 682380 141520 682620
rect 141610 682380 141850 682620
rect 141960 682380 142200 682620
rect 142290 682380 142530 682620
rect 142620 682380 142860 682620
rect 142950 682380 143190 682620
rect 143300 682380 143540 682620
rect 143630 682380 143870 682620
rect 143960 682380 144200 682620
rect 144290 682380 144530 682620
rect 133570 682050 133810 682290
rect 133920 682050 134160 682290
rect 134250 682050 134490 682290
rect 134580 682050 134820 682290
rect 134910 682050 135150 682290
rect 135260 682050 135500 682290
rect 135590 682050 135830 682290
rect 135920 682050 136160 682290
rect 136250 682050 136490 682290
rect 136600 682050 136840 682290
rect 136930 682050 137170 682290
rect 137260 682050 137500 682290
rect 137590 682050 137830 682290
rect 137940 682050 138180 682290
rect 138270 682050 138510 682290
rect 138600 682050 138840 682290
rect 138930 682050 139170 682290
rect 139280 682050 139520 682290
rect 139610 682050 139850 682290
rect 139940 682050 140180 682290
rect 140270 682050 140510 682290
rect 140620 682050 140860 682290
rect 140950 682050 141190 682290
rect 141280 682050 141520 682290
rect 141610 682050 141850 682290
rect 141960 682050 142200 682290
rect 142290 682050 142530 682290
rect 142620 682050 142860 682290
rect 142950 682050 143190 682290
rect 143300 682050 143540 682290
rect 143630 682050 143870 682290
rect 143960 682050 144200 682290
rect 144290 682050 144530 682290
rect 133570 681700 133810 681940
rect 133920 681700 134160 681940
rect 134250 681700 134490 681940
rect 134580 681700 134820 681940
rect 134910 681700 135150 681940
rect 135260 681700 135500 681940
rect 135590 681700 135830 681940
rect 135920 681700 136160 681940
rect 136250 681700 136490 681940
rect 136600 681700 136840 681940
rect 136930 681700 137170 681940
rect 137260 681700 137500 681940
rect 137590 681700 137830 681940
rect 137940 681700 138180 681940
rect 138270 681700 138510 681940
rect 138600 681700 138840 681940
rect 138930 681700 139170 681940
rect 139280 681700 139520 681940
rect 139610 681700 139850 681940
rect 139940 681700 140180 681940
rect 140270 681700 140510 681940
rect 140620 681700 140860 681940
rect 140950 681700 141190 681940
rect 141280 681700 141520 681940
rect 141610 681700 141850 681940
rect 141960 681700 142200 681940
rect 142290 681700 142530 681940
rect 142620 681700 142860 681940
rect 142950 681700 143190 681940
rect 143300 681700 143540 681940
rect 143630 681700 143870 681940
rect 143960 681700 144200 681940
rect 144290 681700 144530 681940
rect 133570 681370 133810 681610
rect 133920 681370 134160 681610
rect 134250 681370 134490 681610
rect 134580 681370 134820 681610
rect 134910 681370 135150 681610
rect 135260 681370 135500 681610
rect 135590 681370 135830 681610
rect 135920 681370 136160 681610
rect 136250 681370 136490 681610
rect 136600 681370 136840 681610
rect 136930 681370 137170 681610
rect 137260 681370 137500 681610
rect 137590 681370 137830 681610
rect 137940 681370 138180 681610
rect 138270 681370 138510 681610
rect 138600 681370 138840 681610
rect 138930 681370 139170 681610
rect 139280 681370 139520 681610
rect 139610 681370 139850 681610
rect 139940 681370 140180 681610
rect 140270 681370 140510 681610
rect 140620 681370 140860 681610
rect 140950 681370 141190 681610
rect 141280 681370 141520 681610
rect 141610 681370 141850 681610
rect 141960 681370 142200 681610
rect 142290 681370 142530 681610
rect 142620 681370 142860 681610
rect 142950 681370 143190 681610
rect 143300 681370 143540 681610
rect 143630 681370 143870 681610
rect 143960 681370 144200 681610
rect 144290 681370 144530 681610
rect 133570 681040 133810 681280
rect 133920 681040 134160 681280
rect 134250 681040 134490 681280
rect 134580 681040 134820 681280
rect 134910 681040 135150 681280
rect 135260 681040 135500 681280
rect 135590 681040 135830 681280
rect 135920 681040 136160 681280
rect 136250 681040 136490 681280
rect 136600 681040 136840 681280
rect 136930 681040 137170 681280
rect 137260 681040 137500 681280
rect 137590 681040 137830 681280
rect 137940 681040 138180 681280
rect 138270 681040 138510 681280
rect 138600 681040 138840 681280
rect 138930 681040 139170 681280
rect 139280 681040 139520 681280
rect 139610 681040 139850 681280
rect 139940 681040 140180 681280
rect 140270 681040 140510 681280
rect 140620 681040 140860 681280
rect 140950 681040 141190 681280
rect 141280 681040 141520 681280
rect 141610 681040 141850 681280
rect 141960 681040 142200 681280
rect 142290 681040 142530 681280
rect 142620 681040 142860 681280
rect 142950 681040 143190 681280
rect 143300 681040 143540 681280
rect 143630 681040 143870 681280
rect 143960 681040 144200 681280
rect 144290 681040 144530 681280
rect 133570 680710 133810 680950
rect 133920 680710 134160 680950
rect 134250 680710 134490 680950
rect 134580 680710 134820 680950
rect 134910 680710 135150 680950
rect 135260 680710 135500 680950
rect 135590 680710 135830 680950
rect 135920 680710 136160 680950
rect 136250 680710 136490 680950
rect 136600 680710 136840 680950
rect 136930 680710 137170 680950
rect 137260 680710 137500 680950
rect 137590 680710 137830 680950
rect 137940 680710 138180 680950
rect 138270 680710 138510 680950
rect 138600 680710 138840 680950
rect 138930 680710 139170 680950
rect 139280 680710 139520 680950
rect 139610 680710 139850 680950
rect 139940 680710 140180 680950
rect 140270 680710 140510 680950
rect 140620 680710 140860 680950
rect 140950 680710 141190 680950
rect 141280 680710 141520 680950
rect 141610 680710 141850 680950
rect 141960 680710 142200 680950
rect 142290 680710 142530 680950
rect 142620 680710 142860 680950
rect 142950 680710 143190 680950
rect 143300 680710 143540 680950
rect 143630 680710 143870 680950
rect 143960 680710 144200 680950
rect 144290 680710 144530 680950
rect 133570 680360 133810 680600
rect 133920 680360 134160 680600
rect 134250 680360 134490 680600
rect 134580 680360 134820 680600
rect 134910 680360 135150 680600
rect 135260 680360 135500 680600
rect 135590 680360 135830 680600
rect 135920 680360 136160 680600
rect 136250 680360 136490 680600
rect 136600 680360 136840 680600
rect 136930 680360 137170 680600
rect 137260 680360 137500 680600
rect 137590 680360 137830 680600
rect 137940 680360 138180 680600
rect 138270 680360 138510 680600
rect 138600 680360 138840 680600
rect 138930 680360 139170 680600
rect 139280 680360 139520 680600
rect 139610 680360 139850 680600
rect 139940 680360 140180 680600
rect 140270 680360 140510 680600
rect 140620 680360 140860 680600
rect 140950 680360 141190 680600
rect 141280 680360 141520 680600
rect 141610 680360 141850 680600
rect 141960 680360 142200 680600
rect 142290 680360 142530 680600
rect 142620 680360 142860 680600
rect 142950 680360 143190 680600
rect 143300 680360 143540 680600
rect 143630 680360 143870 680600
rect 143960 680360 144200 680600
rect 144290 680360 144530 680600
rect 133570 680030 133810 680270
rect 133920 680030 134160 680270
rect 134250 680030 134490 680270
rect 134580 680030 134820 680270
rect 134910 680030 135150 680270
rect 135260 680030 135500 680270
rect 135590 680030 135830 680270
rect 135920 680030 136160 680270
rect 136250 680030 136490 680270
rect 136600 680030 136840 680270
rect 136930 680030 137170 680270
rect 137260 680030 137500 680270
rect 137590 680030 137830 680270
rect 137940 680030 138180 680270
rect 138270 680030 138510 680270
rect 138600 680030 138840 680270
rect 138930 680030 139170 680270
rect 139280 680030 139520 680270
rect 139610 680030 139850 680270
rect 139940 680030 140180 680270
rect 140270 680030 140510 680270
rect 140620 680030 140860 680270
rect 140950 680030 141190 680270
rect 141280 680030 141520 680270
rect 141610 680030 141850 680270
rect 141960 680030 142200 680270
rect 142290 680030 142530 680270
rect 142620 680030 142860 680270
rect 142950 680030 143190 680270
rect 143300 680030 143540 680270
rect 143630 680030 143870 680270
rect 143960 680030 144200 680270
rect 144290 680030 144530 680270
rect 133570 679700 133810 679940
rect 133920 679700 134160 679940
rect 134250 679700 134490 679940
rect 134580 679700 134820 679940
rect 134910 679700 135150 679940
rect 135260 679700 135500 679940
rect 135590 679700 135830 679940
rect 135920 679700 136160 679940
rect 136250 679700 136490 679940
rect 136600 679700 136840 679940
rect 136930 679700 137170 679940
rect 137260 679700 137500 679940
rect 137590 679700 137830 679940
rect 137940 679700 138180 679940
rect 138270 679700 138510 679940
rect 138600 679700 138840 679940
rect 138930 679700 139170 679940
rect 139280 679700 139520 679940
rect 139610 679700 139850 679940
rect 139940 679700 140180 679940
rect 140270 679700 140510 679940
rect 140620 679700 140860 679940
rect 140950 679700 141190 679940
rect 141280 679700 141520 679940
rect 141610 679700 141850 679940
rect 141960 679700 142200 679940
rect 142290 679700 142530 679940
rect 142620 679700 142860 679940
rect 142950 679700 143190 679940
rect 143300 679700 143540 679940
rect 143630 679700 143870 679940
rect 143960 679700 144200 679940
rect 144290 679700 144530 679940
rect 133570 679370 133810 679610
rect 133920 679370 134160 679610
rect 134250 679370 134490 679610
rect 134580 679370 134820 679610
rect 134910 679370 135150 679610
rect 135260 679370 135500 679610
rect 135590 679370 135830 679610
rect 135920 679370 136160 679610
rect 136250 679370 136490 679610
rect 136600 679370 136840 679610
rect 136930 679370 137170 679610
rect 137260 679370 137500 679610
rect 137590 679370 137830 679610
rect 137940 679370 138180 679610
rect 138270 679370 138510 679610
rect 138600 679370 138840 679610
rect 138930 679370 139170 679610
rect 139280 679370 139520 679610
rect 139610 679370 139850 679610
rect 139940 679370 140180 679610
rect 140270 679370 140510 679610
rect 140620 679370 140860 679610
rect 140950 679370 141190 679610
rect 141280 679370 141520 679610
rect 141610 679370 141850 679610
rect 141960 679370 142200 679610
rect 142290 679370 142530 679610
rect 142620 679370 142860 679610
rect 142950 679370 143190 679610
rect 143300 679370 143540 679610
rect 143630 679370 143870 679610
rect 143960 679370 144200 679610
rect 144290 679370 144530 679610
rect 133570 679020 133810 679260
rect 133920 679020 134160 679260
rect 134250 679020 134490 679260
rect 134580 679020 134820 679260
rect 134910 679020 135150 679260
rect 135260 679020 135500 679260
rect 135590 679020 135830 679260
rect 135920 679020 136160 679260
rect 136250 679020 136490 679260
rect 136600 679020 136840 679260
rect 136930 679020 137170 679260
rect 137260 679020 137500 679260
rect 137590 679020 137830 679260
rect 137940 679020 138180 679260
rect 138270 679020 138510 679260
rect 138600 679020 138840 679260
rect 138930 679020 139170 679260
rect 139280 679020 139520 679260
rect 139610 679020 139850 679260
rect 139940 679020 140180 679260
rect 140270 679020 140510 679260
rect 140620 679020 140860 679260
rect 140950 679020 141190 679260
rect 141280 679020 141520 679260
rect 141610 679020 141850 679260
rect 141960 679020 142200 679260
rect 142290 679020 142530 679260
rect 142620 679020 142860 679260
rect 142950 679020 143190 679260
rect 143300 679020 143540 679260
rect 143630 679020 143870 679260
rect 143960 679020 144200 679260
rect 144290 679020 144530 679260
rect 133570 678690 133810 678930
rect 133920 678690 134160 678930
rect 134250 678690 134490 678930
rect 134580 678690 134820 678930
rect 134910 678690 135150 678930
rect 135260 678690 135500 678930
rect 135590 678690 135830 678930
rect 135920 678690 136160 678930
rect 136250 678690 136490 678930
rect 136600 678690 136840 678930
rect 136930 678690 137170 678930
rect 137260 678690 137500 678930
rect 137590 678690 137830 678930
rect 137940 678690 138180 678930
rect 138270 678690 138510 678930
rect 138600 678690 138840 678930
rect 138930 678690 139170 678930
rect 139280 678690 139520 678930
rect 139610 678690 139850 678930
rect 139940 678690 140180 678930
rect 140270 678690 140510 678930
rect 140620 678690 140860 678930
rect 140950 678690 141190 678930
rect 141280 678690 141520 678930
rect 141610 678690 141850 678930
rect 141960 678690 142200 678930
rect 142290 678690 142530 678930
rect 142620 678690 142860 678930
rect 142950 678690 143190 678930
rect 143300 678690 143540 678930
rect 143630 678690 143870 678930
rect 143960 678690 144200 678930
rect 144290 678690 144530 678930
rect 133570 678360 133810 678600
rect 133920 678360 134160 678600
rect 134250 678360 134490 678600
rect 134580 678360 134820 678600
rect 134910 678360 135150 678600
rect 135260 678360 135500 678600
rect 135590 678360 135830 678600
rect 135920 678360 136160 678600
rect 136250 678360 136490 678600
rect 136600 678360 136840 678600
rect 136930 678360 137170 678600
rect 137260 678360 137500 678600
rect 137590 678360 137830 678600
rect 137940 678360 138180 678600
rect 138270 678360 138510 678600
rect 138600 678360 138840 678600
rect 138930 678360 139170 678600
rect 139280 678360 139520 678600
rect 139610 678360 139850 678600
rect 139940 678360 140180 678600
rect 140270 678360 140510 678600
rect 140620 678360 140860 678600
rect 140950 678360 141190 678600
rect 141280 678360 141520 678600
rect 141610 678360 141850 678600
rect 141960 678360 142200 678600
rect 142290 678360 142530 678600
rect 142620 678360 142860 678600
rect 142950 678360 143190 678600
rect 143300 678360 143540 678600
rect 143630 678360 143870 678600
rect 143960 678360 144200 678600
rect 144290 678360 144530 678600
rect 133570 678030 133810 678270
rect 133920 678030 134160 678270
rect 134250 678030 134490 678270
rect 134580 678030 134820 678270
rect 134910 678030 135150 678270
rect 135260 678030 135500 678270
rect 135590 678030 135830 678270
rect 135920 678030 136160 678270
rect 136250 678030 136490 678270
rect 136600 678030 136840 678270
rect 136930 678030 137170 678270
rect 137260 678030 137500 678270
rect 137590 678030 137830 678270
rect 137940 678030 138180 678270
rect 138270 678030 138510 678270
rect 138600 678030 138840 678270
rect 138930 678030 139170 678270
rect 139280 678030 139520 678270
rect 139610 678030 139850 678270
rect 139940 678030 140180 678270
rect 140270 678030 140510 678270
rect 140620 678030 140860 678270
rect 140950 678030 141190 678270
rect 141280 678030 141520 678270
rect 141610 678030 141850 678270
rect 141960 678030 142200 678270
rect 142290 678030 142530 678270
rect 142620 678030 142860 678270
rect 142950 678030 143190 678270
rect 143300 678030 143540 678270
rect 143630 678030 143870 678270
rect 143960 678030 144200 678270
rect 144290 678030 144530 678270
rect 133570 677680 133810 677920
rect 133920 677680 134160 677920
rect 134250 677680 134490 677920
rect 134580 677680 134820 677920
rect 134910 677680 135150 677920
rect 135260 677680 135500 677920
rect 135590 677680 135830 677920
rect 135920 677680 136160 677920
rect 136250 677680 136490 677920
rect 136600 677680 136840 677920
rect 136930 677680 137170 677920
rect 137260 677680 137500 677920
rect 137590 677680 137830 677920
rect 137940 677680 138180 677920
rect 138270 677680 138510 677920
rect 138600 677680 138840 677920
rect 138930 677680 139170 677920
rect 139280 677680 139520 677920
rect 139610 677680 139850 677920
rect 139940 677680 140180 677920
rect 140270 677680 140510 677920
rect 140620 677680 140860 677920
rect 140950 677680 141190 677920
rect 141280 677680 141520 677920
rect 141610 677680 141850 677920
rect 141960 677680 142200 677920
rect 142290 677680 142530 677920
rect 142620 677680 142860 677920
rect 142950 677680 143190 677920
rect 143300 677680 143540 677920
rect 143630 677680 143870 677920
rect 143960 677680 144200 677920
rect 144290 677680 144530 677920
rect 133570 677350 133810 677590
rect 133920 677350 134160 677590
rect 134250 677350 134490 677590
rect 134580 677350 134820 677590
rect 134910 677350 135150 677590
rect 135260 677350 135500 677590
rect 135590 677350 135830 677590
rect 135920 677350 136160 677590
rect 136250 677350 136490 677590
rect 136600 677350 136840 677590
rect 136930 677350 137170 677590
rect 137260 677350 137500 677590
rect 137590 677350 137830 677590
rect 137940 677350 138180 677590
rect 138270 677350 138510 677590
rect 138600 677350 138840 677590
rect 138930 677350 139170 677590
rect 139280 677350 139520 677590
rect 139610 677350 139850 677590
rect 139940 677350 140180 677590
rect 140270 677350 140510 677590
rect 140620 677350 140860 677590
rect 140950 677350 141190 677590
rect 141280 677350 141520 677590
rect 141610 677350 141850 677590
rect 141960 677350 142200 677590
rect 142290 677350 142530 677590
rect 142620 677350 142860 677590
rect 142950 677350 143190 677590
rect 143300 677350 143540 677590
rect 143630 677350 143870 677590
rect 143960 677350 144200 677590
rect 144290 677350 144530 677590
rect 133570 677020 133810 677260
rect 133920 677020 134160 677260
rect 134250 677020 134490 677260
rect 134580 677020 134820 677260
rect 134910 677020 135150 677260
rect 135260 677020 135500 677260
rect 135590 677020 135830 677260
rect 135920 677020 136160 677260
rect 136250 677020 136490 677260
rect 136600 677020 136840 677260
rect 136930 677020 137170 677260
rect 137260 677020 137500 677260
rect 137590 677020 137830 677260
rect 137940 677020 138180 677260
rect 138270 677020 138510 677260
rect 138600 677020 138840 677260
rect 138930 677020 139170 677260
rect 139280 677020 139520 677260
rect 139610 677020 139850 677260
rect 139940 677020 140180 677260
rect 140270 677020 140510 677260
rect 140620 677020 140860 677260
rect 140950 677020 141190 677260
rect 141280 677020 141520 677260
rect 141610 677020 141850 677260
rect 141960 677020 142200 677260
rect 142290 677020 142530 677260
rect 142620 677020 142860 677260
rect 142950 677020 143190 677260
rect 143300 677020 143540 677260
rect 143630 677020 143870 677260
rect 143960 677020 144200 677260
rect 144290 677020 144530 677260
rect 133570 676690 133810 676930
rect 133920 676690 134160 676930
rect 134250 676690 134490 676930
rect 134580 676690 134820 676930
rect 134910 676690 135150 676930
rect 135260 676690 135500 676930
rect 135590 676690 135830 676930
rect 135920 676690 136160 676930
rect 136250 676690 136490 676930
rect 136600 676690 136840 676930
rect 136930 676690 137170 676930
rect 137260 676690 137500 676930
rect 137590 676690 137830 676930
rect 137940 676690 138180 676930
rect 138270 676690 138510 676930
rect 138600 676690 138840 676930
rect 138930 676690 139170 676930
rect 139280 676690 139520 676930
rect 139610 676690 139850 676930
rect 139940 676690 140180 676930
rect 140270 676690 140510 676930
rect 140620 676690 140860 676930
rect 140950 676690 141190 676930
rect 141280 676690 141520 676930
rect 141610 676690 141850 676930
rect 141960 676690 142200 676930
rect 142290 676690 142530 676930
rect 142620 676690 142860 676930
rect 142950 676690 143190 676930
rect 143300 676690 143540 676930
rect 143630 676690 143870 676930
rect 143960 676690 144200 676930
rect 144290 676690 144530 676930
rect 133570 676340 133810 676580
rect 133920 676340 134160 676580
rect 134250 676340 134490 676580
rect 134580 676340 134820 676580
rect 134910 676340 135150 676580
rect 135260 676340 135500 676580
rect 135590 676340 135830 676580
rect 135920 676340 136160 676580
rect 136250 676340 136490 676580
rect 136600 676340 136840 676580
rect 136930 676340 137170 676580
rect 137260 676340 137500 676580
rect 137590 676340 137830 676580
rect 137940 676340 138180 676580
rect 138270 676340 138510 676580
rect 138600 676340 138840 676580
rect 138930 676340 139170 676580
rect 139280 676340 139520 676580
rect 139610 676340 139850 676580
rect 139940 676340 140180 676580
rect 140270 676340 140510 676580
rect 140620 676340 140860 676580
rect 140950 676340 141190 676580
rect 141280 676340 141520 676580
rect 141610 676340 141850 676580
rect 141960 676340 142200 676580
rect 142290 676340 142530 676580
rect 142620 676340 142860 676580
rect 142950 676340 143190 676580
rect 143300 676340 143540 676580
rect 143630 676340 143870 676580
rect 143960 676340 144200 676580
rect 144290 676340 144530 676580
rect 133570 676010 133810 676250
rect 133920 676010 134160 676250
rect 134250 676010 134490 676250
rect 134580 676010 134820 676250
rect 134910 676010 135150 676250
rect 135260 676010 135500 676250
rect 135590 676010 135830 676250
rect 135920 676010 136160 676250
rect 136250 676010 136490 676250
rect 136600 676010 136840 676250
rect 136930 676010 137170 676250
rect 137260 676010 137500 676250
rect 137590 676010 137830 676250
rect 137940 676010 138180 676250
rect 138270 676010 138510 676250
rect 138600 676010 138840 676250
rect 138930 676010 139170 676250
rect 139280 676010 139520 676250
rect 139610 676010 139850 676250
rect 139940 676010 140180 676250
rect 140270 676010 140510 676250
rect 140620 676010 140860 676250
rect 140950 676010 141190 676250
rect 141280 676010 141520 676250
rect 141610 676010 141850 676250
rect 141960 676010 142200 676250
rect 142290 676010 142530 676250
rect 142620 676010 142860 676250
rect 142950 676010 143190 676250
rect 143300 676010 143540 676250
rect 143630 676010 143870 676250
rect 143960 676010 144200 676250
rect 144290 676010 144530 676250
rect 133570 675680 133810 675920
rect 133920 675680 134160 675920
rect 134250 675680 134490 675920
rect 134580 675680 134820 675920
rect 134910 675680 135150 675920
rect 135260 675680 135500 675920
rect 135590 675680 135830 675920
rect 135920 675680 136160 675920
rect 136250 675680 136490 675920
rect 136600 675680 136840 675920
rect 136930 675680 137170 675920
rect 137260 675680 137500 675920
rect 137590 675680 137830 675920
rect 137940 675680 138180 675920
rect 138270 675680 138510 675920
rect 138600 675680 138840 675920
rect 138930 675680 139170 675920
rect 139280 675680 139520 675920
rect 139610 675680 139850 675920
rect 139940 675680 140180 675920
rect 140270 675680 140510 675920
rect 140620 675680 140860 675920
rect 140950 675680 141190 675920
rect 141280 675680 141520 675920
rect 141610 675680 141850 675920
rect 141960 675680 142200 675920
rect 142290 675680 142530 675920
rect 142620 675680 142860 675920
rect 142950 675680 143190 675920
rect 143300 675680 143540 675920
rect 143630 675680 143870 675920
rect 143960 675680 144200 675920
rect 144290 675680 144530 675920
rect 133570 675350 133810 675590
rect 133920 675350 134160 675590
rect 134250 675350 134490 675590
rect 134580 675350 134820 675590
rect 134910 675350 135150 675590
rect 135260 675350 135500 675590
rect 135590 675350 135830 675590
rect 135920 675350 136160 675590
rect 136250 675350 136490 675590
rect 136600 675350 136840 675590
rect 136930 675350 137170 675590
rect 137260 675350 137500 675590
rect 137590 675350 137830 675590
rect 137940 675350 138180 675590
rect 138270 675350 138510 675590
rect 138600 675350 138840 675590
rect 138930 675350 139170 675590
rect 139280 675350 139520 675590
rect 139610 675350 139850 675590
rect 139940 675350 140180 675590
rect 140270 675350 140510 675590
rect 140620 675350 140860 675590
rect 140950 675350 141190 675590
rect 141280 675350 141520 675590
rect 141610 675350 141850 675590
rect 141960 675350 142200 675590
rect 142290 675350 142530 675590
rect 142620 675350 142860 675590
rect 142950 675350 143190 675590
rect 143300 675350 143540 675590
rect 143630 675350 143870 675590
rect 143960 675350 144200 675590
rect 144290 675350 144530 675590
rect 133570 675000 133810 675240
rect 133920 675000 134160 675240
rect 134250 675000 134490 675240
rect 134580 675000 134820 675240
rect 134910 675000 135150 675240
rect 135260 675000 135500 675240
rect 135590 675000 135830 675240
rect 135920 675000 136160 675240
rect 136250 675000 136490 675240
rect 136600 675000 136840 675240
rect 136930 675000 137170 675240
rect 137260 675000 137500 675240
rect 137590 675000 137830 675240
rect 137940 675000 138180 675240
rect 138270 675000 138510 675240
rect 138600 675000 138840 675240
rect 138930 675000 139170 675240
rect 139280 675000 139520 675240
rect 139610 675000 139850 675240
rect 139940 675000 140180 675240
rect 140270 675000 140510 675240
rect 140620 675000 140860 675240
rect 140950 675000 141190 675240
rect 141280 675000 141520 675240
rect 141610 675000 141850 675240
rect 141960 675000 142200 675240
rect 142290 675000 142530 675240
rect 142620 675000 142860 675240
rect 142950 675000 143190 675240
rect 143300 675000 143540 675240
rect 143630 675000 143870 675240
rect 143960 675000 144200 675240
rect 144290 675000 144530 675240
rect 133570 674670 133810 674910
rect 133920 674670 134160 674910
rect 134250 674670 134490 674910
rect 134580 674670 134820 674910
rect 134910 674670 135150 674910
rect 135260 674670 135500 674910
rect 135590 674670 135830 674910
rect 135920 674670 136160 674910
rect 136250 674670 136490 674910
rect 136600 674670 136840 674910
rect 136930 674670 137170 674910
rect 137260 674670 137500 674910
rect 137590 674670 137830 674910
rect 137940 674670 138180 674910
rect 138270 674670 138510 674910
rect 138600 674670 138840 674910
rect 138930 674670 139170 674910
rect 139280 674670 139520 674910
rect 139610 674670 139850 674910
rect 139940 674670 140180 674910
rect 140270 674670 140510 674910
rect 140620 674670 140860 674910
rect 140950 674670 141190 674910
rect 141280 674670 141520 674910
rect 141610 674670 141850 674910
rect 141960 674670 142200 674910
rect 142290 674670 142530 674910
rect 142620 674670 142860 674910
rect 142950 674670 143190 674910
rect 143300 674670 143540 674910
rect 143630 674670 143870 674910
rect 143960 674670 144200 674910
rect 144290 674670 144530 674910
rect 133570 674340 133810 674580
rect 133920 674340 134160 674580
rect 134250 674340 134490 674580
rect 134580 674340 134820 674580
rect 134910 674340 135150 674580
rect 135260 674340 135500 674580
rect 135590 674340 135830 674580
rect 135920 674340 136160 674580
rect 136250 674340 136490 674580
rect 136600 674340 136840 674580
rect 136930 674340 137170 674580
rect 137260 674340 137500 674580
rect 137590 674340 137830 674580
rect 137940 674340 138180 674580
rect 138270 674340 138510 674580
rect 138600 674340 138840 674580
rect 138930 674340 139170 674580
rect 139280 674340 139520 674580
rect 139610 674340 139850 674580
rect 139940 674340 140180 674580
rect 140270 674340 140510 674580
rect 140620 674340 140860 674580
rect 140950 674340 141190 674580
rect 141280 674340 141520 674580
rect 141610 674340 141850 674580
rect 141960 674340 142200 674580
rect 142290 674340 142530 674580
rect 142620 674340 142860 674580
rect 142950 674340 143190 674580
rect 143300 674340 143540 674580
rect 143630 674340 143870 674580
rect 143960 674340 144200 674580
rect 144290 674340 144530 674580
rect 133570 674010 133810 674250
rect 133920 674010 134160 674250
rect 134250 674010 134490 674250
rect 134580 674010 134820 674250
rect 134910 674010 135150 674250
rect 135260 674010 135500 674250
rect 135590 674010 135830 674250
rect 135920 674010 136160 674250
rect 136250 674010 136490 674250
rect 136600 674010 136840 674250
rect 136930 674010 137170 674250
rect 137260 674010 137500 674250
rect 137590 674010 137830 674250
rect 137940 674010 138180 674250
rect 138270 674010 138510 674250
rect 138600 674010 138840 674250
rect 138930 674010 139170 674250
rect 139280 674010 139520 674250
rect 139610 674010 139850 674250
rect 139940 674010 140180 674250
rect 140270 674010 140510 674250
rect 140620 674010 140860 674250
rect 140950 674010 141190 674250
rect 141280 674010 141520 674250
rect 141610 674010 141850 674250
rect 141960 674010 142200 674250
rect 142290 674010 142530 674250
rect 142620 674010 142860 674250
rect 142950 674010 143190 674250
rect 143300 674010 143540 674250
rect 143630 674010 143870 674250
rect 143960 674010 144200 674250
rect 144290 674010 144530 674250
rect 133570 673660 133810 673900
rect 133920 673660 134160 673900
rect 134250 673660 134490 673900
rect 134580 673660 134820 673900
rect 134910 673660 135150 673900
rect 135260 673660 135500 673900
rect 135590 673660 135830 673900
rect 135920 673660 136160 673900
rect 136250 673660 136490 673900
rect 136600 673660 136840 673900
rect 136930 673660 137170 673900
rect 137260 673660 137500 673900
rect 137590 673660 137830 673900
rect 137940 673660 138180 673900
rect 138270 673660 138510 673900
rect 138600 673660 138840 673900
rect 138930 673660 139170 673900
rect 139280 673660 139520 673900
rect 139610 673660 139850 673900
rect 139940 673660 140180 673900
rect 140270 673660 140510 673900
rect 140620 673660 140860 673900
rect 140950 673660 141190 673900
rect 141280 673660 141520 673900
rect 141610 673660 141850 673900
rect 141960 673660 142200 673900
rect 142290 673660 142530 673900
rect 142620 673660 142860 673900
rect 142950 673660 143190 673900
rect 143300 673660 143540 673900
rect 143630 673660 143870 673900
rect 143960 673660 144200 673900
rect 144290 673660 144530 673900
rect 133570 673330 133810 673570
rect 133920 673330 134160 673570
rect 134250 673330 134490 673570
rect 134580 673330 134820 673570
rect 134910 673330 135150 673570
rect 135260 673330 135500 673570
rect 135590 673330 135830 673570
rect 135920 673330 136160 673570
rect 136250 673330 136490 673570
rect 136600 673330 136840 673570
rect 136930 673330 137170 673570
rect 137260 673330 137500 673570
rect 137590 673330 137830 673570
rect 137940 673330 138180 673570
rect 138270 673330 138510 673570
rect 138600 673330 138840 673570
rect 138930 673330 139170 673570
rect 139280 673330 139520 673570
rect 139610 673330 139850 673570
rect 139940 673330 140180 673570
rect 140270 673330 140510 673570
rect 140620 673330 140860 673570
rect 140950 673330 141190 673570
rect 141280 673330 141520 673570
rect 141610 673330 141850 673570
rect 141960 673330 142200 673570
rect 142290 673330 142530 673570
rect 142620 673330 142860 673570
rect 142950 673330 143190 673570
rect 143300 673330 143540 673570
rect 143630 673330 143870 673570
rect 143960 673330 144200 673570
rect 144290 673330 144530 673570
rect 133570 673000 133810 673240
rect 133920 673000 134160 673240
rect 134250 673000 134490 673240
rect 134580 673000 134820 673240
rect 134910 673000 135150 673240
rect 135260 673000 135500 673240
rect 135590 673000 135830 673240
rect 135920 673000 136160 673240
rect 136250 673000 136490 673240
rect 136600 673000 136840 673240
rect 136930 673000 137170 673240
rect 137260 673000 137500 673240
rect 137590 673000 137830 673240
rect 137940 673000 138180 673240
rect 138270 673000 138510 673240
rect 138600 673000 138840 673240
rect 138930 673000 139170 673240
rect 139280 673000 139520 673240
rect 139610 673000 139850 673240
rect 139940 673000 140180 673240
rect 140270 673000 140510 673240
rect 140620 673000 140860 673240
rect 140950 673000 141190 673240
rect 141280 673000 141520 673240
rect 141610 673000 141850 673240
rect 141960 673000 142200 673240
rect 142290 673000 142530 673240
rect 142620 673000 142860 673240
rect 142950 673000 143190 673240
rect 143300 673000 143540 673240
rect 143630 673000 143870 673240
rect 143960 673000 144200 673240
rect 144290 673000 144530 673240
rect 133570 672670 133810 672910
rect 133920 672670 134160 672910
rect 134250 672670 134490 672910
rect 134580 672670 134820 672910
rect 134910 672670 135150 672910
rect 135260 672670 135500 672910
rect 135590 672670 135830 672910
rect 135920 672670 136160 672910
rect 136250 672670 136490 672910
rect 136600 672670 136840 672910
rect 136930 672670 137170 672910
rect 137260 672670 137500 672910
rect 137590 672670 137830 672910
rect 137940 672670 138180 672910
rect 138270 672670 138510 672910
rect 138600 672670 138840 672910
rect 138930 672670 139170 672910
rect 139280 672670 139520 672910
rect 139610 672670 139850 672910
rect 139940 672670 140180 672910
rect 140270 672670 140510 672910
rect 140620 672670 140860 672910
rect 140950 672670 141190 672910
rect 141280 672670 141520 672910
rect 141610 672670 141850 672910
rect 141960 672670 142200 672910
rect 142290 672670 142530 672910
rect 142620 672670 142860 672910
rect 142950 672670 143190 672910
rect 143300 672670 143540 672910
rect 143630 672670 143870 672910
rect 143960 672670 144200 672910
rect 144290 672670 144530 672910
rect 133570 672320 133810 672560
rect 133920 672320 134160 672560
rect 134250 672320 134490 672560
rect 134580 672320 134820 672560
rect 134910 672320 135150 672560
rect 135260 672320 135500 672560
rect 135590 672320 135830 672560
rect 135920 672320 136160 672560
rect 136250 672320 136490 672560
rect 136600 672320 136840 672560
rect 136930 672320 137170 672560
rect 137260 672320 137500 672560
rect 137590 672320 137830 672560
rect 137940 672320 138180 672560
rect 138270 672320 138510 672560
rect 138600 672320 138840 672560
rect 138930 672320 139170 672560
rect 139280 672320 139520 672560
rect 139610 672320 139850 672560
rect 139940 672320 140180 672560
rect 140270 672320 140510 672560
rect 140620 672320 140860 672560
rect 140950 672320 141190 672560
rect 141280 672320 141520 672560
rect 141610 672320 141850 672560
rect 141960 672320 142200 672560
rect 142290 672320 142530 672560
rect 142620 672320 142860 672560
rect 142950 672320 143190 672560
rect 143300 672320 143540 672560
rect 143630 672320 143870 672560
rect 143960 672320 144200 672560
rect 144290 672320 144530 672560
rect 144950 683040 145190 683280
rect 145300 683040 145540 683280
rect 145630 683040 145870 683280
rect 145960 683040 146200 683280
rect 146290 683040 146530 683280
rect 146640 683040 146880 683280
rect 146970 683040 147210 683280
rect 147300 683040 147540 683280
rect 147630 683040 147870 683280
rect 147980 683040 148220 683280
rect 148310 683040 148550 683280
rect 148640 683040 148880 683280
rect 148970 683040 149210 683280
rect 149320 683040 149560 683280
rect 149650 683040 149890 683280
rect 149980 683040 150220 683280
rect 150310 683040 150550 683280
rect 150660 683040 150900 683280
rect 150990 683040 151230 683280
rect 151320 683040 151560 683280
rect 151650 683040 151890 683280
rect 152000 683040 152240 683280
rect 152330 683040 152570 683280
rect 152660 683040 152900 683280
rect 152990 683040 153230 683280
rect 153340 683040 153580 683280
rect 153670 683040 153910 683280
rect 154000 683040 154240 683280
rect 154330 683040 154570 683280
rect 154680 683040 154920 683280
rect 155010 683040 155250 683280
rect 155340 683040 155580 683280
rect 155670 683040 155910 683280
rect 144950 682710 145190 682950
rect 145300 682710 145540 682950
rect 145630 682710 145870 682950
rect 145960 682710 146200 682950
rect 146290 682710 146530 682950
rect 146640 682710 146880 682950
rect 146970 682710 147210 682950
rect 147300 682710 147540 682950
rect 147630 682710 147870 682950
rect 147980 682710 148220 682950
rect 148310 682710 148550 682950
rect 148640 682710 148880 682950
rect 148970 682710 149210 682950
rect 149320 682710 149560 682950
rect 149650 682710 149890 682950
rect 149980 682710 150220 682950
rect 150310 682710 150550 682950
rect 150660 682710 150900 682950
rect 150990 682710 151230 682950
rect 151320 682710 151560 682950
rect 151650 682710 151890 682950
rect 152000 682710 152240 682950
rect 152330 682710 152570 682950
rect 152660 682710 152900 682950
rect 152990 682710 153230 682950
rect 153340 682710 153580 682950
rect 153670 682710 153910 682950
rect 154000 682710 154240 682950
rect 154330 682710 154570 682950
rect 154680 682710 154920 682950
rect 155010 682710 155250 682950
rect 155340 682710 155580 682950
rect 155670 682710 155910 682950
rect 144950 682380 145190 682620
rect 145300 682380 145540 682620
rect 145630 682380 145870 682620
rect 145960 682380 146200 682620
rect 146290 682380 146530 682620
rect 146640 682380 146880 682620
rect 146970 682380 147210 682620
rect 147300 682380 147540 682620
rect 147630 682380 147870 682620
rect 147980 682380 148220 682620
rect 148310 682380 148550 682620
rect 148640 682380 148880 682620
rect 148970 682380 149210 682620
rect 149320 682380 149560 682620
rect 149650 682380 149890 682620
rect 149980 682380 150220 682620
rect 150310 682380 150550 682620
rect 150660 682380 150900 682620
rect 150990 682380 151230 682620
rect 151320 682380 151560 682620
rect 151650 682380 151890 682620
rect 152000 682380 152240 682620
rect 152330 682380 152570 682620
rect 152660 682380 152900 682620
rect 152990 682380 153230 682620
rect 153340 682380 153580 682620
rect 153670 682380 153910 682620
rect 154000 682380 154240 682620
rect 154330 682380 154570 682620
rect 154680 682380 154920 682620
rect 155010 682380 155250 682620
rect 155340 682380 155580 682620
rect 155670 682380 155910 682620
rect 144950 682050 145190 682290
rect 145300 682050 145540 682290
rect 145630 682050 145870 682290
rect 145960 682050 146200 682290
rect 146290 682050 146530 682290
rect 146640 682050 146880 682290
rect 146970 682050 147210 682290
rect 147300 682050 147540 682290
rect 147630 682050 147870 682290
rect 147980 682050 148220 682290
rect 148310 682050 148550 682290
rect 148640 682050 148880 682290
rect 148970 682050 149210 682290
rect 149320 682050 149560 682290
rect 149650 682050 149890 682290
rect 149980 682050 150220 682290
rect 150310 682050 150550 682290
rect 150660 682050 150900 682290
rect 150990 682050 151230 682290
rect 151320 682050 151560 682290
rect 151650 682050 151890 682290
rect 152000 682050 152240 682290
rect 152330 682050 152570 682290
rect 152660 682050 152900 682290
rect 152990 682050 153230 682290
rect 153340 682050 153580 682290
rect 153670 682050 153910 682290
rect 154000 682050 154240 682290
rect 154330 682050 154570 682290
rect 154680 682050 154920 682290
rect 155010 682050 155250 682290
rect 155340 682050 155580 682290
rect 155670 682050 155910 682290
rect 144950 681700 145190 681940
rect 145300 681700 145540 681940
rect 145630 681700 145870 681940
rect 145960 681700 146200 681940
rect 146290 681700 146530 681940
rect 146640 681700 146880 681940
rect 146970 681700 147210 681940
rect 147300 681700 147540 681940
rect 147630 681700 147870 681940
rect 147980 681700 148220 681940
rect 148310 681700 148550 681940
rect 148640 681700 148880 681940
rect 148970 681700 149210 681940
rect 149320 681700 149560 681940
rect 149650 681700 149890 681940
rect 149980 681700 150220 681940
rect 150310 681700 150550 681940
rect 150660 681700 150900 681940
rect 150990 681700 151230 681940
rect 151320 681700 151560 681940
rect 151650 681700 151890 681940
rect 152000 681700 152240 681940
rect 152330 681700 152570 681940
rect 152660 681700 152900 681940
rect 152990 681700 153230 681940
rect 153340 681700 153580 681940
rect 153670 681700 153910 681940
rect 154000 681700 154240 681940
rect 154330 681700 154570 681940
rect 154680 681700 154920 681940
rect 155010 681700 155250 681940
rect 155340 681700 155580 681940
rect 155670 681700 155910 681940
rect 144950 681370 145190 681610
rect 145300 681370 145540 681610
rect 145630 681370 145870 681610
rect 145960 681370 146200 681610
rect 146290 681370 146530 681610
rect 146640 681370 146880 681610
rect 146970 681370 147210 681610
rect 147300 681370 147540 681610
rect 147630 681370 147870 681610
rect 147980 681370 148220 681610
rect 148310 681370 148550 681610
rect 148640 681370 148880 681610
rect 148970 681370 149210 681610
rect 149320 681370 149560 681610
rect 149650 681370 149890 681610
rect 149980 681370 150220 681610
rect 150310 681370 150550 681610
rect 150660 681370 150900 681610
rect 150990 681370 151230 681610
rect 151320 681370 151560 681610
rect 151650 681370 151890 681610
rect 152000 681370 152240 681610
rect 152330 681370 152570 681610
rect 152660 681370 152900 681610
rect 152990 681370 153230 681610
rect 153340 681370 153580 681610
rect 153670 681370 153910 681610
rect 154000 681370 154240 681610
rect 154330 681370 154570 681610
rect 154680 681370 154920 681610
rect 155010 681370 155250 681610
rect 155340 681370 155580 681610
rect 155670 681370 155910 681610
rect 144950 681040 145190 681280
rect 145300 681040 145540 681280
rect 145630 681040 145870 681280
rect 145960 681040 146200 681280
rect 146290 681040 146530 681280
rect 146640 681040 146880 681280
rect 146970 681040 147210 681280
rect 147300 681040 147540 681280
rect 147630 681040 147870 681280
rect 147980 681040 148220 681280
rect 148310 681040 148550 681280
rect 148640 681040 148880 681280
rect 148970 681040 149210 681280
rect 149320 681040 149560 681280
rect 149650 681040 149890 681280
rect 149980 681040 150220 681280
rect 150310 681040 150550 681280
rect 150660 681040 150900 681280
rect 150990 681040 151230 681280
rect 151320 681040 151560 681280
rect 151650 681040 151890 681280
rect 152000 681040 152240 681280
rect 152330 681040 152570 681280
rect 152660 681040 152900 681280
rect 152990 681040 153230 681280
rect 153340 681040 153580 681280
rect 153670 681040 153910 681280
rect 154000 681040 154240 681280
rect 154330 681040 154570 681280
rect 154680 681040 154920 681280
rect 155010 681040 155250 681280
rect 155340 681040 155580 681280
rect 155670 681040 155910 681280
rect 144950 680710 145190 680950
rect 145300 680710 145540 680950
rect 145630 680710 145870 680950
rect 145960 680710 146200 680950
rect 146290 680710 146530 680950
rect 146640 680710 146880 680950
rect 146970 680710 147210 680950
rect 147300 680710 147540 680950
rect 147630 680710 147870 680950
rect 147980 680710 148220 680950
rect 148310 680710 148550 680950
rect 148640 680710 148880 680950
rect 148970 680710 149210 680950
rect 149320 680710 149560 680950
rect 149650 680710 149890 680950
rect 149980 680710 150220 680950
rect 150310 680710 150550 680950
rect 150660 680710 150900 680950
rect 150990 680710 151230 680950
rect 151320 680710 151560 680950
rect 151650 680710 151890 680950
rect 152000 680710 152240 680950
rect 152330 680710 152570 680950
rect 152660 680710 152900 680950
rect 152990 680710 153230 680950
rect 153340 680710 153580 680950
rect 153670 680710 153910 680950
rect 154000 680710 154240 680950
rect 154330 680710 154570 680950
rect 154680 680710 154920 680950
rect 155010 680710 155250 680950
rect 155340 680710 155580 680950
rect 155670 680710 155910 680950
rect 144950 680360 145190 680600
rect 145300 680360 145540 680600
rect 145630 680360 145870 680600
rect 145960 680360 146200 680600
rect 146290 680360 146530 680600
rect 146640 680360 146880 680600
rect 146970 680360 147210 680600
rect 147300 680360 147540 680600
rect 147630 680360 147870 680600
rect 147980 680360 148220 680600
rect 148310 680360 148550 680600
rect 148640 680360 148880 680600
rect 148970 680360 149210 680600
rect 149320 680360 149560 680600
rect 149650 680360 149890 680600
rect 149980 680360 150220 680600
rect 150310 680360 150550 680600
rect 150660 680360 150900 680600
rect 150990 680360 151230 680600
rect 151320 680360 151560 680600
rect 151650 680360 151890 680600
rect 152000 680360 152240 680600
rect 152330 680360 152570 680600
rect 152660 680360 152900 680600
rect 152990 680360 153230 680600
rect 153340 680360 153580 680600
rect 153670 680360 153910 680600
rect 154000 680360 154240 680600
rect 154330 680360 154570 680600
rect 154680 680360 154920 680600
rect 155010 680360 155250 680600
rect 155340 680360 155580 680600
rect 155670 680360 155910 680600
rect 144950 680030 145190 680270
rect 145300 680030 145540 680270
rect 145630 680030 145870 680270
rect 145960 680030 146200 680270
rect 146290 680030 146530 680270
rect 146640 680030 146880 680270
rect 146970 680030 147210 680270
rect 147300 680030 147540 680270
rect 147630 680030 147870 680270
rect 147980 680030 148220 680270
rect 148310 680030 148550 680270
rect 148640 680030 148880 680270
rect 148970 680030 149210 680270
rect 149320 680030 149560 680270
rect 149650 680030 149890 680270
rect 149980 680030 150220 680270
rect 150310 680030 150550 680270
rect 150660 680030 150900 680270
rect 150990 680030 151230 680270
rect 151320 680030 151560 680270
rect 151650 680030 151890 680270
rect 152000 680030 152240 680270
rect 152330 680030 152570 680270
rect 152660 680030 152900 680270
rect 152990 680030 153230 680270
rect 153340 680030 153580 680270
rect 153670 680030 153910 680270
rect 154000 680030 154240 680270
rect 154330 680030 154570 680270
rect 154680 680030 154920 680270
rect 155010 680030 155250 680270
rect 155340 680030 155580 680270
rect 155670 680030 155910 680270
rect 144950 679700 145190 679940
rect 145300 679700 145540 679940
rect 145630 679700 145870 679940
rect 145960 679700 146200 679940
rect 146290 679700 146530 679940
rect 146640 679700 146880 679940
rect 146970 679700 147210 679940
rect 147300 679700 147540 679940
rect 147630 679700 147870 679940
rect 147980 679700 148220 679940
rect 148310 679700 148550 679940
rect 148640 679700 148880 679940
rect 148970 679700 149210 679940
rect 149320 679700 149560 679940
rect 149650 679700 149890 679940
rect 149980 679700 150220 679940
rect 150310 679700 150550 679940
rect 150660 679700 150900 679940
rect 150990 679700 151230 679940
rect 151320 679700 151560 679940
rect 151650 679700 151890 679940
rect 152000 679700 152240 679940
rect 152330 679700 152570 679940
rect 152660 679700 152900 679940
rect 152990 679700 153230 679940
rect 153340 679700 153580 679940
rect 153670 679700 153910 679940
rect 154000 679700 154240 679940
rect 154330 679700 154570 679940
rect 154680 679700 154920 679940
rect 155010 679700 155250 679940
rect 155340 679700 155580 679940
rect 155670 679700 155910 679940
rect 144950 679370 145190 679610
rect 145300 679370 145540 679610
rect 145630 679370 145870 679610
rect 145960 679370 146200 679610
rect 146290 679370 146530 679610
rect 146640 679370 146880 679610
rect 146970 679370 147210 679610
rect 147300 679370 147540 679610
rect 147630 679370 147870 679610
rect 147980 679370 148220 679610
rect 148310 679370 148550 679610
rect 148640 679370 148880 679610
rect 148970 679370 149210 679610
rect 149320 679370 149560 679610
rect 149650 679370 149890 679610
rect 149980 679370 150220 679610
rect 150310 679370 150550 679610
rect 150660 679370 150900 679610
rect 150990 679370 151230 679610
rect 151320 679370 151560 679610
rect 151650 679370 151890 679610
rect 152000 679370 152240 679610
rect 152330 679370 152570 679610
rect 152660 679370 152900 679610
rect 152990 679370 153230 679610
rect 153340 679370 153580 679610
rect 153670 679370 153910 679610
rect 154000 679370 154240 679610
rect 154330 679370 154570 679610
rect 154680 679370 154920 679610
rect 155010 679370 155250 679610
rect 155340 679370 155580 679610
rect 155670 679370 155910 679610
rect 144950 679020 145190 679260
rect 145300 679020 145540 679260
rect 145630 679020 145870 679260
rect 145960 679020 146200 679260
rect 146290 679020 146530 679260
rect 146640 679020 146880 679260
rect 146970 679020 147210 679260
rect 147300 679020 147540 679260
rect 147630 679020 147870 679260
rect 147980 679020 148220 679260
rect 148310 679020 148550 679260
rect 148640 679020 148880 679260
rect 148970 679020 149210 679260
rect 149320 679020 149560 679260
rect 149650 679020 149890 679260
rect 149980 679020 150220 679260
rect 150310 679020 150550 679260
rect 150660 679020 150900 679260
rect 150990 679020 151230 679260
rect 151320 679020 151560 679260
rect 151650 679020 151890 679260
rect 152000 679020 152240 679260
rect 152330 679020 152570 679260
rect 152660 679020 152900 679260
rect 152990 679020 153230 679260
rect 153340 679020 153580 679260
rect 153670 679020 153910 679260
rect 154000 679020 154240 679260
rect 154330 679020 154570 679260
rect 154680 679020 154920 679260
rect 155010 679020 155250 679260
rect 155340 679020 155580 679260
rect 155670 679020 155910 679260
rect 144950 678690 145190 678930
rect 145300 678690 145540 678930
rect 145630 678690 145870 678930
rect 145960 678690 146200 678930
rect 146290 678690 146530 678930
rect 146640 678690 146880 678930
rect 146970 678690 147210 678930
rect 147300 678690 147540 678930
rect 147630 678690 147870 678930
rect 147980 678690 148220 678930
rect 148310 678690 148550 678930
rect 148640 678690 148880 678930
rect 148970 678690 149210 678930
rect 149320 678690 149560 678930
rect 149650 678690 149890 678930
rect 149980 678690 150220 678930
rect 150310 678690 150550 678930
rect 150660 678690 150900 678930
rect 150990 678690 151230 678930
rect 151320 678690 151560 678930
rect 151650 678690 151890 678930
rect 152000 678690 152240 678930
rect 152330 678690 152570 678930
rect 152660 678690 152900 678930
rect 152990 678690 153230 678930
rect 153340 678690 153580 678930
rect 153670 678690 153910 678930
rect 154000 678690 154240 678930
rect 154330 678690 154570 678930
rect 154680 678690 154920 678930
rect 155010 678690 155250 678930
rect 155340 678690 155580 678930
rect 155670 678690 155910 678930
rect 144950 678360 145190 678600
rect 145300 678360 145540 678600
rect 145630 678360 145870 678600
rect 145960 678360 146200 678600
rect 146290 678360 146530 678600
rect 146640 678360 146880 678600
rect 146970 678360 147210 678600
rect 147300 678360 147540 678600
rect 147630 678360 147870 678600
rect 147980 678360 148220 678600
rect 148310 678360 148550 678600
rect 148640 678360 148880 678600
rect 148970 678360 149210 678600
rect 149320 678360 149560 678600
rect 149650 678360 149890 678600
rect 149980 678360 150220 678600
rect 150310 678360 150550 678600
rect 150660 678360 150900 678600
rect 150990 678360 151230 678600
rect 151320 678360 151560 678600
rect 151650 678360 151890 678600
rect 152000 678360 152240 678600
rect 152330 678360 152570 678600
rect 152660 678360 152900 678600
rect 152990 678360 153230 678600
rect 153340 678360 153580 678600
rect 153670 678360 153910 678600
rect 154000 678360 154240 678600
rect 154330 678360 154570 678600
rect 154680 678360 154920 678600
rect 155010 678360 155250 678600
rect 155340 678360 155580 678600
rect 155670 678360 155910 678600
rect 144950 678030 145190 678270
rect 145300 678030 145540 678270
rect 145630 678030 145870 678270
rect 145960 678030 146200 678270
rect 146290 678030 146530 678270
rect 146640 678030 146880 678270
rect 146970 678030 147210 678270
rect 147300 678030 147540 678270
rect 147630 678030 147870 678270
rect 147980 678030 148220 678270
rect 148310 678030 148550 678270
rect 148640 678030 148880 678270
rect 148970 678030 149210 678270
rect 149320 678030 149560 678270
rect 149650 678030 149890 678270
rect 149980 678030 150220 678270
rect 150310 678030 150550 678270
rect 150660 678030 150900 678270
rect 150990 678030 151230 678270
rect 151320 678030 151560 678270
rect 151650 678030 151890 678270
rect 152000 678030 152240 678270
rect 152330 678030 152570 678270
rect 152660 678030 152900 678270
rect 152990 678030 153230 678270
rect 153340 678030 153580 678270
rect 153670 678030 153910 678270
rect 154000 678030 154240 678270
rect 154330 678030 154570 678270
rect 154680 678030 154920 678270
rect 155010 678030 155250 678270
rect 155340 678030 155580 678270
rect 155670 678030 155910 678270
rect 144950 677680 145190 677920
rect 145300 677680 145540 677920
rect 145630 677680 145870 677920
rect 145960 677680 146200 677920
rect 146290 677680 146530 677920
rect 146640 677680 146880 677920
rect 146970 677680 147210 677920
rect 147300 677680 147540 677920
rect 147630 677680 147870 677920
rect 147980 677680 148220 677920
rect 148310 677680 148550 677920
rect 148640 677680 148880 677920
rect 148970 677680 149210 677920
rect 149320 677680 149560 677920
rect 149650 677680 149890 677920
rect 149980 677680 150220 677920
rect 150310 677680 150550 677920
rect 150660 677680 150900 677920
rect 150990 677680 151230 677920
rect 151320 677680 151560 677920
rect 151650 677680 151890 677920
rect 152000 677680 152240 677920
rect 152330 677680 152570 677920
rect 152660 677680 152900 677920
rect 152990 677680 153230 677920
rect 153340 677680 153580 677920
rect 153670 677680 153910 677920
rect 154000 677680 154240 677920
rect 154330 677680 154570 677920
rect 154680 677680 154920 677920
rect 155010 677680 155250 677920
rect 155340 677680 155580 677920
rect 155670 677680 155910 677920
rect 144950 677350 145190 677590
rect 145300 677350 145540 677590
rect 145630 677350 145870 677590
rect 145960 677350 146200 677590
rect 146290 677350 146530 677590
rect 146640 677350 146880 677590
rect 146970 677350 147210 677590
rect 147300 677350 147540 677590
rect 147630 677350 147870 677590
rect 147980 677350 148220 677590
rect 148310 677350 148550 677590
rect 148640 677350 148880 677590
rect 148970 677350 149210 677590
rect 149320 677350 149560 677590
rect 149650 677350 149890 677590
rect 149980 677350 150220 677590
rect 150310 677350 150550 677590
rect 150660 677350 150900 677590
rect 150990 677350 151230 677590
rect 151320 677350 151560 677590
rect 151650 677350 151890 677590
rect 152000 677350 152240 677590
rect 152330 677350 152570 677590
rect 152660 677350 152900 677590
rect 152990 677350 153230 677590
rect 153340 677350 153580 677590
rect 153670 677350 153910 677590
rect 154000 677350 154240 677590
rect 154330 677350 154570 677590
rect 154680 677350 154920 677590
rect 155010 677350 155250 677590
rect 155340 677350 155580 677590
rect 155670 677350 155910 677590
rect 144950 677020 145190 677260
rect 145300 677020 145540 677260
rect 145630 677020 145870 677260
rect 145960 677020 146200 677260
rect 146290 677020 146530 677260
rect 146640 677020 146880 677260
rect 146970 677020 147210 677260
rect 147300 677020 147540 677260
rect 147630 677020 147870 677260
rect 147980 677020 148220 677260
rect 148310 677020 148550 677260
rect 148640 677020 148880 677260
rect 148970 677020 149210 677260
rect 149320 677020 149560 677260
rect 149650 677020 149890 677260
rect 149980 677020 150220 677260
rect 150310 677020 150550 677260
rect 150660 677020 150900 677260
rect 150990 677020 151230 677260
rect 151320 677020 151560 677260
rect 151650 677020 151890 677260
rect 152000 677020 152240 677260
rect 152330 677020 152570 677260
rect 152660 677020 152900 677260
rect 152990 677020 153230 677260
rect 153340 677020 153580 677260
rect 153670 677020 153910 677260
rect 154000 677020 154240 677260
rect 154330 677020 154570 677260
rect 154680 677020 154920 677260
rect 155010 677020 155250 677260
rect 155340 677020 155580 677260
rect 155670 677020 155910 677260
rect 144950 676690 145190 676930
rect 145300 676690 145540 676930
rect 145630 676690 145870 676930
rect 145960 676690 146200 676930
rect 146290 676690 146530 676930
rect 146640 676690 146880 676930
rect 146970 676690 147210 676930
rect 147300 676690 147540 676930
rect 147630 676690 147870 676930
rect 147980 676690 148220 676930
rect 148310 676690 148550 676930
rect 148640 676690 148880 676930
rect 148970 676690 149210 676930
rect 149320 676690 149560 676930
rect 149650 676690 149890 676930
rect 149980 676690 150220 676930
rect 150310 676690 150550 676930
rect 150660 676690 150900 676930
rect 150990 676690 151230 676930
rect 151320 676690 151560 676930
rect 151650 676690 151890 676930
rect 152000 676690 152240 676930
rect 152330 676690 152570 676930
rect 152660 676690 152900 676930
rect 152990 676690 153230 676930
rect 153340 676690 153580 676930
rect 153670 676690 153910 676930
rect 154000 676690 154240 676930
rect 154330 676690 154570 676930
rect 154680 676690 154920 676930
rect 155010 676690 155250 676930
rect 155340 676690 155580 676930
rect 155670 676690 155910 676930
rect 144950 676340 145190 676580
rect 145300 676340 145540 676580
rect 145630 676340 145870 676580
rect 145960 676340 146200 676580
rect 146290 676340 146530 676580
rect 146640 676340 146880 676580
rect 146970 676340 147210 676580
rect 147300 676340 147540 676580
rect 147630 676340 147870 676580
rect 147980 676340 148220 676580
rect 148310 676340 148550 676580
rect 148640 676340 148880 676580
rect 148970 676340 149210 676580
rect 149320 676340 149560 676580
rect 149650 676340 149890 676580
rect 149980 676340 150220 676580
rect 150310 676340 150550 676580
rect 150660 676340 150900 676580
rect 150990 676340 151230 676580
rect 151320 676340 151560 676580
rect 151650 676340 151890 676580
rect 152000 676340 152240 676580
rect 152330 676340 152570 676580
rect 152660 676340 152900 676580
rect 152990 676340 153230 676580
rect 153340 676340 153580 676580
rect 153670 676340 153910 676580
rect 154000 676340 154240 676580
rect 154330 676340 154570 676580
rect 154680 676340 154920 676580
rect 155010 676340 155250 676580
rect 155340 676340 155580 676580
rect 155670 676340 155910 676580
rect 144950 676010 145190 676250
rect 145300 676010 145540 676250
rect 145630 676010 145870 676250
rect 145960 676010 146200 676250
rect 146290 676010 146530 676250
rect 146640 676010 146880 676250
rect 146970 676010 147210 676250
rect 147300 676010 147540 676250
rect 147630 676010 147870 676250
rect 147980 676010 148220 676250
rect 148310 676010 148550 676250
rect 148640 676010 148880 676250
rect 148970 676010 149210 676250
rect 149320 676010 149560 676250
rect 149650 676010 149890 676250
rect 149980 676010 150220 676250
rect 150310 676010 150550 676250
rect 150660 676010 150900 676250
rect 150990 676010 151230 676250
rect 151320 676010 151560 676250
rect 151650 676010 151890 676250
rect 152000 676010 152240 676250
rect 152330 676010 152570 676250
rect 152660 676010 152900 676250
rect 152990 676010 153230 676250
rect 153340 676010 153580 676250
rect 153670 676010 153910 676250
rect 154000 676010 154240 676250
rect 154330 676010 154570 676250
rect 154680 676010 154920 676250
rect 155010 676010 155250 676250
rect 155340 676010 155580 676250
rect 155670 676010 155910 676250
rect 144950 675680 145190 675920
rect 145300 675680 145540 675920
rect 145630 675680 145870 675920
rect 145960 675680 146200 675920
rect 146290 675680 146530 675920
rect 146640 675680 146880 675920
rect 146970 675680 147210 675920
rect 147300 675680 147540 675920
rect 147630 675680 147870 675920
rect 147980 675680 148220 675920
rect 148310 675680 148550 675920
rect 148640 675680 148880 675920
rect 148970 675680 149210 675920
rect 149320 675680 149560 675920
rect 149650 675680 149890 675920
rect 149980 675680 150220 675920
rect 150310 675680 150550 675920
rect 150660 675680 150900 675920
rect 150990 675680 151230 675920
rect 151320 675680 151560 675920
rect 151650 675680 151890 675920
rect 152000 675680 152240 675920
rect 152330 675680 152570 675920
rect 152660 675680 152900 675920
rect 152990 675680 153230 675920
rect 153340 675680 153580 675920
rect 153670 675680 153910 675920
rect 154000 675680 154240 675920
rect 154330 675680 154570 675920
rect 154680 675680 154920 675920
rect 155010 675680 155250 675920
rect 155340 675680 155580 675920
rect 155670 675680 155910 675920
rect 144950 675350 145190 675590
rect 145300 675350 145540 675590
rect 145630 675350 145870 675590
rect 145960 675350 146200 675590
rect 146290 675350 146530 675590
rect 146640 675350 146880 675590
rect 146970 675350 147210 675590
rect 147300 675350 147540 675590
rect 147630 675350 147870 675590
rect 147980 675350 148220 675590
rect 148310 675350 148550 675590
rect 148640 675350 148880 675590
rect 148970 675350 149210 675590
rect 149320 675350 149560 675590
rect 149650 675350 149890 675590
rect 149980 675350 150220 675590
rect 150310 675350 150550 675590
rect 150660 675350 150900 675590
rect 150990 675350 151230 675590
rect 151320 675350 151560 675590
rect 151650 675350 151890 675590
rect 152000 675350 152240 675590
rect 152330 675350 152570 675590
rect 152660 675350 152900 675590
rect 152990 675350 153230 675590
rect 153340 675350 153580 675590
rect 153670 675350 153910 675590
rect 154000 675350 154240 675590
rect 154330 675350 154570 675590
rect 154680 675350 154920 675590
rect 155010 675350 155250 675590
rect 155340 675350 155580 675590
rect 155670 675350 155910 675590
rect 144950 675000 145190 675240
rect 145300 675000 145540 675240
rect 145630 675000 145870 675240
rect 145960 675000 146200 675240
rect 146290 675000 146530 675240
rect 146640 675000 146880 675240
rect 146970 675000 147210 675240
rect 147300 675000 147540 675240
rect 147630 675000 147870 675240
rect 147980 675000 148220 675240
rect 148310 675000 148550 675240
rect 148640 675000 148880 675240
rect 148970 675000 149210 675240
rect 149320 675000 149560 675240
rect 149650 675000 149890 675240
rect 149980 675000 150220 675240
rect 150310 675000 150550 675240
rect 150660 675000 150900 675240
rect 150990 675000 151230 675240
rect 151320 675000 151560 675240
rect 151650 675000 151890 675240
rect 152000 675000 152240 675240
rect 152330 675000 152570 675240
rect 152660 675000 152900 675240
rect 152990 675000 153230 675240
rect 153340 675000 153580 675240
rect 153670 675000 153910 675240
rect 154000 675000 154240 675240
rect 154330 675000 154570 675240
rect 154680 675000 154920 675240
rect 155010 675000 155250 675240
rect 155340 675000 155580 675240
rect 155670 675000 155910 675240
rect 144950 674670 145190 674910
rect 145300 674670 145540 674910
rect 145630 674670 145870 674910
rect 145960 674670 146200 674910
rect 146290 674670 146530 674910
rect 146640 674670 146880 674910
rect 146970 674670 147210 674910
rect 147300 674670 147540 674910
rect 147630 674670 147870 674910
rect 147980 674670 148220 674910
rect 148310 674670 148550 674910
rect 148640 674670 148880 674910
rect 148970 674670 149210 674910
rect 149320 674670 149560 674910
rect 149650 674670 149890 674910
rect 149980 674670 150220 674910
rect 150310 674670 150550 674910
rect 150660 674670 150900 674910
rect 150990 674670 151230 674910
rect 151320 674670 151560 674910
rect 151650 674670 151890 674910
rect 152000 674670 152240 674910
rect 152330 674670 152570 674910
rect 152660 674670 152900 674910
rect 152990 674670 153230 674910
rect 153340 674670 153580 674910
rect 153670 674670 153910 674910
rect 154000 674670 154240 674910
rect 154330 674670 154570 674910
rect 154680 674670 154920 674910
rect 155010 674670 155250 674910
rect 155340 674670 155580 674910
rect 155670 674670 155910 674910
rect 144950 674340 145190 674580
rect 145300 674340 145540 674580
rect 145630 674340 145870 674580
rect 145960 674340 146200 674580
rect 146290 674340 146530 674580
rect 146640 674340 146880 674580
rect 146970 674340 147210 674580
rect 147300 674340 147540 674580
rect 147630 674340 147870 674580
rect 147980 674340 148220 674580
rect 148310 674340 148550 674580
rect 148640 674340 148880 674580
rect 148970 674340 149210 674580
rect 149320 674340 149560 674580
rect 149650 674340 149890 674580
rect 149980 674340 150220 674580
rect 150310 674340 150550 674580
rect 150660 674340 150900 674580
rect 150990 674340 151230 674580
rect 151320 674340 151560 674580
rect 151650 674340 151890 674580
rect 152000 674340 152240 674580
rect 152330 674340 152570 674580
rect 152660 674340 152900 674580
rect 152990 674340 153230 674580
rect 153340 674340 153580 674580
rect 153670 674340 153910 674580
rect 154000 674340 154240 674580
rect 154330 674340 154570 674580
rect 154680 674340 154920 674580
rect 155010 674340 155250 674580
rect 155340 674340 155580 674580
rect 155670 674340 155910 674580
rect 144950 674010 145190 674250
rect 145300 674010 145540 674250
rect 145630 674010 145870 674250
rect 145960 674010 146200 674250
rect 146290 674010 146530 674250
rect 146640 674010 146880 674250
rect 146970 674010 147210 674250
rect 147300 674010 147540 674250
rect 147630 674010 147870 674250
rect 147980 674010 148220 674250
rect 148310 674010 148550 674250
rect 148640 674010 148880 674250
rect 148970 674010 149210 674250
rect 149320 674010 149560 674250
rect 149650 674010 149890 674250
rect 149980 674010 150220 674250
rect 150310 674010 150550 674250
rect 150660 674010 150900 674250
rect 150990 674010 151230 674250
rect 151320 674010 151560 674250
rect 151650 674010 151890 674250
rect 152000 674010 152240 674250
rect 152330 674010 152570 674250
rect 152660 674010 152900 674250
rect 152990 674010 153230 674250
rect 153340 674010 153580 674250
rect 153670 674010 153910 674250
rect 154000 674010 154240 674250
rect 154330 674010 154570 674250
rect 154680 674010 154920 674250
rect 155010 674010 155250 674250
rect 155340 674010 155580 674250
rect 155670 674010 155910 674250
rect 144950 673660 145190 673900
rect 145300 673660 145540 673900
rect 145630 673660 145870 673900
rect 145960 673660 146200 673900
rect 146290 673660 146530 673900
rect 146640 673660 146880 673900
rect 146970 673660 147210 673900
rect 147300 673660 147540 673900
rect 147630 673660 147870 673900
rect 147980 673660 148220 673900
rect 148310 673660 148550 673900
rect 148640 673660 148880 673900
rect 148970 673660 149210 673900
rect 149320 673660 149560 673900
rect 149650 673660 149890 673900
rect 149980 673660 150220 673900
rect 150310 673660 150550 673900
rect 150660 673660 150900 673900
rect 150990 673660 151230 673900
rect 151320 673660 151560 673900
rect 151650 673660 151890 673900
rect 152000 673660 152240 673900
rect 152330 673660 152570 673900
rect 152660 673660 152900 673900
rect 152990 673660 153230 673900
rect 153340 673660 153580 673900
rect 153670 673660 153910 673900
rect 154000 673660 154240 673900
rect 154330 673660 154570 673900
rect 154680 673660 154920 673900
rect 155010 673660 155250 673900
rect 155340 673660 155580 673900
rect 155670 673660 155910 673900
rect 144950 673330 145190 673570
rect 145300 673330 145540 673570
rect 145630 673330 145870 673570
rect 145960 673330 146200 673570
rect 146290 673330 146530 673570
rect 146640 673330 146880 673570
rect 146970 673330 147210 673570
rect 147300 673330 147540 673570
rect 147630 673330 147870 673570
rect 147980 673330 148220 673570
rect 148310 673330 148550 673570
rect 148640 673330 148880 673570
rect 148970 673330 149210 673570
rect 149320 673330 149560 673570
rect 149650 673330 149890 673570
rect 149980 673330 150220 673570
rect 150310 673330 150550 673570
rect 150660 673330 150900 673570
rect 150990 673330 151230 673570
rect 151320 673330 151560 673570
rect 151650 673330 151890 673570
rect 152000 673330 152240 673570
rect 152330 673330 152570 673570
rect 152660 673330 152900 673570
rect 152990 673330 153230 673570
rect 153340 673330 153580 673570
rect 153670 673330 153910 673570
rect 154000 673330 154240 673570
rect 154330 673330 154570 673570
rect 154680 673330 154920 673570
rect 155010 673330 155250 673570
rect 155340 673330 155580 673570
rect 155670 673330 155910 673570
rect 144950 673000 145190 673240
rect 145300 673000 145540 673240
rect 145630 673000 145870 673240
rect 145960 673000 146200 673240
rect 146290 673000 146530 673240
rect 146640 673000 146880 673240
rect 146970 673000 147210 673240
rect 147300 673000 147540 673240
rect 147630 673000 147870 673240
rect 147980 673000 148220 673240
rect 148310 673000 148550 673240
rect 148640 673000 148880 673240
rect 148970 673000 149210 673240
rect 149320 673000 149560 673240
rect 149650 673000 149890 673240
rect 149980 673000 150220 673240
rect 150310 673000 150550 673240
rect 150660 673000 150900 673240
rect 150990 673000 151230 673240
rect 151320 673000 151560 673240
rect 151650 673000 151890 673240
rect 152000 673000 152240 673240
rect 152330 673000 152570 673240
rect 152660 673000 152900 673240
rect 152990 673000 153230 673240
rect 153340 673000 153580 673240
rect 153670 673000 153910 673240
rect 154000 673000 154240 673240
rect 154330 673000 154570 673240
rect 154680 673000 154920 673240
rect 155010 673000 155250 673240
rect 155340 673000 155580 673240
rect 155670 673000 155910 673240
rect 144950 672670 145190 672910
rect 145300 672670 145540 672910
rect 145630 672670 145870 672910
rect 145960 672670 146200 672910
rect 146290 672670 146530 672910
rect 146640 672670 146880 672910
rect 146970 672670 147210 672910
rect 147300 672670 147540 672910
rect 147630 672670 147870 672910
rect 147980 672670 148220 672910
rect 148310 672670 148550 672910
rect 148640 672670 148880 672910
rect 148970 672670 149210 672910
rect 149320 672670 149560 672910
rect 149650 672670 149890 672910
rect 149980 672670 150220 672910
rect 150310 672670 150550 672910
rect 150660 672670 150900 672910
rect 150990 672670 151230 672910
rect 151320 672670 151560 672910
rect 151650 672670 151890 672910
rect 152000 672670 152240 672910
rect 152330 672670 152570 672910
rect 152660 672670 152900 672910
rect 152990 672670 153230 672910
rect 153340 672670 153580 672910
rect 153670 672670 153910 672910
rect 154000 672670 154240 672910
rect 154330 672670 154570 672910
rect 154680 672670 154920 672910
rect 155010 672670 155250 672910
rect 155340 672670 155580 672910
rect 155670 672670 155910 672910
rect 144950 672320 145190 672560
rect 145300 672320 145540 672560
rect 145630 672320 145870 672560
rect 145960 672320 146200 672560
rect 146290 672320 146530 672560
rect 146640 672320 146880 672560
rect 146970 672320 147210 672560
rect 147300 672320 147540 672560
rect 147630 672320 147870 672560
rect 147980 672320 148220 672560
rect 148310 672320 148550 672560
rect 148640 672320 148880 672560
rect 148970 672320 149210 672560
rect 149320 672320 149560 672560
rect 149650 672320 149890 672560
rect 149980 672320 150220 672560
rect 150310 672320 150550 672560
rect 150660 672320 150900 672560
rect 150990 672320 151230 672560
rect 151320 672320 151560 672560
rect 151650 672320 151890 672560
rect 152000 672320 152240 672560
rect 152330 672320 152570 672560
rect 152660 672320 152900 672560
rect 152990 672320 153230 672560
rect 153340 672320 153580 672560
rect 153670 672320 153910 672560
rect 154000 672320 154240 672560
rect 154330 672320 154570 672560
rect 154680 672320 154920 672560
rect 155010 672320 155250 672560
rect 155340 672320 155580 672560
rect 155670 672320 155910 672560
rect 110810 671660 111050 671900
rect 111140 671660 111380 671900
rect 111470 671660 111710 671900
rect 111800 671660 112040 671900
rect 112150 671660 112390 671900
rect 112480 671660 112720 671900
rect 112810 671660 113050 671900
rect 113140 671660 113380 671900
rect 113490 671660 113730 671900
rect 113820 671660 114060 671900
rect 114150 671660 114390 671900
rect 114480 671660 114720 671900
rect 114830 671660 115070 671900
rect 115160 671660 115400 671900
rect 115490 671660 115730 671900
rect 115820 671660 116060 671900
rect 116170 671660 116410 671900
rect 116500 671660 116740 671900
rect 116830 671660 117070 671900
rect 117160 671660 117400 671900
rect 117510 671660 117750 671900
rect 117840 671660 118080 671900
rect 118170 671660 118410 671900
rect 118500 671660 118740 671900
rect 118850 671660 119090 671900
rect 119180 671660 119420 671900
rect 119510 671660 119750 671900
rect 119840 671660 120080 671900
rect 120190 671660 120430 671900
rect 120520 671660 120760 671900
rect 120850 671660 121090 671900
rect 121180 671660 121420 671900
rect 121530 671660 121770 671900
rect 110810 671310 111050 671550
rect 111140 671310 111380 671550
rect 111470 671310 111710 671550
rect 111800 671310 112040 671550
rect 112150 671310 112390 671550
rect 112480 671310 112720 671550
rect 112810 671310 113050 671550
rect 113140 671310 113380 671550
rect 113490 671310 113730 671550
rect 113820 671310 114060 671550
rect 114150 671310 114390 671550
rect 114480 671310 114720 671550
rect 114830 671310 115070 671550
rect 115160 671310 115400 671550
rect 115490 671310 115730 671550
rect 115820 671310 116060 671550
rect 116170 671310 116410 671550
rect 116500 671310 116740 671550
rect 116830 671310 117070 671550
rect 117160 671310 117400 671550
rect 117510 671310 117750 671550
rect 117840 671310 118080 671550
rect 118170 671310 118410 671550
rect 118500 671310 118740 671550
rect 118850 671310 119090 671550
rect 119180 671310 119420 671550
rect 119510 671310 119750 671550
rect 119840 671310 120080 671550
rect 120190 671310 120430 671550
rect 120520 671310 120760 671550
rect 120850 671310 121090 671550
rect 121180 671310 121420 671550
rect 121530 671310 121770 671550
rect 110810 670980 111050 671220
rect 111140 670980 111380 671220
rect 111470 670980 111710 671220
rect 111800 670980 112040 671220
rect 112150 670980 112390 671220
rect 112480 670980 112720 671220
rect 112810 670980 113050 671220
rect 113140 670980 113380 671220
rect 113490 670980 113730 671220
rect 113820 670980 114060 671220
rect 114150 670980 114390 671220
rect 114480 670980 114720 671220
rect 114830 670980 115070 671220
rect 115160 670980 115400 671220
rect 115490 670980 115730 671220
rect 115820 670980 116060 671220
rect 116170 670980 116410 671220
rect 116500 670980 116740 671220
rect 116830 670980 117070 671220
rect 117160 670980 117400 671220
rect 117510 670980 117750 671220
rect 117840 670980 118080 671220
rect 118170 670980 118410 671220
rect 118500 670980 118740 671220
rect 118850 670980 119090 671220
rect 119180 670980 119420 671220
rect 119510 670980 119750 671220
rect 119840 670980 120080 671220
rect 120190 670980 120430 671220
rect 120520 670980 120760 671220
rect 120850 670980 121090 671220
rect 121180 670980 121420 671220
rect 121530 670980 121770 671220
rect 110810 670650 111050 670890
rect 111140 670650 111380 670890
rect 111470 670650 111710 670890
rect 111800 670650 112040 670890
rect 112150 670650 112390 670890
rect 112480 670650 112720 670890
rect 112810 670650 113050 670890
rect 113140 670650 113380 670890
rect 113490 670650 113730 670890
rect 113820 670650 114060 670890
rect 114150 670650 114390 670890
rect 114480 670650 114720 670890
rect 114830 670650 115070 670890
rect 115160 670650 115400 670890
rect 115490 670650 115730 670890
rect 115820 670650 116060 670890
rect 116170 670650 116410 670890
rect 116500 670650 116740 670890
rect 116830 670650 117070 670890
rect 117160 670650 117400 670890
rect 117510 670650 117750 670890
rect 117840 670650 118080 670890
rect 118170 670650 118410 670890
rect 118500 670650 118740 670890
rect 118850 670650 119090 670890
rect 119180 670650 119420 670890
rect 119510 670650 119750 670890
rect 119840 670650 120080 670890
rect 120190 670650 120430 670890
rect 120520 670650 120760 670890
rect 120850 670650 121090 670890
rect 121180 670650 121420 670890
rect 121530 670650 121770 670890
rect 110810 670320 111050 670560
rect 111140 670320 111380 670560
rect 111470 670320 111710 670560
rect 111800 670320 112040 670560
rect 112150 670320 112390 670560
rect 112480 670320 112720 670560
rect 112810 670320 113050 670560
rect 113140 670320 113380 670560
rect 113490 670320 113730 670560
rect 113820 670320 114060 670560
rect 114150 670320 114390 670560
rect 114480 670320 114720 670560
rect 114830 670320 115070 670560
rect 115160 670320 115400 670560
rect 115490 670320 115730 670560
rect 115820 670320 116060 670560
rect 116170 670320 116410 670560
rect 116500 670320 116740 670560
rect 116830 670320 117070 670560
rect 117160 670320 117400 670560
rect 117510 670320 117750 670560
rect 117840 670320 118080 670560
rect 118170 670320 118410 670560
rect 118500 670320 118740 670560
rect 118850 670320 119090 670560
rect 119180 670320 119420 670560
rect 119510 670320 119750 670560
rect 119840 670320 120080 670560
rect 120190 670320 120430 670560
rect 120520 670320 120760 670560
rect 120850 670320 121090 670560
rect 121180 670320 121420 670560
rect 121530 670320 121770 670560
rect 110810 669970 111050 670210
rect 111140 669970 111380 670210
rect 111470 669970 111710 670210
rect 111800 669970 112040 670210
rect 112150 669970 112390 670210
rect 112480 669970 112720 670210
rect 112810 669970 113050 670210
rect 113140 669970 113380 670210
rect 113490 669970 113730 670210
rect 113820 669970 114060 670210
rect 114150 669970 114390 670210
rect 114480 669970 114720 670210
rect 114830 669970 115070 670210
rect 115160 669970 115400 670210
rect 115490 669970 115730 670210
rect 115820 669970 116060 670210
rect 116170 669970 116410 670210
rect 116500 669970 116740 670210
rect 116830 669970 117070 670210
rect 117160 669970 117400 670210
rect 117510 669970 117750 670210
rect 117840 669970 118080 670210
rect 118170 669970 118410 670210
rect 118500 669970 118740 670210
rect 118850 669970 119090 670210
rect 119180 669970 119420 670210
rect 119510 669970 119750 670210
rect 119840 669970 120080 670210
rect 120190 669970 120430 670210
rect 120520 669970 120760 670210
rect 120850 669970 121090 670210
rect 121180 669970 121420 670210
rect 121530 669970 121770 670210
rect 110810 669640 111050 669880
rect 111140 669640 111380 669880
rect 111470 669640 111710 669880
rect 111800 669640 112040 669880
rect 112150 669640 112390 669880
rect 112480 669640 112720 669880
rect 112810 669640 113050 669880
rect 113140 669640 113380 669880
rect 113490 669640 113730 669880
rect 113820 669640 114060 669880
rect 114150 669640 114390 669880
rect 114480 669640 114720 669880
rect 114830 669640 115070 669880
rect 115160 669640 115400 669880
rect 115490 669640 115730 669880
rect 115820 669640 116060 669880
rect 116170 669640 116410 669880
rect 116500 669640 116740 669880
rect 116830 669640 117070 669880
rect 117160 669640 117400 669880
rect 117510 669640 117750 669880
rect 117840 669640 118080 669880
rect 118170 669640 118410 669880
rect 118500 669640 118740 669880
rect 118850 669640 119090 669880
rect 119180 669640 119420 669880
rect 119510 669640 119750 669880
rect 119840 669640 120080 669880
rect 120190 669640 120430 669880
rect 120520 669640 120760 669880
rect 120850 669640 121090 669880
rect 121180 669640 121420 669880
rect 121530 669640 121770 669880
rect 110810 669310 111050 669550
rect 111140 669310 111380 669550
rect 111470 669310 111710 669550
rect 111800 669310 112040 669550
rect 112150 669310 112390 669550
rect 112480 669310 112720 669550
rect 112810 669310 113050 669550
rect 113140 669310 113380 669550
rect 113490 669310 113730 669550
rect 113820 669310 114060 669550
rect 114150 669310 114390 669550
rect 114480 669310 114720 669550
rect 114830 669310 115070 669550
rect 115160 669310 115400 669550
rect 115490 669310 115730 669550
rect 115820 669310 116060 669550
rect 116170 669310 116410 669550
rect 116500 669310 116740 669550
rect 116830 669310 117070 669550
rect 117160 669310 117400 669550
rect 117510 669310 117750 669550
rect 117840 669310 118080 669550
rect 118170 669310 118410 669550
rect 118500 669310 118740 669550
rect 118850 669310 119090 669550
rect 119180 669310 119420 669550
rect 119510 669310 119750 669550
rect 119840 669310 120080 669550
rect 120190 669310 120430 669550
rect 120520 669310 120760 669550
rect 120850 669310 121090 669550
rect 121180 669310 121420 669550
rect 121530 669310 121770 669550
rect 110810 668980 111050 669220
rect 111140 668980 111380 669220
rect 111470 668980 111710 669220
rect 111800 668980 112040 669220
rect 112150 668980 112390 669220
rect 112480 668980 112720 669220
rect 112810 668980 113050 669220
rect 113140 668980 113380 669220
rect 113490 668980 113730 669220
rect 113820 668980 114060 669220
rect 114150 668980 114390 669220
rect 114480 668980 114720 669220
rect 114830 668980 115070 669220
rect 115160 668980 115400 669220
rect 115490 668980 115730 669220
rect 115820 668980 116060 669220
rect 116170 668980 116410 669220
rect 116500 668980 116740 669220
rect 116830 668980 117070 669220
rect 117160 668980 117400 669220
rect 117510 668980 117750 669220
rect 117840 668980 118080 669220
rect 118170 668980 118410 669220
rect 118500 668980 118740 669220
rect 118850 668980 119090 669220
rect 119180 668980 119420 669220
rect 119510 668980 119750 669220
rect 119840 668980 120080 669220
rect 120190 668980 120430 669220
rect 120520 668980 120760 669220
rect 120850 668980 121090 669220
rect 121180 668980 121420 669220
rect 121530 668980 121770 669220
rect 110810 668630 111050 668870
rect 111140 668630 111380 668870
rect 111470 668630 111710 668870
rect 111800 668630 112040 668870
rect 112150 668630 112390 668870
rect 112480 668630 112720 668870
rect 112810 668630 113050 668870
rect 113140 668630 113380 668870
rect 113490 668630 113730 668870
rect 113820 668630 114060 668870
rect 114150 668630 114390 668870
rect 114480 668630 114720 668870
rect 114830 668630 115070 668870
rect 115160 668630 115400 668870
rect 115490 668630 115730 668870
rect 115820 668630 116060 668870
rect 116170 668630 116410 668870
rect 116500 668630 116740 668870
rect 116830 668630 117070 668870
rect 117160 668630 117400 668870
rect 117510 668630 117750 668870
rect 117840 668630 118080 668870
rect 118170 668630 118410 668870
rect 118500 668630 118740 668870
rect 118850 668630 119090 668870
rect 119180 668630 119420 668870
rect 119510 668630 119750 668870
rect 119840 668630 120080 668870
rect 120190 668630 120430 668870
rect 120520 668630 120760 668870
rect 120850 668630 121090 668870
rect 121180 668630 121420 668870
rect 121530 668630 121770 668870
rect 110810 668300 111050 668540
rect 111140 668300 111380 668540
rect 111470 668300 111710 668540
rect 111800 668300 112040 668540
rect 112150 668300 112390 668540
rect 112480 668300 112720 668540
rect 112810 668300 113050 668540
rect 113140 668300 113380 668540
rect 113490 668300 113730 668540
rect 113820 668300 114060 668540
rect 114150 668300 114390 668540
rect 114480 668300 114720 668540
rect 114830 668300 115070 668540
rect 115160 668300 115400 668540
rect 115490 668300 115730 668540
rect 115820 668300 116060 668540
rect 116170 668300 116410 668540
rect 116500 668300 116740 668540
rect 116830 668300 117070 668540
rect 117160 668300 117400 668540
rect 117510 668300 117750 668540
rect 117840 668300 118080 668540
rect 118170 668300 118410 668540
rect 118500 668300 118740 668540
rect 118850 668300 119090 668540
rect 119180 668300 119420 668540
rect 119510 668300 119750 668540
rect 119840 668300 120080 668540
rect 120190 668300 120430 668540
rect 120520 668300 120760 668540
rect 120850 668300 121090 668540
rect 121180 668300 121420 668540
rect 121530 668300 121770 668540
rect 110810 667970 111050 668210
rect 111140 667970 111380 668210
rect 111470 667970 111710 668210
rect 111800 667970 112040 668210
rect 112150 667970 112390 668210
rect 112480 667970 112720 668210
rect 112810 667970 113050 668210
rect 113140 667970 113380 668210
rect 113490 667970 113730 668210
rect 113820 667970 114060 668210
rect 114150 667970 114390 668210
rect 114480 667970 114720 668210
rect 114830 667970 115070 668210
rect 115160 667970 115400 668210
rect 115490 667970 115730 668210
rect 115820 667970 116060 668210
rect 116170 667970 116410 668210
rect 116500 667970 116740 668210
rect 116830 667970 117070 668210
rect 117160 667970 117400 668210
rect 117510 667970 117750 668210
rect 117840 667970 118080 668210
rect 118170 667970 118410 668210
rect 118500 667970 118740 668210
rect 118850 667970 119090 668210
rect 119180 667970 119420 668210
rect 119510 667970 119750 668210
rect 119840 667970 120080 668210
rect 120190 667970 120430 668210
rect 120520 667970 120760 668210
rect 120850 667970 121090 668210
rect 121180 667970 121420 668210
rect 121530 667970 121770 668210
rect 110810 667640 111050 667880
rect 111140 667640 111380 667880
rect 111470 667640 111710 667880
rect 111800 667640 112040 667880
rect 112150 667640 112390 667880
rect 112480 667640 112720 667880
rect 112810 667640 113050 667880
rect 113140 667640 113380 667880
rect 113490 667640 113730 667880
rect 113820 667640 114060 667880
rect 114150 667640 114390 667880
rect 114480 667640 114720 667880
rect 114830 667640 115070 667880
rect 115160 667640 115400 667880
rect 115490 667640 115730 667880
rect 115820 667640 116060 667880
rect 116170 667640 116410 667880
rect 116500 667640 116740 667880
rect 116830 667640 117070 667880
rect 117160 667640 117400 667880
rect 117510 667640 117750 667880
rect 117840 667640 118080 667880
rect 118170 667640 118410 667880
rect 118500 667640 118740 667880
rect 118850 667640 119090 667880
rect 119180 667640 119420 667880
rect 119510 667640 119750 667880
rect 119840 667640 120080 667880
rect 120190 667640 120430 667880
rect 120520 667640 120760 667880
rect 120850 667640 121090 667880
rect 121180 667640 121420 667880
rect 121530 667640 121770 667880
rect 110810 667290 111050 667530
rect 111140 667290 111380 667530
rect 111470 667290 111710 667530
rect 111800 667290 112040 667530
rect 112150 667290 112390 667530
rect 112480 667290 112720 667530
rect 112810 667290 113050 667530
rect 113140 667290 113380 667530
rect 113490 667290 113730 667530
rect 113820 667290 114060 667530
rect 114150 667290 114390 667530
rect 114480 667290 114720 667530
rect 114830 667290 115070 667530
rect 115160 667290 115400 667530
rect 115490 667290 115730 667530
rect 115820 667290 116060 667530
rect 116170 667290 116410 667530
rect 116500 667290 116740 667530
rect 116830 667290 117070 667530
rect 117160 667290 117400 667530
rect 117510 667290 117750 667530
rect 117840 667290 118080 667530
rect 118170 667290 118410 667530
rect 118500 667290 118740 667530
rect 118850 667290 119090 667530
rect 119180 667290 119420 667530
rect 119510 667290 119750 667530
rect 119840 667290 120080 667530
rect 120190 667290 120430 667530
rect 120520 667290 120760 667530
rect 120850 667290 121090 667530
rect 121180 667290 121420 667530
rect 121530 667290 121770 667530
rect 110810 666960 111050 667200
rect 111140 666960 111380 667200
rect 111470 666960 111710 667200
rect 111800 666960 112040 667200
rect 112150 666960 112390 667200
rect 112480 666960 112720 667200
rect 112810 666960 113050 667200
rect 113140 666960 113380 667200
rect 113490 666960 113730 667200
rect 113820 666960 114060 667200
rect 114150 666960 114390 667200
rect 114480 666960 114720 667200
rect 114830 666960 115070 667200
rect 115160 666960 115400 667200
rect 115490 666960 115730 667200
rect 115820 666960 116060 667200
rect 116170 666960 116410 667200
rect 116500 666960 116740 667200
rect 116830 666960 117070 667200
rect 117160 666960 117400 667200
rect 117510 666960 117750 667200
rect 117840 666960 118080 667200
rect 118170 666960 118410 667200
rect 118500 666960 118740 667200
rect 118850 666960 119090 667200
rect 119180 666960 119420 667200
rect 119510 666960 119750 667200
rect 119840 666960 120080 667200
rect 120190 666960 120430 667200
rect 120520 666960 120760 667200
rect 120850 666960 121090 667200
rect 121180 666960 121420 667200
rect 121530 666960 121770 667200
rect 110810 666630 111050 666870
rect 111140 666630 111380 666870
rect 111470 666630 111710 666870
rect 111800 666630 112040 666870
rect 112150 666630 112390 666870
rect 112480 666630 112720 666870
rect 112810 666630 113050 666870
rect 113140 666630 113380 666870
rect 113490 666630 113730 666870
rect 113820 666630 114060 666870
rect 114150 666630 114390 666870
rect 114480 666630 114720 666870
rect 114830 666630 115070 666870
rect 115160 666630 115400 666870
rect 115490 666630 115730 666870
rect 115820 666630 116060 666870
rect 116170 666630 116410 666870
rect 116500 666630 116740 666870
rect 116830 666630 117070 666870
rect 117160 666630 117400 666870
rect 117510 666630 117750 666870
rect 117840 666630 118080 666870
rect 118170 666630 118410 666870
rect 118500 666630 118740 666870
rect 118850 666630 119090 666870
rect 119180 666630 119420 666870
rect 119510 666630 119750 666870
rect 119840 666630 120080 666870
rect 120190 666630 120430 666870
rect 120520 666630 120760 666870
rect 120850 666630 121090 666870
rect 121180 666630 121420 666870
rect 121530 666630 121770 666870
rect 110810 666300 111050 666540
rect 111140 666300 111380 666540
rect 111470 666300 111710 666540
rect 111800 666300 112040 666540
rect 112150 666300 112390 666540
rect 112480 666300 112720 666540
rect 112810 666300 113050 666540
rect 113140 666300 113380 666540
rect 113490 666300 113730 666540
rect 113820 666300 114060 666540
rect 114150 666300 114390 666540
rect 114480 666300 114720 666540
rect 114830 666300 115070 666540
rect 115160 666300 115400 666540
rect 115490 666300 115730 666540
rect 115820 666300 116060 666540
rect 116170 666300 116410 666540
rect 116500 666300 116740 666540
rect 116830 666300 117070 666540
rect 117160 666300 117400 666540
rect 117510 666300 117750 666540
rect 117840 666300 118080 666540
rect 118170 666300 118410 666540
rect 118500 666300 118740 666540
rect 118850 666300 119090 666540
rect 119180 666300 119420 666540
rect 119510 666300 119750 666540
rect 119840 666300 120080 666540
rect 120190 666300 120430 666540
rect 120520 666300 120760 666540
rect 120850 666300 121090 666540
rect 121180 666300 121420 666540
rect 121530 666300 121770 666540
rect 110810 665950 111050 666190
rect 111140 665950 111380 666190
rect 111470 665950 111710 666190
rect 111800 665950 112040 666190
rect 112150 665950 112390 666190
rect 112480 665950 112720 666190
rect 112810 665950 113050 666190
rect 113140 665950 113380 666190
rect 113490 665950 113730 666190
rect 113820 665950 114060 666190
rect 114150 665950 114390 666190
rect 114480 665950 114720 666190
rect 114830 665950 115070 666190
rect 115160 665950 115400 666190
rect 115490 665950 115730 666190
rect 115820 665950 116060 666190
rect 116170 665950 116410 666190
rect 116500 665950 116740 666190
rect 116830 665950 117070 666190
rect 117160 665950 117400 666190
rect 117510 665950 117750 666190
rect 117840 665950 118080 666190
rect 118170 665950 118410 666190
rect 118500 665950 118740 666190
rect 118850 665950 119090 666190
rect 119180 665950 119420 666190
rect 119510 665950 119750 666190
rect 119840 665950 120080 666190
rect 120190 665950 120430 666190
rect 120520 665950 120760 666190
rect 120850 665950 121090 666190
rect 121180 665950 121420 666190
rect 121530 665950 121770 666190
rect 110810 665620 111050 665860
rect 111140 665620 111380 665860
rect 111470 665620 111710 665860
rect 111800 665620 112040 665860
rect 112150 665620 112390 665860
rect 112480 665620 112720 665860
rect 112810 665620 113050 665860
rect 113140 665620 113380 665860
rect 113490 665620 113730 665860
rect 113820 665620 114060 665860
rect 114150 665620 114390 665860
rect 114480 665620 114720 665860
rect 114830 665620 115070 665860
rect 115160 665620 115400 665860
rect 115490 665620 115730 665860
rect 115820 665620 116060 665860
rect 116170 665620 116410 665860
rect 116500 665620 116740 665860
rect 116830 665620 117070 665860
rect 117160 665620 117400 665860
rect 117510 665620 117750 665860
rect 117840 665620 118080 665860
rect 118170 665620 118410 665860
rect 118500 665620 118740 665860
rect 118850 665620 119090 665860
rect 119180 665620 119420 665860
rect 119510 665620 119750 665860
rect 119840 665620 120080 665860
rect 120190 665620 120430 665860
rect 120520 665620 120760 665860
rect 120850 665620 121090 665860
rect 121180 665620 121420 665860
rect 121530 665620 121770 665860
rect 110810 665290 111050 665530
rect 111140 665290 111380 665530
rect 111470 665290 111710 665530
rect 111800 665290 112040 665530
rect 112150 665290 112390 665530
rect 112480 665290 112720 665530
rect 112810 665290 113050 665530
rect 113140 665290 113380 665530
rect 113490 665290 113730 665530
rect 113820 665290 114060 665530
rect 114150 665290 114390 665530
rect 114480 665290 114720 665530
rect 114830 665290 115070 665530
rect 115160 665290 115400 665530
rect 115490 665290 115730 665530
rect 115820 665290 116060 665530
rect 116170 665290 116410 665530
rect 116500 665290 116740 665530
rect 116830 665290 117070 665530
rect 117160 665290 117400 665530
rect 117510 665290 117750 665530
rect 117840 665290 118080 665530
rect 118170 665290 118410 665530
rect 118500 665290 118740 665530
rect 118850 665290 119090 665530
rect 119180 665290 119420 665530
rect 119510 665290 119750 665530
rect 119840 665290 120080 665530
rect 120190 665290 120430 665530
rect 120520 665290 120760 665530
rect 120850 665290 121090 665530
rect 121180 665290 121420 665530
rect 121530 665290 121770 665530
rect 110810 664960 111050 665200
rect 111140 664960 111380 665200
rect 111470 664960 111710 665200
rect 111800 664960 112040 665200
rect 112150 664960 112390 665200
rect 112480 664960 112720 665200
rect 112810 664960 113050 665200
rect 113140 664960 113380 665200
rect 113490 664960 113730 665200
rect 113820 664960 114060 665200
rect 114150 664960 114390 665200
rect 114480 664960 114720 665200
rect 114830 664960 115070 665200
rect 115160 664960 115400 665200
rect 115490 664960 115730 665200
rect 115820 664960 116060 665200
rect 116170 664960 116410 665200
rect 116500 664960 116740 665200
rect 116830 664960 117070 665200
rect 117160 664960 117400 665200
rect 117510 664960 117750 665200
rect 117840 664960 118080 665200
rect 118170 664960 118410 665200
rect 118500 664960 118740 665200
rect 118850 664960 119090 665200
rect 119180 664960 119420 665200
rect 119510 664960 119750 665200
rect 119840 664960 120080 665200
rect 120190 664960 120430 665200
rect 120520 664960 120760 665200
rect 120850 664960 121090 665200
rect 121180 664960 121420 665200
rect 121530 664960 121770 665200
rect 110810 664610 111050 664850
rect 111140 664610 111380 664850
rect 111470 664610 111710 664850
rect 111800 664610 112040 664850
rect 112150 664610 112390 664850
rect 112480 664610 112720 664850
rect 112810 664610 113050 664850
rect 113140 664610 113380 664850
rect 113490 664610 113730 664850
rect 113820 664610 114060 664850
rect 114150 664610 114390 664850
rect 114480 664610 114720 664850
rect 114830 664610 115070 664850
rect 115160 664610 115400 664850
rect 115490 664610 115730 664850
rect 115820 664610 116060 664850
rect 116170 664610 116410 664850
rect 116500 664610 116740 664850
rect 116830 664610 117070 664850
rect 117160 664610 117400 664850
rect 117510 664610 117750 664850
rect 117840 664610 118080 664850
rect 118170 664610 118410 664850
rect 118500 664610 118740 664850
rect 118850 664610 119090 664850
rect 119180 664610 119420 664850
rect 119510 664610 119750 664850
rect 119840 664610 120080 664850
rect 120190 664610 120430 664850
rect 120520 664610 120760 664850
rect 120850 664610 121090 664850
rect 121180 664610 121420 664850
rect 121530 664610 121770 664850
rect 110810 664280 111050 664520
rect 111140 664280 111380 664520
rect 111470 664280 111710 664520
rect 111800 664280 112040 664520
rect 112150 664280 112390 664520
rect 112480 664280 112720 664520
rect 112810 664280 113050 664520
rect 113140 664280 113380 664520
rect 113490 664280 113730 664520
rect 113820 664280 114060 664520
rect 114150 664280 114390 664520
rect 114480 664280 114720 664520
rect 114830 664280 115070 664520
rect 115160 664280 115400 664520
rect 115490 664280 115730 664520
rect 115820 664280 116060 664520
rect 116170 664280 116410 664520
rect 116500 664280 116740 664520
rect 116830 664280 117070 664520
rect 117160 664280 117400 664520
rect 117510 664280 117750 664520
rect 117840 664280 118080 664520
rect 118170 664280 118410 664520
rect 118500 664280 118740 664520
rect 118850 664280 119090 664520
rect 119180 664280 119420 664520
rect 119510 664280 119750 664520
rect 119840 664280 120080 664520
rect 120190 664280 120430 664520
rect 120520 664280 120760 664520
rect 120850 664280 121090 664520
rect 121180 664280 121420 664520
rect 121530 664280 121770 664520
rect 110810 663950 111050 664190
rect 111140 663950 111380 664190
rect 111470 663950 111710 664190
rect 111800 663950 112040 664190
rect 112150 663950 112390 664190
rect 112480 663950 112720 664190
rect 112810 663950 113050 664190
rect 113140 663950 113380 664190
rect 113490 663950 113730 664190
rect 113820 663950 114060 664190
rect 114150 663950 114390 664190
rect 114480 663950 114720 664190
rect 114830 663950 115070 664190
rect 115160 663950 115400 664190
rect 115490 663950 115730 664190
rect 115820 663950 116060 664190
rect 116170 663950 116410 664190
rect 116500 663950 116740 664190
rect 116830 663950 117070 664190
rect 117160 663950 117400 664190
rect 117510 663950 117750 664190
rect 117840 663950 118080 664190
rect 118170 663950 118410 664190
rect 118500 663950 118740 664190
rect 118850 663950 119090 664190
rect 119180 663950 119420 664190
rect 119510 663950 119750 664190
rect 119840 663950 120080 664190
rect 120190 663950 120430 664190
rect 120520 663950 120760 664190
rect 120850 663950 121090 664190
rect 121180 663950 121420 664190
rect 121530 663950 121770 664190
rect 110810 663620 111050 663860
rect 111140 663620 111380 663860
rect 111470 663620 111710 663860
rect 111800 663620 112040 663860
rect 112150 663620 112390 663860
rect 112480 663620 112720 663860
rect 112810 663620 113050 663860
rect 113140 663620 113380 663860
rect 113490 663620 113730 663860
rect 113820 663620 114060 663860
rect 114150 663620 114390 663860
rect 114480 663620 114720 663860
rect 114830 663620 115070 663860
rect 115160 663620 115400 663860
rect 115490 663620 115730 663860
rect 115820 663620 116060 663860
rect 116170 663620 116410 663860
rect 116500 663620 116740 663860
rect 116830 663620 117070 663860
rect 117160 663620 117400 663860
rect 117510 663620 117750 663860
rect 117840 663620 118080 663860
rect 118170 663620 118410 663860
rect 118500 663620 118740 663860
rect 118850 663620 119090 663860
rect 119180 663620 119420 663860
rect 119510 663620 119750 663860
rect 119840 663620 120080 663860
rect 120190 663620 120430 663860
rect 120520 663620 120760 663860
rect 120850 663620 121090 663860
rect 121180 663620 121420 663860
rect 121530 663620 121770 663860
rect 110810 663270 111050 663510
rect 111140 663270 111380 663510
rect 111470 663270 111710 663510
rect 111800 663270 112040 663510
rect 112150 663270 112390 663510
rect 112480 663270 112720 663510
rect 112810 663270 113050 663510
rect 113140 663270 113380 663510
rect 113490 663270 113730 663510
rect 113820 663270 114060 663510
rect 114150 663270 114390 663510
rect 114480 663270 114720 663510
rect 114830 663270 115070 663510
rect 115160 663270 115400 663510
rect 115490 663270 115730 663510
rect 115820 663270 116060 663510
rect 116170 663270 116410 663510
rect 116500 663270 116740 663510
rect 116830 663270 117070 663510
rect 117160 663270 117400 663510
rect 117510 663270 117750 663510
rect 117840 663270 118080 663510
rect 118170 663270 118410 663510
rect 118500 663270 118740 663510
rect 118850 663270 119090 663510
rect 119180 663270 119420 663510
rect 119510 663270 119750 663510
rect 119840 663270 120080 663510
rect 120190 663270 120430 663510
rect 120520 663270 120760 663510
rect 120850 663270 121090 663510
rect 121180 663270 121420 663510
rect 121530 663270 121770 663510
rect 110810 662940 111050 663180
rect 111140 662940 111380 663180
rect 111470 662940 111710 663180
rect 111800 662940 112040 663180
rect 112150 662940 112390 663180
rect 112480 662940 112720 663180
rect 112810 662940 113050 663180
rect 113140 662940 113380 663180
rect 113490 662940 113730 663180
rect 113820 662940 114060 663180
rect 114150 662940 114390 663180
rect 114480 662940 114720 663180
rect 114830 662940 115070 663180
rect 115160 662940 115400 663180
rect 115490 662940 115730 663180
rect 115820 662940 116060 663180
rect 116170 662940 116410 663180
rect 116500 662940 116740 663180
rect 116830 662940 117070 663180
rect 117160 662940 117400 663180
rect 117510 662940 117750 663180
rect 117840 662940 118080 663180
rect 118170 662940 118410 663180
rect 118500 662940 118740 663180
rect 118850 662940 119090 663180
rect 119180 662940 119420 663180
rect 119510 662940 119750 663180
rect 119840 662940 120080 663180
rect 120190 662940 120430 663180
rect 120520 662940 120760 663180
rect 120850 662940 121090 663180
rect 121180 662940 121420 663180
rect 121530 662940 121770 663180
rect 110810 662610 111050 662850
rect 111140 662610 111380 662850
rect 111470 662610 111710 662850
rect 111800 662610 112040 662850
rect 112150 662610 112390 662850
rect 112480 662610 112720 662850
rect 112810 662610 113050 662850
rect 113140 662610 113380 662850
rect 113490 662610 113730 662850
rect 113820 662610 114060 662850
rect 114150 662610 114390 662850
rect 114480 662610 114720 662850
rect 114830 662610 115070 662850
rect 115160 662610 115400 662850
rect 115490 662610 115730 662850
rect 115820 662610 116060 662850
rect 116170 662610 116410 662850
rect 116500 662610 116740 662850
rect 116830 662610 117070 662850
rect 117160 662610 117400 662850
rect 117510 662610 117750 662850
rect 117840 662610 118080 662850
rect 118170 662610 118410 662850
rect 118500 662610 118740 662850
rect 118850 662610 119090 662850
rect 119180 662610 119420 662850
rect 119510 662610 119750 662850
rect 119840 662610 120080 662850
rect 120190 662610 120430 662850
rect 120520 662610 120760 662850
rect 120850 662610 121090 662850
rect 121180 662610 121420 662850
rect 121530 662610 121770 662850
rect 110810 662280 111050 662520
rect 111140 662280 111380 662520
rect 111470 662280 111710 662520
rect 111800 662280 112040 662520
rect 112150 662280 112390 662520
rect 112480 662280 112720 662520
rect 112810 662280 113050 662520
rect 113140 662280 113380 662520
rect 113490 662280 113730 662520
rect 113820 662280 114060 662520
rect 114150 662280 114390 662520
rect 114480 662280 114720 662520
rect 114830 662280 115070 662520
rect 115160 662280 115400 662520
rect 115490 662280 115730 662520
rect 115820 662280 116060 662520
rect 116170 662280 116410 662520
rect 116500 662280 116740 662520
rect 116830 662280 117070 662520
rect 117160 662280 117400 662520
rect 117510 662280 117750 662520
rect 117840 662280 118080 662520
rect 118170 662280 118410 662520
rect 118500 662280 118740 662520
rect 118850 662280 119090 662520
rect 119180 662280 119420 662520
rect 119510 662280 119750 662520
rect 119840 662280 120080 662520
rect 120190 662280 120430 662520
rect 120520 662280 120760 662520
rect 120850 662280 121090 662520
rect 121180 662280 121420 662520
rect 121530 662280 121770 662520
rect 110810 661930 111050 662170
rect 111140 661930 111380 662170
rect 111470 661930 111710 662170
rect 111800 661930 112040 662170
rect 112150 661930 112390 662170
rect 112480 661930 112720 662170
rect 112810 661930 113050 662170
rect 113140 661930 113380 662170
rect 113490 661930 113730 662170
rect 113820 661930 114060 662170
rect 114150 661930 114390 662170
rect 114480 661930 114720 662170
rect 114830 661930 115070 662170
rect 115160 661930 115400 662170
rect 115490 661930 115730 662170
rect 115820 661930 116060 662170
rect 116170 661930 116410 662170
rect 116500 661930 116740 662170
rect 116830 661930 117070 662170
rect 117160 661930 117400 662170
rect 117510 661930 117750 662170
rect 117840 661930 118080 662170
rect 118170 661930 118410 662170
rect 118500 661930 118740 662170
rect 118850 661930 119090 662170
rect 119180 661930 119420 662170
rect 119510 661930 119750 662170
rect 119840 661930 120080 662170
rect 120190 661930 120430 662170
rect 120520 661930 120760 662170
rect 120850 661930 121090 662170
rect 121180 661930 121420 662170
rect 121530 661930 121770 662170
rect 110810 661600 111050 661840
rect 111140 661600 111380 661840
rect 111470 661600 111710 661840
rect 111800 661600 112040 661840
rect 112150 661600 112390 661840
rect 112480 661600 112720 661840
rect 112810 661600 113050 661840
rect 113140 661600 113380 661840
rect 113490 661600 113730 661840
rect 113820 661600 114060 661840
rect 114150 661600 114390 661840
rect 114480 661600 114720 661840
rect 114830 661600 115070 661840
rect 115160 661600 115400 661840
rect 115490 661600 115730 661840
rect 115820 661600 116060 661840
rect 116170 661600 116410 661840
rect 116500 661600 116740 661840
rect 116830 661600 117070 661840
rect 117160 661600 117400 661840
rect 117510 661600 117750 661840
rect 117840 661600 118080 661840
rect 118170 661600 118410 661840
rect 118500 661600 118740 661840
rect 118850 661600 119090 661840
rect 119180 661600 119420 661840
rect 119510 661600 119750 661840
rect 119840 661600 120080 661840
rect 120190 661600 120430 661840
rect 120520 661600 120760 661840
rect 120850 661600 121090 661840
rect 121180 661600 121420 661840
rect 121530 661600 121770 661840
rect 110810 661270 111050 661510
rect 111140 661270 111380 661510
rect 111470 661270 111710 661510
rect 111800 661270 112040 661510
rect 112150 661270 112390 661510
rect 112480 661270 112720 661510
rect 112810 661270 113050 661510
rect 113140 661270 113380 661510
rect 113490 661270 113730 661510
rect 113820 661270 114060 661510
rect 114150 661270 114390 661510
rect 114480 661270 114720 661510
rect 114830 661270 115070 661510
rect 115160 661270 115400 661510
rect 115490 661270 115730 661510
rect 115820 661270 116060 661510
rect 116170 661270 116410 661510
rect 116500 661270 116740 661510
rect 116830 661270 117070 661510
rect 117160 661270 117400 661510
rect 117510 661270 117750 661510
rect 117840 661270 118080 661510
rect 118170 661270 118410 661510
rect 118500 661270 118740 661510
rect 118850 661270 119090 661510
rect 119180 661270 119420 661510
rect 119510 661270 119750 661510
rect 119840 661270 120080 661510
rect 120190 661270 120430 661510
rect 120520 661270 120760 661510
rect 120850 661270 121090 661510
rect 121180 661270 121420 661510
rect 121530 661270 121770 661510
rect 110810 660940 111050 661180
rect 111140 660940 111380 661180
rect 111470 660940 111710 661180
rect 111800 660940 112040 661180
rect 112150 660940 112390 661180
rect 112480 660940 112720 661180
rect 112810 660940 113050 661180
rect 113140 660940 113380 661180
rect 113490 660940 113730 661180
rect 113820 660940 114060 661180
rect 114150 660940 114390 661180
rect 114480 660940 114720 661180
rect 114830 660940 115070 661180
rect 115160 660940 115400 661180
rect 115490 660940 115730 661180
rect 115820 660940 116060 661180
rect 116170 660940 116410 661180
rect 116500 660940 116740 661180
rect 116830 660940 117070 661180
rect 117160 660940 117400 661180
rect 117510 660940 117750 661180
rect 117840 660940 118080 661180
rect 118170 660940 118410 661180
rect 118500 660940 118740 661180
rect 118850 660940 119090 661180
rect 119180 660940 119420 661180
rect 119510 660940 119750 661180
rect 119840 660940 120080 661180
rect 120190 660940 120430 661180
rect 120520 660940 120760 661180
rect 120850 660940 121090 661180
rect 121180 660940 121420 661180
rect 121530 660940 121770 661180
rect 122190 671660 122430 671900
rect 122520 671660 122760 671900
rect 122850 671660 123090 671900
rect 123180 671660 123420 671900
rect 123530 671660 123770 671900
rect 123860 671660 124100 671900
rect 124190 671660 124430 671900
rect 124520 671660 124760 671900
rect 124870 671660 125110 671900
rect 125200 671660 125440 671900
rect 125530 671660 125770 671900
rect 125860 671660 126100 671900
rect 126210 671660 126450 671900
rect 126540 671660 126780 671900
rect 126870 671660 127110 671900
rect 127200 671660 127440 671900
rect 127550 671660 127790 671900
rect 127880 671660 128120 671900
rect 128210 671660 128450 671900
rect 128540 671660 128780 671900
rect 128890 671660 129130 671900
rect 129220 671660 129460 671900
rect 129550 671660 129790 671900
rect 129880 671660 130120 671900
rect 130230 671660 130470 671900
rect 130560 671660 130800 671900
rect 130890 671660 131130 671900
rect 131220 671660 131460 671900
rect 131570 671660 131810 671900
rect 131900 671660 132140 671900
rect 132230 671660 132470 671900
rect 132560 671660 132800 671900
rect 132910 671660 133150 671900
rect 122190 671310 122430 671550
rect 122520 671310 122760 671550
rect 122850 671310 123090 671550
rect 123180 671310 123420 671550
rect 123530 671310 123770 671550
rect 123860 671310 124100 671550
rect 124190 671310 124430 671550
rect 124520 671310 124760 671550
rect 124870 671310 125110 671550
rect 125200 671310 125440 671550
rect 125530 671310 125770 671550
rect 125860 671310 126100 671550
rect 126210 671310 126450 671550
rect 126540 671310 126780 671550
rect 126870 671310 127110 671550
rect 127200 671310 127440 671550
rect 127550 671310 127790 671550
rect 127880 671310 128120 671550
rect 128210 671310 128450 671550
rect 128540 671310 128780 671550
rect 128890 671310 129130 671550
rect 129220 671310 129460 671550
rect 129550 671310 129790 671550
rect 129880 671310 130120 671550
rect 130230 671310 130470 671550
rect 130560 671310 130800 671550
rect 130890 671310 131130 671550
rect 131220 671310 131460 671550
rect 131570 671310 131810 671550
rect 131900 671310 132140 671550
rect 132230 671310 132470 671550
rect 132560 671310 132800 671550
rect 132910 671310 133150 671550
rect 122190 670980 122430 671220
rect 122520 670980 122760 671220
rect 122850 670980 123090 671220
rect 123180 670980 123420 671220
rect 123530 670980 123770 671220
rect 123860 670980 124100 671220
rect 124190 670980 124430 671220
rect 124520 670980 124760 671220
rect 124870 670980 125110 671220
rect 125200 670980 125440 671220
rect 125530 670980 125770 671220
rect 125860 670980 126100 671220
rect 126210 670980 126450 671220
rect 126540 670980 126780 671220
rect 126870 670980 127110 671220
rect 127200 670980 127440 671220
rect 127550 670980 127790 671220
rect 127880 670980 128120 671220
rect 128210 670980 128450 671220
rect 128540 670980 128780 671220
rect 128890 670980 129130 671220
rect 129220 670980 129460 671220
rect 129550 670980 129790 671220
rect 129880 670980 130120 671220
rect 130230 670980 130470 671220
rect 130560 670980 130800 671220
rect 130890 670980 131130 671220
rect 131220 670980 131460 671220
rect 131570 670980 131810 671220
rect 131900 670980 132140 671220
rect 132230 670980 132470 671220
rect 132560 670980 132800 671220
rect 132910 670980 133150 671220
rect 122190 670650 122430 670890
rect 122520 670650 122760 670890
rect 122850 670650 123090 670890
rect 123180 670650 123420 670890
rect 123530 670650 123770 670890
rect 123860 670650 124100 670890
rect 124190 670650 124430 670890
rect 124520 670650 124760 670890
rect 124870 670650 125110 670890
rect 125200 670650 125440 670890
rect 125530 670650 125770 670890
rect 125860 670650 126100 670890
rect 126210 670650 126450 670890
rect 126540 670650 126780 670890
rect 126870 670650 127110 670890
rect 127200 670650 127440 670890
rect 127550 670650 127790 670890
rect 127880 670650 128120 670890
rect 128210 670650 128450 670890
rect 128540 670650 128780 670890
rect 128890 670650 129130 670890
rect 129220 670650 129460 670890
rect 129550 670650 129790 670890
rect 129880 670650 130120 670890
rect 130230 670650 130470 670890
rect 130560 670650 130800 670890
rect 130890 670650 131130 670890
rect 131220 670650 131460 670890
rect 131570 670650 131810 670890
rect 131900 670650 132140 670890
rect 132230 670650 132470 670890
rect 132560 670650 132800 670890
rect 132910 670650 133150 670890
rect 122190 670320 122430 670560
rect 122520 670320 122760 670560
rect 122850 670320 123090 670560
rect 123180 670320 123420 670560
rect 123530 670320 123770 670560
rect 123860 670320 124100 670560
rect 124190 670320 124430 670560
rect 124520 670320 124760 670560
rect 124870 670320 125110 670560
rect 125200 670320 125440 670560
rect 125530 670320 125770 670560
rect 125860 670320 126100 670560
rect 126210 670320 126450 670560
rect 126540 670320 126780 670560
rect 126870 670320 127110 670560
rect 127200 670320 127440 670560
rect 127550 670320 127790 670560
rect 127880 670320 128120 670560
rect 128210 670320 128450 670560
rect 128540 670320 128780 670560
rect 128890 670320 129130 670560
rect 129220 670320 129460 670560
rect 129550 670320 129790 670560
rect 129880 670320 130120 670560
rect 130230 670320 130470 670560
rect 130560 670320 130800 670560
rect 130890 670320 131130 670560
rect 131220 670320 131460 670560
rect 131570 670320 131810 670560
rect 131900 670320 132140 670560
rect 132230 670320 132470 670560
rect 132560 670320 132800 670560
rect 132910 670320 133150 670560
rect 122190 669970 122430 670210
rect 122520 669970 122760 670210
rect 122850 669970 123090 670210
rect 123180 669970 123420 670210
rect 123530 669970 123770 670210
rect 123860 669970 124100 670210
rect 124190 669970 124430 670210
rect 124520 669970 124760 670210
rect 124870 669970 125110 670210
rect 125200 669970 125440 670210
rect 125530 669970 125770 670210
rect 125860 669970 126100 670210
rect 126210 669970 126450 670210
rect 126540 669970 126780 670210
rect 126870 669970 127110 670210
rect 127200 669970 127440 670210
rect 127550 669970 127790 670210
rect 127880 669970 128120 670210
rect 128210 669970 128450 670210
rect 128540 669970 128780 670210
rect 128890 669970 129130 670210
rect 129220 669970 129460 670210
rect 129550 669970 129790 670210
rect 129880 669970 130120 670210
rect 130230 669970 130470 670210
rect 130560 669970 130800 670210
rect 130890 669970 131130 670210
rect 131220 669970 131460 670210
rect 131570 669970 131810 670210
rect 131900 669970 132140 670210
rect 132230 669970 132470 670210
rect 132560 669970 132800 670210
rect 132910 669970 133150 670210
rect 122190 669640 122430 669880
rect 122520 669640 122760 669880
rect 122850 669640 123090 669880
rect 123180 669640 123420 669880
rect 123530 669640 123770 669880
rect 123860 669640 124100 669880
rect 124190 669640 124430 669880
rect 124520 669640 124760 669880
rect 124870 669640 125110 669880
rect 125200 669640 125440 669880
rect 125530 669640 125770 669880
rect 125860 669640 126100 669880
rect 126210 669640 126450 669880
rect 126540 669640 126780 669880
rect 126870 669640 127110 669880
rect 127200 669640 127440 669880
rect 127550 669640 127790 669880
rect 127880 669640 128120 669880
rect 128210 669640 128450 669880
rect 128540 669640 128780 669880
rect 128890 669640 129130 669880
rect 129220 669640 129460 669880
rect 129550 669640 129790 669880
rect 129880 669640 130120 669880
rect 130230 669640 130470 669880
rect 130560 669640 130800 669880
rect 130890 669640 131130 669880
rect 131220 669640 131460 669880
rect 131570 669640 131810 669880
rect 131900 669640 132140 669880
rect 132230 669640 132470 669880
rect 132560 669640 132800 669880
rect 132910 669640 133150 669880
rect 122190 669310 122430 669550
rect 122520 669310 122760 669550
rect 122850 669310 123090 669550
rect 123180 669310 123420 669550
rect 123530 669310 123770 669550
rect 123860 669310 124100 669550
rect 124190 669310 124430 669550
rect 124520 669310 124760 669550
rect 124870 669310 125110 669550
rect 125200 669310 125440 669550
rect 125530 669310 125770 669550
rect 125860 669310 126100 669550
rect 126210 669310 126450 669550
rect 126540 669310 126780 669550
rect 126870 669310 127110 669550
rect 127200 669310 127440 669550
rect 127550 669310 127790 669550
rect 127880 669310 128120 669550
rect 128210 669310 128450 669550
rect 128540 669310 128780 669550
rect 128890 669310 129130 669550
rect 129220 669310 129460 669550
rect 129550 669310 129790 669550
rect 129880 669310 130120 669550
rect 130230 669310 130470 669550
rect 130560 669310 130800 669550
rect 130890 669310 131130 669550
rect 131220 669310 131460 669550
rect 131570 669310 131810 669550
rect 131900 669310 132140 669550
rect 132230 669310 132470 669550
rect 132560 669310 132800 669550
rect 132910 669310 133150 669550
rect 122190 668980 122430 669220
rect 122520 668980 122760 669220
rect 122850 668980 123090 669220
rect 123180 668980 123420 669220
rect 123530 668980 123770 669220
rect 123860 668980 124100 669220
rect 124190 668980 124430 669220
rect 124520 668980 124760 669220
rect 124870 668980 125110 669220
rect 125200 668980 125440 669220
rect 125530 668980 125770 669220
rect 125860 668980 126100 669220
rect 126210 668980 126450 669220
rect 126540 668980 126780 669220
rect 126870 668980 127110 669220
rect 127200 668980 127440 669220
rect 127550 668980 127790 669220
rect 127880 668980 128120 669220
rect 128210 668980 128450 669220
rect 128540 668980 128780 669220
rect 128890 668980 129130 669220
rect 129220 668980 129460 669220
rect 129550 668980 129790 669220
rect 129880 668980 130120 669220
rect 130230 668980 130470 669220
rect 130560 668980 130800 669220
rect 130890 668980 131130 669220
rect 131220 668980 131460 669220
rect 131570 668980 131810 669220
rect 131900 668980 132140 669220
rect 132230 668980 132470 669220
rect 132560 668980 132800 669220
rect 132910 668980 133150 669220
rect 122190 668630 122430 668870
rect 122520 668630 122760 668870
rect 122850 668630 123090 668870
rect 123180 668630 123420 668870
rect 123530 668630 123770 668870
rect 123860 668630 124100 668870
rect 124190 668630 124430 668870
rect 124520 668630 124760 668870
rect 124870 668630 125110 668870
rect 125200 668630 125440 668870
rect 125530 668630 125770 668870
rect 125860 668630 126100 668870
rect 126210 668630 126450 668870
rect 126540 668630 126780 668870
rect 126870 668630 127110 668870
rect 127200 668630 127440 668870
rect 127550 668630 127790 668870
rect 127880 668630 128120 668870
rect 128210 668630 128450 668870
rect 128540 668630 128780 668870
rect 128890 668630 129130 668870
rect 129220 668630 129460 668870
rect 129550 668630 129790 668870
rect 129880 668630 130120 668870
rect 130230 668630 130470 668870
rect 130560 668630 130800 668870
rect 130890 668630 131130 668870
rect 131220 668630 131460 668870
rect 131570 668630 131810 668870
rect 131900 668630 132140 668870
rect 132230 668630 132470 668870
rect 132560 668630 132800 668870
rect 132910 668630 133150 668870
rect 122190 668300 122430 668540
rect 122520 668300 122760 668540
rect 122850 668300 123090 668540
rect 123180 668300 123420 668540
rect 123530 668300 123770 668540
rect 123860 668300 124100 668540
rect 124190 668300 124430 668540
rect 124520 668300 124760 668540
rect 124870 668300 125110 668540
rect 125200 668300 125440 668540
rect 125530 668300 125770 668540
rect 125860 668300 126100 668540
rect 126210 668300 126450 668540
rect 126540 668300 126780 668540
rect 126870 668300 127110 668540
rect 127200 668300 127440 668540
rect 127550 668300 127790 668540
rect 127880 668300 128120 668540
rect 128210 668300 128450 668540
rect 128540 668300 128780 668540
rect 128890 668300 129130 668540
rect 129220 668300 129460 668540
rect 129550 668300 129790 668540
rect 129880 668300 130120 668540
rect 130230 668300 130470 668540
rect 130560 668300 130800 668540
rect 130890 668300 131130 668540
rect 131220 668300 131460 668540
rect 131570 668300 131810 668540
rect 131900 668300 132140 668540
rect 132230 668300 132470 668540
rect 132560 668300 132800 668540
rect 132910 668300 133150 668540
rect 122190 667970 122430 668210
rect 122520 667970 122760 668210
rect 122850 667970 123090 668210
rect 123180 667970 123420 668210
rect 123530 667970 123770 668210
rect 123860 667970 124100 668210
rect 124190 667970 124430 668210
rect 124520 667970 124760 668210
rect 124870 667970 125110 668210
rect 125200 667970 125440 668210
rect 125530 667970 125770 668210
rect 125860 667970 126100 668210
rect 126210 667970 126450 668210
rect 126540 667970 126780 668210
rect 126870 667970 127110 668210
rect 127200 667970 127440 668210
rect 127550 667970 127790 668210
rect 127880 667970 128120 668210
rect 128210 667970 128450 668210
rect 128540 667970 128780 668210
rect 128890 667970 129130 668210
rect 129220 667970 129460 668210
rect 129550 667970 129790 668210
rect 129880 667970 130120 668210
rect 130230 667970 130470 668210
rect 130560 667970 130800 668210
rect 130890 667970 131130 668210
rect 131220 667970 131460 668210
rect 131570 667970 131810 668210
rect 131900 667970 132140 668210
rect 132230 667970 132470 668210
rect 132560 667970 132800 668210
rect 132910 667970 133150 668210
rect 122190 667640 122430 667880
rect 122520 667640 122760 667880
rect 122850 667640 123090 667880
rect 123180 667640 123420 667880
rect 123530 667640 123770 667880
rect 123860 667640 124100 667880
rect 124190 667640 124430 667880
rect 124520 667640 124760 667880
rect 124870 667640 125110 667880
rect 125200 667640 125440 667880
rect 125530 667640 125770 667880
rect 125860 667640 126100 667880
rect 126210 667640 126450 667880
rect 126540 667640 126780 667880
rect 126870 667640 127110 667880
rect 127200 667640 127440 667880
rect 127550 667640 127790 667880
rect 127880 667640 128120 667880
rect 128210 667640 128450 667880
rect 128540 667640 128780 667880
rect 128890 667640 129130 667880
rect 129220 667640 129460 667880
rect 129550 667640 129790 667880
rect 129880 667640 130120 667880
rect 130230 667640 130470 667880
rect 130560 667640 130800 667880
rect 130890 667640 131130 667880
rect 131220 667640 131460 667880
rect 131570 667640 131810 667880
rect 131900 667640 132140 667880
rect 132230 667640 132470 667880
rect 132560 667640 132800 667880
rect 132910 667640 133150 667880
rect 122190 667290 122430 667530
rect 122520 667290 122760 667530
rect 122850 667290 123090 667530
rect 123180 667290 123420 667530
rect 123530 667290 123770 667530
rect 123860 667290 124100 667530
rect 124190 667290 124430 667530
rect 124520 667290 124760 667530
rect 124870 667290 125110 667530
rect 125200 667290 125440 667530
rect 125530 667290 125770 667530
rect 125860 667290 126100 667530
rect 126210 667290 126450 667530
rect 126540 667290 126780 667530
rect 126870 667290 127110 667530
rect 127200 667290 127440 667530
rect 127550 667290 127790 667530
rect 127880 667290 128120 667530
rect 128210 667290 128450 667530
rect 128540 667290 128780 667530
rect 128890 667290 129130 667530
rect 129220 667290 129460 667530
rect 129550 667290 129790 667530
rect 129880 667290 130120 667530
rect 130230 667290 130470 667530
rect 130560 667290 130800 667530
rect 130890 667290 131130 667530
rect 131220 667290 131460 667530
rect 131570 667290 131810 667530
rect 131900 667290 132140 667530
rect 132230 667290 132470 667530
rect 132560 667290 132800 667530
rect 132910 667290 133150 667530
rect 122190 666960 122430 667200
rect 122520 666960 122760 667200
rect 122850 666960 123090 667200
rect 123180 666960 123420 667200
rect 123530 666960 123770 667200
rect 123860 666960 124100 667200
rect 124190 666960 124430 667200
rect 124520 666960 124760 667200
rect 124870 666960 125110 667200
rect 125200 666960 125440 667200
rect 125530 666960 125770 667200
rect 125860 666960 126100 667200
rect 126210 666960 126450 667200
rect 126540 666960 126780 667200
rect 126870 666960 127110 667200
rect 127200 666960 127440 667200
rect 127550 666960 127790 667200
rect 127880 666960 128120 667200
rect 128210 666960 128450 667200
rect 128540 666960 128780 667200
rect 128890 666960 129130 667200
rect 129220 666960 129460 667200
rect 129550 666960 129790 667200
rect 129880 666960 130120 667200
rect 130230 666960 130470 667200
rect 130560 666960 130800 667200
rect 130890 666960 131130 667200
rect 131220 666960 131460 667200
rect 131570 666960 131810 667200
rect 131900 666960 132140 667200
rect 132230 666960 132470 667200
rect 132560 666960 132800 667200
rect 132910 666960 133150 667200
rect 122190 666630 122430 666870
rect 122520 666630 122760 666870
rect 122850 666630 123090 666870
rect 123180 666630 123420 666870
rect 123530 666630 123770 666870
rect 123860 666630 124100 666870
rect 124190 666630 124430 666870
rect 124520 666630 124760 666870
rect 124870 666630 125110 666870
rect 125200 666630 125440 666870
rect 125530 666630 125770 666870
rect 125860 666630 126100 666870
rect 126210 666630 126450 666870
rect 126540 666630 126780 666870
rect 126870 666630 127110 666870
rect 127200 666630 127440 666870
rect 127550 666630 127790 666870
rect 127880 666630 128120 666870
rect 128210 666630 128450 666870
rect 128540 666630 128780 666870
rect 128890 666630 129130 666870
rect 129220 666630 129460 666870
rect 129550 666630 129790 666870
rect 129880 666630 130120 666870
rect 130230 666630 130470 666870
rect 130560 666630 130800 666870
rect 130890 666630 131130 666870
rect 131220 666630 131460 666870
rect 131570 666630 131810 666870
rect 131900 666630 132140 666870
rect 132230 666630 132470 666870
rect 132560 666630 132800 666870
rect 132910 666630 133150 666870
rect 122190 666300 122430 666540
rect 122520 666300 122760 666540
rect 122850 666300 123090 666540
rect 123180 666300 123420 666540
rect 123530 666300 123770 666540
rect 123860 666300 124100 666540
rect 124190 666300 124430 666540
rect 124520 666300 124760 666540
rect 124870 666300 125110 666540
rect 125200 666300 125440 666540
rect 125530 666300 125770 666540
rect 125860 666300 126100 666540
rect 126210 666300 126450 666540
rect 126540 666300 126780 666540
rect 126870 666300 127110 666540
rect 127200 666300 127440 666540
rect 127550 666300 127790 666540
rect 127880 666300 128120 666540
rect 128210 666300 128450 666540
rect 128540 666300 128780 666540
rect 128890 666300 129130 666540
rect 129220 666300 129460 666540
rect 129550 666300 129790 666540
rect 129880 666300 130120 666540
rect 130230 666300 130470 666540
rect 130560 666300 130800 666540
rect 130890 666300 131130 666540
rect 131220 666300 131460 666540
rect 131570 666300 131810 666540
rect 131900 666300 132140 666540
rect 132230 666300 132470 666540
rect 132560 666300 132800 666540
rect 132910 666300 133150 666540
rect 122190 665950 122430 666190
rect 122520 665950 122760 666190
rect 122850 665950 123090 666190
rect 123180 665950 123420 666190
rect 123530 665950 123770 666190
rect 123860 665950 124100 666190
rect 124190 665950 124430 666190
rect 124520 665950 124760 666190
rect 124870 665950 125110 666190
rect 125200 665950 125440 666190
rect 125530 665950 125770 666190
rect 125860 665950 126100 666190
rect 126210 665950 126450 666190
rect 126540 665950 126780 666190
rect 126870 665950 127110 666190
rect 127200 665950 127440 666190
rect 127550 665950 127790 666190
rect 127880 665950 128120 666190
rect 128210 665950 128450 666190
rect 128540 665950 128780 666190
rect 128890 665950 129130 666190
rect 129220 665950 129460 666190
rect 129550 665950 129790 666190
rect 129880 665950 130120 666190
rect 130230 665950 130470 666190
rect 130560 665950 130800 666190
rect 130890 665950 131130 666190
rect 131220 665950 131460 666190
rect 131570 665950 131810 666190
rect 131900 665950 132140 666190
rect 132230 665950 132470 666190
rect 132560 665950 132800 666190
rect 132910 665950 133150 666190
rect 122190 665620 122430 665860
rect 122520 665620 122760 665860
rect 122850 665620 123090 665860
rect 123180 665620 123420 665860
rect 123530 665620 123770 665860
rect 123860 665620 124100 665860
rect 124190 665620 124430 665860
rect 124520 665620 124760 665860
rect 124870 665620 125110 665860
rect 125200 665620 125440 665860
rect 125530 665620 125770 665860
rect 125860 665620 126100 665860
rect 126210 665620 126450 665860
rect 126540 665620 126780 665860
rect 126870 665620 127110 665860
rect 127200 665620 127440 665860
rect 127550 665620 127790 665860
rect 127880 665620 128120 665860
rect 128210 665620 128450 665860
rect 128540 665620 128780 665860
rect 128890 665620 129130 665860
rect 129220 665620 129460 665860
rect 129550 665620 129790 665860
rect 129880 665620 130120 665860
rect 130230 665620 130470 665860
rect 130560 665620 130800 665860
rect 130890 665620 131130 665860
rect 131220 665620 131460 665860
rect 131570 665620 131810 665860
rect 131900 665620 132140 665860
rect 132230 665620 132470 665860
rect 132560 665620 132800 665860
rect 132910 665620 133150 665860
rect 122190 665290 122430 665530
rect 122520 665290 122760 665530
rect 122850 665290 123090 665530
rect 123180 665290 123420 665530
rect 123530 665290 123770 665530
rect 123860 665290 124100 665530
rect 124190 665290 124430 665530
rect 124520 665290 124760 665530
rect 124870 665290 125110 665530
rect 125200 665290 125440 665530
rect 125530 665290 125770 665530
rect 125860 665290 126100 665530
rect 126210 665290 126450 665530
rect 126540 665290 126780 665530
rect 126870 665290 127110 665530
rect 127200 665290 127440 665530
rect 127550 665290 127790 665530
rect 127880 665290 128120 665530
rect 128210 665290 128450 665530
rect 128540 665290 128780 665530
rect 128890 665290 129130 665530
rect 129220 665290 129460 665530
rect 129550 665290 129790 665530
rect 129880 665290 130120 665530
rect 130230 665290 130470 665530
rect 130560 665290 130800 665530
rect 130890 665290 131130 665530
rect 131220 665290 131460 665530
rect 131570 665290 131810 665530
rect 131900 665290 132140 665530
rect 132230 665290 132470 665530
rect 132560 665290 132800 665530
rect 132910 665290 133150 665530
rect 122190 664960 122430 665200
rect 122520 664960 122760 665200
rect 122850 664960 123090 665200
rect 123180 664960 123420 665200
rect 123530 664960 123770 665200
rect 123860 664960 124100 665200
rect 124190 664960 124430 665200
rect 124520 664960 124760 665200
rect 124870 664960 125110 665200
rect 125200 664960 125440 665200
rect 125530 664960 125770 665200
rect 125860 664960 126100 665200
rect 126210 664960 126450 665200
rect 126540 664960 126780 665200
rect 126870 664960 127110 665200
rect 127200 664960 127440 665200
rect 127550 664960 127790 665200
rect 127880 664960 128120 665200
rect 128210 664960 128450 665200
rect 128540 664960 128780 665200
rect 128890 664960 129130 665200
rect 129220 664960 129460 665200
rect 129550 664960 129790 665200
rect 129880 664960 130120 665200
rect 130230 664960 130470 665200
rect 130560 664960 130800 665200
rect 130890 664960 131130 665200
rect 131220 664960 131460 665200
rect 131570 664960 131810 665200
rect 131900 664960 132140 665200
rect 132230 664960 132470 665200
rect 132560 664960 132800 665200
rect 132910 664960 133150 665200
rect 122190 664610 122430 664850
rect 122520 664610 122760 664850
rect 122850 664610 123090 664850
rect 123180 664610 123420 664850
rect 123530 664610 123770 664850
rect 123860 664610 124100 664850
rect 124190 664610 124430 664850
rect 124520 664610 124760 664850
rect 124870 664610 125110 664850
rect 125200 664610 125440 664850
rect 125530 664610 125770 664850
rect 125860 664610 126100 664850
rect 126210 664610 126450 664850
rect 126540 664610 126780 664850
rect 126870 664610 127110 664850
rect 127200 664610 127440 664850
rect 127550 664610 127790 664850
rect 127880 664610 128120 664850
rect 128210 664610 128450 664850
rect 128540 664610 128780 664850
rect 128890 664610 129130 664850
rect 129220 664610 129460 664850
rect 129550 664610 129790 664850
rect 129880 664610 130120 664850
rect 130230 664610 130470 664850
rect 130560 664610 130800 664850
rect 130890 664610 131130 664850
rect 131220 664610 131460 664850
rect 131570 664610 131810 664850
rect 131900 664610 132140 664850
rect 132230 664610 132470 664850
rect 132560 664610 132800 664850
rect 132910 664610 133150 664850
rect 122190 664280 122430 664520
rect 122520 664280 122760 664520
rect 122850 664280 123090 664520
rect 123180 664280 123420 664520
rect 123530 664280 123770 664520
rect 123860 664280 124100 664520
rect 124190 664280 124430 664520
rect 124520 664280 124760 664520
rect 124870 664280 125110 664520
rect 125200 664280 125440 664520
rect 125530 664280 125770 664520
rect 125860 664280 126100 664520
rect 126210 664280 126450 664520
rect 126540 664280 126780 664520
rect 126870 664280 127110 664520
rect 127200 664280 127440 664520
rect 127550 664280 127790 664520
rect 127880 664280 128120 664520
rect 128210 664280 128450 664520
rect 128540 664280 128780 664520
rect 128890 664280 129130 664520
rect 129220 664280 129460 664520
rect 129550 664280 129790 664520
rect 129880 664280 130120 664520
rect 130230 664280 130470 664520
rect 130560 664280 130800 664520
rect 130890 664280 131130 664520
rect 131220 664280 131460 664520
rect 131570 664280 131810 664520
rect 131900 664280 132140 664520
rect 132230 664280 132470 664520
rect 132560 664280 132800 664520
rect 132910 664280 133150 664520
rect 122190 663950 122430 664190
rect 122520 663950 122760 664190
rect 122850 663950 123090 664190
rect 123180 663950 123420 664190
rect 123530 663950 123770 664190
rect 123860 663950 124100 664190
rect 124190 663950 124430 664190
rect 124520 663950 124760 664190
rect 124870 663950 125110 664190
rect 125200 663950 125440 664190
rect 125530 663950 125770 664190
rect 125860 663950 126100 664190
rect 126210 663950 126450 664190
rect 126540 663950 126780 664190
rect 126870 663950 127110 664190
rect 127200 663950 127440 664190
rect 127550 663950 127790 664190
rect 127880 663950 128120 664190
rect 128210 663950 128450 664190
rect 128540 663950 128780 664190
rect 128890 663950 129130 664190
rect 129220 663950 129460 664190
rect 129550 663950 129790 664190
rect 129880 663950 130120 664190
rect 130230 663950 130470 664190
rect 130560 663950 130800 664190
rect 130890 663950 131130 664190
rect 131220 663950 131460 664190
rect 131570 663950 131810 664190
rect 131900 663950 132140 664190
rect 132230 663950 132470 664190
rect 132560 663950 132800 664190
rect 132910 663950 133150 664190
rect 122190 663620 122430 663860
rect 122520 663620 122760 663860
rect 122850 663620 123090 663860
rect 123180 663620 123420 663860
rect 123530 663620 123770 663860
rect 123860 663620 124100 663860
rect 124190 663620 124430 663860
rect 124520 663620 124760 663860
rect 124870 663620 125110 663860
rect 125200 663620 125440 663860
rect 125530 663620 125770 663860
rect 125860 663620 126100 663860
rect 126210 663620 126450 663860
rect 126540 663620 126780 663860
rect 126870 663620 127110 663860
rect 127200 663620 127440 663860
rect 127550 663620 127790 663860
rect 127880 663620 128120 663860
rect 128210 663620 128450 663860
rect 128540 663620 128780 663860
rect 128890 663620 129130 663860
rect 129220 663620 129460 663860
rect 129550 663620 129790 663860
rect 129880 663620 130120 663860
rect 130230 663620 130470 663860
rect 130560 663620 130800 663860
rect 130890 663620 131130 663860
rect 131220 663620 131460 663860
rect 131570 663620 131810 663860
rect 131900 663620 132140 663860
rect 132230 663620 132470 663860
rect 132560 663620 132800 663860
rect 132910 663620 133150 663860
rect 122190 663270 122430 663510
rect 122520 663270 122760 663510
rect 122850 663270 123090 663510
rect 123180 663270 123420 663510
rect 123530 663270 123770 663510
rect 123860 663270 124100 663510
rect 124190 663270 124430 663510
rect 124520 663270 124760 663510
rect 124870 663270 125110 663510
rect 125200 663270 125440 663510
rect 125530 663270 125770 663510
rect 125860 663270 126100 663510
rect 126210 663270 126450 663510
rect 126540 663270 126780 663510
rect 126870 663270 127110 663510
rect 127200 663270 127440 663510
rect 127550 663270 127790 663510
rect 127880 663270 128120 663510
rect 128210 663270 128450 663510
rect 128540 663270 128780 663510
rect 128890 663270 129130 663510
rect 129220 663270 129460 663510
rect 129550 663270 129790 663510
rect 129880 663270 130120 663510
rect 130230 663270 130470 663510
rect 130560 663270 130800 663510
rect 130890 663270 131130 663510
rect 131220 663270 131460 663510
rect 131570 663270 131810 663510
rect 131900 663270 132140 663510
rect 132230 663270 132470 663510
rect 132560 663270 132800 663510
rect 132910 663270 133150 663510
rect 122190 662940 122430 663180
rect 122520 662940 122760 663180
rect 122850 662940 123090 663180
rect 123180 662940 123420 663180
rect 123530 662940 123770 663180
rect 123860 662940 124100 663180
rect 124190 662940 124430 663180
rect 124520 662940 124760 663180
rect 124870 662940 125110 663180
rect 125200 662940 125440 663180
rect 125530 662940 125770 663180
rect 125860 662940 126100 663180
rect 126210 662940 126450 663180
rect 126540 662940 126780 663180
rect 126870 662940 127110 663180
rect 127200 662940 127440 663180
rect 127550 662940 127790 663180
rect 127880 662940 128120 663180
rect 128210 662940 128450 663180
rect 128540 662940 128780 663180
rect 128890 662940 129130 663180
rect 129220 662940 129460 663180
rect 129550 662940 129790 663180
rect 129880 662940 130120 663180
rect 130230 662940 130470 663180
rect 130560 662940 130800 663180
rect 130890 662940 131130 663180
rect 131220 662940 131460 663180
rect 131570 662940 131810 663180
rect 131900 662940 132140 663180
rect 132230 662940 132470 663180
rect 132560 662940 132800 663180
rect 132910 662940 133150 663180
rect 122190 662610 122430 662850
rect 122520 662610 122760 662850
rect 122850 662610 123090 662850
rect 123180 662610 123420 662850
rect 123530 662610 123770 662850
rect 123860 662610 124100 662850
rect 124190 662610 124430 662850
rect 124520 662610 124760 662850
rect 124870 662610 125110 662850
rect 125200 662610 125440 662850
rect 125530 662610 125770 662850
rect 125860 662610 126100 662850
rect 126210 662610 126450 662850
rect 126540 662610 126780 662850
rect 126870 662610 127110 662850
rect 127200 662610 127440 662850
rect 127550 662610 127790 662850
rect 127880 662610 128120 662850
rect 128210 662610 128450 662850
rect 128540 662610 128780 662850
rect 128890 662610 129130 662850
rect 129220 662610 129460 662850
rect 129550 662610 129790 662850
rect 129880 662610 130120 662850
rect 130230 662610 130470 662850
rect 130560 662610 130800 662850
rect 130890 662610 131130 662850
rect 131220 662610 131460 662850
rect 131570 662610 131810 662850
rect 131900 662610 132140 662850
rect 132230 662610 132470 662850
rect 132560 662610 132800 662850
rect 132910 662610 133150 662850
rect 122190 662280 122430 662520
rect 122520 662280 122760 662520
rect 122850 662280 123090 662520
rect 123180 662280 123420 662520
rect 123530 662280 123770 662520
rect 123860 662280 124100 662520
rect 124190 662280 124430 662520
rect 124520 662280 124760 662520
rect 124870 662280 125110 662520
rect 125200 662280 125440 662520
rect 125530 662280 125770 662520
rect 125860 662280 126100 662520
rect 126210 662280 126450 662520
rect 126540 662280 126780 662520
rect 126870 662280 127110 662520
rect 127200 662280 127440 662520
rect 127550 662280 127790 662520
rect 127880 662280 128120 662520
rect 128210 662280 128450 662520
rect 128540 662280 128780 662520
rect 128890 662280 129130 662520
rect 129220 662280 129460 662520
rect 129550 662280 129790 662520
rect 129880 662280 130120 662520
rect 130230 662280 130470 662520
rect 130560 662280 130800 662520
rect 130890 662280 131130 662520
rect 131220 662280 131460 662520
rect 131570 662280 131810 662520
rect 131900 662280 132140 662520
rect 132230 662280 132470 662520
rect 132560 662280 132800 662520
rect 132910 662280 133150 662520
rect 122190 661930 122430 662170
rect 122520 661930 122760 662170
rect 122850 661930 123090 662170
rect 123180 661930 123420 662170
rect 123530 661930 123770 662170
rect 123860 661930 124100 662170
rect 124190 661930 124430 662170
rect 124520 661930 124760 662170
rect 124870 661930 125110 662170
rect 125200 661930 125440 662170
rect 125530 661930 125770 662170
rect 125860 661930 126100 662170
rect 126210 661930 126450 662170
rect 126540 661930 126780 662170
rect 126870 661930 127110 662170
rect 127200 661930 127440 662170
rect 127550 661930 127790 662170
rect 127880 661930 128120 662170
rect 128210 661930 128450 662170
rect 128540 661930 128780 662170
rect 128890 661930 129130 662170
rect 129220 661930 129460 662170
rect 129550 661930 129790 662170
rect 129880 661930 130120 662170
rect 130230 661930 130470 662170
rect 130560 661930 130800 662170
rect 130890 661930 131130 662170
rect 131220 661930 131460 662170
rect 131570 661930 131810 662170
rect 131900 661930 132140 662170
rect 132230 661930 132470 662170
rect 132560 661930 132800 662170
rect 132910 661930 133150 662170
rect 122190 661600 122430 661840
rect 122520 661600 122760 661840
rect 122850 661600 123090 661840
rect 123180 661600 123420 661840
rect 123530 661600 123770 661840
rect 123860 661600 124100 661840
rect 124190 661600 124430 661840
rect 124520 661600 124760 661840
rect 124870 661600 125110 661840
rect 125200 661600 125440 661840
rect 125530 661600 125770 661840
rect 125860 661600 126100 661840
rect 126210 661600 126450 661840
rect 126540 661600 126780 661840
rect 126870 661600 127110 661840
rect 127200 661600 127440 661840
rect 127550 661600 127790 661840
rect 127880 661600 128120 661840
rect 128210 661600 128450 661840
rect 128540 661600 128780 661840
rect 128890 661600 129130 661840
rect 129220 661600 129460 661840
rect 129550 661600 129790 661840
rect 129880 661600 130120 661840
rect 130230 661600 130470 661840
rect 130560 661600 130800 661840
rect 130890 661600 131130 661840
rect 131220 661600 131460 661840
rect 131570 661600 131810 661840
rect 131900 661600 132140 661840
rect 132230 661600 132470 661840
rect 132560 661600 132800 661840
rect 132910 661600 133150 661840
rect 122190 661270 122430 661510
rect 122520 661270 122760 661510
rect 122850 661270 123090 661510
rect 123180 661270 123420 661510
rect 123530 661270 123770 661510
rect 123860 661270 124100 661510
rect 124190 661270 124430 661510
rect 124520 661270 124760 661510
rect 124870 661270 125110 661510
rect 125200 661270 125440 661510
rect 125530 661270 125770 661510
rect 125860 661270 126100 661510
rect 126210 661270 126450 661510
rect 126540 661270 126780 661510
rect 126870 661270 127110 661510
rect 127200 661270 127440 661510
rect 127550 661270 127790 661510
rect 127880 661270 128120 661510
rect 128210 661270 128450 661510
rect 128540 661270 128780 661510
rect 128890 661270 129130 661510
rect 129220 661270 129460 661510
rect 129550 661270 129790 661510
rect 129880 661270 130120 661510
rect 130230 661270 130470 661510
rect 130560 661270 130800 661510
rect 130890 661270 131130 661510
rect 131220 661270 131460 661510
rect 131570 661270 131810 661510
rect 131900 661270 132140 661510
rect 132230 661270 132470 661510
rect 132560 661270 132800 661510
rect 132910 661270 133150 661510
rect 122190 660940 122430 661180
rect 122520 660940 122760 661180
rect 122850 660940 123090 661180
rect 123180 660940 123420 661180
rect 123530 660940 123770 661180
rect 123860 660940 124100 661180
rect 124190 660940 124430 661180
rect 124520 660940 124760 661180
rect 124870 660940 125110 661180
rect 125200 660940 125440 661180
rect 125530 660940 125770 661180
rect 125860 660940 126100 661180
rect 126210 660940 126450 661180
rect 126540 660940 126780 661180
rect 126870 660940 127110 661180
rect 127200 660940 127440 661180
rect 127550 660940 127790 661180
rect 127880 660940 128120 661180
rect 128210 660940 128450 661180
rect 128540 660940 128780 661180
rect 128890 660940 129130 661180
rect 129220 660940 129460 661180
rect 129550 660940 129790 661180
rect 129880 660940 130120 661180
rect 130230 660940 130470 661180
rect 130560 660940 130800 661180
rect 130890 660940 131130 661180
rect 131220 660940 131460 661180
rect 131570 660940 131810 661180
rect 131900 660940 132140 661180
rect 132230 660940 132470 661180
rect 132560 660940 132800 661180
rect 132910 660940 133150 661180
rect 133570 671660 133810 671900
rect 133900 671660 134140 671900
rect 134230 671660 134470 671900
rect 134560 671660 134800 671900
rect 134910 671660 135150 671900
rect 135240 671660 135480 671900
rect 135570 671660 135810 671900
rect 135900 671660 136140 671900
rect 136250 671660 136490 671900
rect 136580 671660 136820 671900
rect 136910 671660 137150 671900
rect 137240 671660 137480 671900
rect 137590 671660 137830 671900
rect 137920 671660 138160 671900
rect 138250 671660 138490 671900
rect 138580 671660 138820 671900
rect 138930 671660 139170 671900
rect 139260 671660 139500 671900
rect 139590 671660 139830 671900
rect 139920 671660 140160 671900
rect 140270 671660 140510 671900
rect 140600 671660 140840 671900
rect 140930 671660 141170 671900
rect 141260 671660 141500 671900
rect 141610 671660 141850 671900
rect 141940 671660 142180 671900
rect 142270 671660 142510 671900
rect 142600 671660 142840 671900
rect 142950 671660 143190 671900
rect 143280 671660 143520 671900
rect 143610 671660 143850 671900
rect 143940 671660 144180 671900
rect 144290 671660 144530 671900
rect 133570 671310 133810 671550
rect 133900 671310 134140 671550
rect 134230 671310 134470 671550
rect 134560 671310 134800 671550
rect 134910 671310 135150 671550
rect 135240 671310 135480 671550
rect 135570 671310 135810 671550
rect 135900 671310 136140 671550
rect 136250 671310 136490 671550
rect 136580 671310 136820 671550
rect 136910 671310 137150 671550
rect 137240 671310 137480 671550
rect 137590 671310 137830 671550
rect 137920 671310 138160 671550
rect 138250 671310 138490 671550
rect 138580 671310 138820 671550
rect 138930 671310 139170 671550
rect 139260 671310 139500 671550
rect 139590 671310 139830 671550
rect 139920 671310 140160 671550
rect 140270 671310 140510 671550
rect 140600 671310 140840 671550
rect 140930 671310 141170 671550
rect 141260 671310 141500 671550
rect 141610 671310 141850 671550
rect 141940 671310 142180 671550
rect 142270 671310 142510 671550
rect 142600 671310 142840 671550
rect 142950 671310 143190 671550
rect 143280 671310 143520 671550
rect 143610 671310 143850 671550
rect 143940 671310 144180 671550
rect 144290 671310 144530 671550
rect 133570 670980 133810 671220
rect 133900 670980 134140 671220
rect 134230 670980 134470 671220
rect 134560 670980 134800 671220
rect 134910 670980 135150 671220
rect 135240 670980 135480 671220
rect 135570 670980 135810 671220
rect 135900 670980 136140 671220
rect 136250 670980 136490 671220
rect 136580 670980 136820 671220
rect 136910 670980 137150 671220
rect 137240 670980 137480 671220
rect 137590 670980 137830 671220
rect 137920 670980 138160 671220
rect 138250 670980 138490 671220
rect 138580 670980 138820 671220
rect 138930 670980 139170 671220
rect 139260 670980 139500 671220
rect 139590 670980 139830 671220
rect 139920 670980 140160 671220
rect 140270 670980 140510 671220
rect 140600 670980 140840 671220
rect 140930 670980 141170 671220
rect 141260 670980 141500 671220
rect 141610 670980 141850 671220
rect 141940 670980 142180 671220
rect 142270 670980 142510 671220
rect 142600 670980 142840 671220
rect 142950 670980 143190 671220
rect 143280 670980 143520 671220
rect 143610 670980 143850 671220
rect 143940 670980 144180 671220
rect 144290 670980 144530 671220
rect 133570 670650 133810 670890
rect 133900 670650 134140 670890
rect 134230 670650 134470 670890
rect 134560 670650 134800 670890
rect 134910 670650 135150 670890
rect 135240 670650 135480 670890
rect 135570 670650 135810 670890
rect 135900 670650 136140 670890
rect 136250 670650 136490 670890
rect 136580 670650 136820 670890
rect 136910 670650 137150 670890
rect 137240 670650 137480 670890
rect 137590 670650 137830 670890
rect 137920 670650 138160 670890
rect 138250 670650 138490 670890
rect 138580 670650 138820 670890
rect 138930 670650 139170 670890
rect 139260 670650 139500 670890
rect 139590 670650 139830 670890
rect 139920 670650 140160 670890
rect 140270 670650 140510 670890
rect 140600 670650 140840 670890
rect 140930 670650 141170 670890
rect 141260 670650 141500 670890
rect 141610 670650 141850 670890
rect 141940 670650 142180 670890
rect 142270 670650 142510 670890
rect 142600 670650 142840 670890
rect 142950 670650 143190 670890
rect 143280 670650 143520 670890
rect 143610 670650 143850 670890
rect 143940 670650 144180 670890
rect 144290 670650 144530 670890
rect 133570 670320 133810 670560
rect 133900 670320 134140 670560
rect 134230 670320 134470 670560
rect 134560 670320 134800 670560
rect 134910 670320 135150 670560
rect 135240 670320 135480 670560
rect 135570 670320 135810 670560
rect 135900 670320 136140 670560
rect 136250 670320 136490 670560
rect 136580 670320 136820 670560
rect 136910 670320 137150 670560
rect 137240 670320 137480 670560
rect 137590 670320 137830 670560
rect 137920 670320 138160 670560
rect 138250 670320 138490 670560
rect 138580 670320 138820 670560
rect 138930 670320 139170 670560
rect 139260 670320 139500 670560
rect 139590 670320 139830 670560
rect 139920 670320 140160 670560
rect 140270 670320 140510 670560
rect 140600 670320 140840 670560
rect 140930 670320 141170 670560
rect 141260 670320 141500 670560
rect 141610 670320 141850 670560
rect 141940 670320 142180 670560
rect 142270 670320 142510 670560
rect 142600 670320 142840 670560
rect 142950 670320 143190 670560
rect 143280 670320 143520 670560
rect 143610 670320 143850 670560
rect 143940 670320 144180 670560
rect 144290 670320 144530 670560
rect 133570 669970 133810 670210
rect 133900 669970 134140 670210
rect 134230 669970 134470 670210
rect 134560 669970 134800 670210
rect 134910 669970 135150 670210
rect 135240 669970 135480 670210
rect 135570 669970 135810 670210
rect 135900 669970 136140 670210
rect 136250 669970 136490 670210
rect 136580 669970 136820 670210
rect 136910 669970 137150 670210
rect 137240 669970 137480 670210
rect 137590 669970 137830 670210
rect 137920 669970 138160 670210
rect 138250 669970 138490 670210
rect 138580 669970 138820 670210
rect 138930 669970 139170 670210
rect 139260 669970 139500 670210
rect 139590 669970 139830 670210
rect 139920 669970 140160 670210
rect 140270 669970 140510 670210
rect 140600 669970 140840 670210
rect 140930 669970 141170 670210
rect 141260 669970 141500 670210
rect 141610 669970 141850 670210
rect 141940 669970 142180 670210
rect 142270 669970 142510 670210
rect 142600 669970 142840 670210
rect 142950 669970 143190 670210
rect 143280 669970 143520 670210
rect 143610 669970 143850 670210
rect 143940 669970 144180 670210
rect 144290 669970 144530 670210
rect 133570 669640 133810 669880
rect 133900 669640 134140 669880
rect 134230 669640 134470 669880
rect 134560 669640 134800 669880
rect 134910 669640 135150 669880
rect 135240 669640 135480 669880
rect 135570 669640 135810 669880
rect 135900 669640 136140 669880
rect 136250 669640 136490 669880
rect 136580 669640 136820 669880
rect 136910 669640 137150 669880
rect 137240 669640 137480 669880
rect 137590 669640 137830 669880
rect 137920 669640 138160 669880
rect 138250 669640 138490 669880
rect 138580 669640 138820 669880
rect 138930 669640 139170 669880
rect 139260 669640 139500 669880
rect 139590 669640 139830 669880
rect 139920 669640 140160 669880
rect 140270 669640 140510 669880
rect 140600 669640 140840 669880
rect 140930 669640 141170 669880
rect 141260 669640 141500 669880
rect 141610 669640 141850 669880
rect 141940 669640 142180 669880
rect 142270 669640 142510 669880
rect 142600 669640 142840 669880
rect 142950 669640 143190 669880
rect 143280 669640 143520 669880
rect 143610 669640 143850 669880
rect 143940 669640 144180 669880
rect 144290 669640 144530 669880
rect 133570 669310 133810 669550
rect 133900 669310 134140 669550
rect 134230 669310 134470 669550
rect 134560 669310 134800 669550
rect 134910 669310 135150 669550
rect 135240 669310 135480 669550
rect 135570 669310 135810 669550
rect 135900 669310 136140 669550
rect 136250 669310 136490 669550
rect 136580 669310 136820 669550
rect 136910 669310 137150 669550
rect 137240 669310 137480 669550
rect 137590 669310 137830 669550
rect 137920 669310 138160 669550
rect 138250 669310 138490 669550
rect 138580 669310 138820 669550
rect 138930 669310 139170 669550
rect 139260 669310 139500 669550
rect 139590 669310 139830 669550
rect 139920 669310 140160 669550
rect 140270 669310 140510 669550
rect 140600 669310 140840 669550
rect 140930 669310 141170 669550
rect 141260 669310 141500 669550
rect 141610 669310 141850 669550
rect 141940 669310 142180 669550
rect 142270 669310 142510 669550
rect 142600 669310 142840 669550
rect 142950 669310 143190 669550
rect 143280 669310 143520 669550
rect 143610 669310 143850 669550
rect 143940 669310 144180 669550
rect 144290 669310 144530 669550
rect 133570 668980 133810 669220
rect 133900 668980 134140 669220
rect 134230 668980 134470 669220
rect 134560 668980 134800 669220
rect 134910 668980 135150 669220
rect 135240 668980 135480 669220
rect 135570 668980 135810 669220
rect 135900 668980 136140 669220
rect 136250 668980 136490 669220
rect 136580 668980 136820 669220
rect 136910 668980 137150 669220
rect 137240 668980 137480 669220
rect 137590 668980 137830 669220
rect 137920 668980 138160 669220
rect 138250 668980 138490 669220
rect 138580 668980 138820 669220
rect 138930 668980 139170 669220
rect 139260 668980 139500 669220
rect 139590 668980 139830 669220
rect 139920 668980 140160 669220
rect 140270 668980 140510 669220
rect 140600 668980 140840 669220
rect 140930 668980 141170 669220
rect 141260 668980 141500 669220
rect 141610 668980 141850 669220
rect 141940 668980 142180 669220
rect 142270 668980 142510 669220
rect 142600 668980 142840 669220
rect 142950 668980 143190 669220
rect 143280 668980 143520 669220
rect 143610 668980 143850 669220
rect 143940 668980 144180 669220
rect 144290 668980 144530 669220
rect 133570 668630 133810 668870
rect 133900 668630 134140 668870
rect 134230 668630 134470 668870
rect 134560 668630 134800 668870
rect 134910 668630 135150 668870
rect 135240 668630 135480 668870
rect 135570 668630 135810 668870
rect 135900 668630 136140 668870
rect 136250 668630 136490 668870
rect 136580 668630 136820 668870
rect 136910 668630 137150 668870
rect 137240 668630 137480 668870
rect 137590 668630 137830 668870
rect 137920 668630 138160 668870
rect 138250 668630 138490 668870
rect 138580 668630 138820 668870
rect 138930 668630 139170 668870
rect 139260 668630 139500 668870
rect 139590 668630 139830 668870
rect 139920 668630 140160 668870
rect 140270 668630 140510 668870
rect 140600 668630 140840 668870
rect 140930 668630 141170 668870
rect 141260 668630 141500 668870
rect 141610 668630 141850 668870
rect 141940 668630 142180 668870
rect 142270 668630 142510 668870
rect 142600 668630 142840 668870
rect 142950 668630 143190 668870
rect 143280 668630 143520 668870
rect 143610 668630 143850 668870
rect 143940 668630 144180 668870
rect 144290 668630 144530 668870
rect 133570 668300 133810 668540
rect 133900 668300 134140 668540
rect 134230 668300 134470 668540
rect 134560 668300 134800 668540
rect 134910 668300 135150 668540
rect 135240 668300 135480 668540
rect 135570 668300 135810 668540
rect 135900 668300 136140 668540
rect 136250 668300 136490 668540
rect 136580 668300 136820 668540
rect 136910 668300 137150 668540
rect 137240 668300 137480 668540
rect 137590 668300 137830 668540
rect 137920 668300 138160 668540
rect 138250 668300 138490 668540
rect 138580 668300 138820 668540
rect 138930 668300 139170 668540
rect 139260 668300 139500 668540
rect 139590 668300 139830 668540
rect 139920 668300 140160 668540
rect 140270 668300 140510 668540
rect 140600 668300 140840 668540
rect 140930 668300 141170 668540
rect 141260 668300 141500 668540
rect 141610 668300 141850 668540
rect 141940 668300 142180 668540
rect 142270 668300 142510 668540
rect 142600 668300 142840 668540
rect 142950 668300 143190 668540
rect 143280 668300 143520 668540
rect 143610 668300 143850 668540
rect 143940 668300 144180 668540
rect 144290 668300 144530 668540
rect 133570 667970 133810 668210
rect 133900 667970 134140 668210
rect 134230 667970 134470 668210
rect 134560 667970 134800 668210
rect 134910 667970 135150 668210
rect 135240 667970 135480 668210
rect 135570 667970 135810 668210
rect 135900 667970 136140 668210
rect 136250 667970 136490 668210
rect 136580 667970 136820 668210
rect 136910 667970 137150 668210
rect 137240 667970 137480 668210
rect 137590 667970 137830 668210
rect 137920 667970 138160 668210
rect 138250 667970 138490 668210
rect 138580 667970 138820 668210
rect 138930 667970 139170 668210
rect 139260 667970 139500 668210
rect 139590 667970 139830 668210
rect 139920 667970 140160 668210
rect 140270 667970 140510 668210
rect 140600 667970 140840 668210
rect 140930 667970 141170 668210
rect 141260 667970 141500 668210
rect 141610 667970 141850 668210
rect 141940 667970 142180 668210
rect 142270 667970 142510 668210
rect 142600 667970 142840 668210
rect 142950 667970 143190 668210
rect 143280 667970 143520 668210
rect 143610 667970 143850 668210
rect 143940 667970 144180 668210
rect 144290 667970 144530 668210
rect 133570 667640 133810 667880
rect 133900 667640 134140 667880
rect 134230 667640 134470 667880
rect 134560 667640 134800 667880
rect 134910 667640 135150 667880
rect 135240 667640 135480 667880
rect 135570 667640 135810 667880
rect 135900 667640 136140 667880
rect 136250 667640 136490 667880
rect 136580 667640 136820 667880
rect 136910 667640 137150 667880
rect 137240 667640 137480 667880
rect 137590 667640 137830 667880
rect 137920 667640 138160 667880
rect 138250 667640 138490 667880
rect 138580 667640 138820 667880
rect 138930 667640 139170 667880
rect 139260 667640 139500 667880
rect 139590 667640 139830 667880
rect 139920 667640 140160 667880
rect 140270 667640 140510 667880
rect 140600 667640 140840 667880
rect 140930 667640 141170 667880
rect 141260 667640 141500 667880
rect 141610 667640 141850 667880
rect 141940 667640 142180 667880
rect 142270 667640 142510 667880
rect 142600 667640 142840 667880
rect 142950 667640 143190 667880
rect 143280 667640 143520 667880
rect 143610 667640 143850 667880
rect 143940 667640 144180 667880
rect 144290 667640 144530 667880
rect 133570 667290 133810 667530
rect 133900 667290 134140 667530
rect 134230 667290 134470 667530
rect 134560 667290 134800 667530
rect 134910 667290 135150 667530
rect 135240 667290 135480 667530
rect 135570 667290 135810 667530
rect 135900 667290 136140 667530
rect 136250 667290 136490 667530
rect 136580 667290 136820 667530
rect 136910 667290 137150 667530
rect 137240 667290 137480 667530
rect 137590 667290 137830 667530
rect 137920 667290 138160 667530
rect 138250 667290 138490 667530
rect 138580 667290 138820 667530
rect 138930 667290 139170 667530
rect 139260 667290 139500 667530
rect 139590 667290 139830 667530
rect 139920 667290 140160 667530
rect 140270 667290 140510 667530
rect 140600 667290 140840 667530
rect 140930 667290 141170 667530
rect 141260 667290 141500 667530
rect 141610 667290 141850 667530
rect 141940 667290 142180 667530
rect 142270 667290 142510 667530
rect 142600 667290 142840 667530
rect 142950 667290 143190 667530
rect 143280 667290 143520 667530
rect 143610 667290 143850 667530
rect 143940 667290 144180 667530
rect 144290 667290 144530 667530
rect 133570 666960 133810 667200
rect 133900 666960 134140 667200
rect 134230 666960 134470 667200
rect 134560 666960 134800 667200
rect 134910 666960 135150 667200
rect 135240 666960 135480 667200
rect 135570 666960 135810 667200
rect 135900 666960 136140 667200
rect 136250 666960 136490 667200
rect 136580 666960 136820 667200
rect 136910 666960 137150 667200
rect 137240 666960 137480 667200
rect 137590 666960 137830 667200
rect 137920 666960 138160 667200
rect 138250 666960 138490 667200
rect 138580 666960 138820 667200
rect 138930 666960 139170 667200
rect 139260 666960 139500 667200
rect 139590 666960 139830 667200
rect 139920 666960 140160 667200
rect 140270 666960 140510 667200
rect 140600 666960 140840 667200
rect 140930 666960 141170 667200
rect 141260 666960 141500 667200
rect 141610 666960 141850 667200
rect 141940 666960 142180 667200
rect 142270 666960 142510 667200
rect 142600 666960 142840 667200
rect 142950 666960 143190 667200
rect 143280 666960 143520 667200
rect 143610 666960 143850 667200
rect 143940 666960 144180 667200
rect 144290 666960 144530 667200
rect 133570 666630 133810 666870
rect 133900 666630 134140 666870
rect 134230 666630 134470 666870
rect 134560 666630 134800 666870
rect 134910 666630 135150 666870
rect 135240 666630 135480 666870
rect 135570 666630 135810 666870
rect 135900 666630 136140 666870
rect 136250 666630 136490 666870
rect 136580 666630 136820 666870
rect 136910 666630 137150 666870
rect 137240 666630 137480 666870
rect 137590 666630 137830 666870
rect 137920 666630 138160 666870
rect 138250 666630 138490 666870
rect 138580 666630 138820 666870
rect 138930 666630 139170 666870
rect 139260 666630 139500 666870
rect 139590 666630 139830 666870
rect 139920 666630 140160 666870
rect 140270 666630 140510 666870
rect 140600 666630 140840 666870
rect 140930 666630 141170 666870
rect 141260 666630 141500 666870
rect 141610 666630 141850 666870
rect 141940 666630 142180 666870
rect 142270 666630 142510 666870
rect 142600 666630 142840 666870
rect 142950 666630 143190 666870
rect 143280 666630 143520 666870
rect 143610 666630 143850 666870
rect 143940 666630 144180 666870
rect 144290 666630 144530 666870
rect 133570 666300 133810 666540
rect 133900 666300 134140 666540
rect 134230 666300 134470 666540
rect 134560 666300 134800 666540
rect 134910 666300 135150 666540
rect 135240 666300 135480 666540
rect 135570 666300 135810 666540
rect 135900 666300 136140 666540
rect 136250 666300 136490 666540
rect 136580 666300 136820 666540
rect 136910 666300 137150 666540
rect 137240 666300 137480 666540
rect 137590 666300 137830 666540
rect 137920 666300 138160 666540
rect 138250 666300 138490 666540
rect 138580 666300 138820 666540
rect 138930 666300 139170 666540
rect 139260 666300 139500 666540
rect 139590 666300 139830 666540
rect 139920 666300 140160 666540
rect 140270 666300 140510 666540
rect 140600 666300 140840 666540
rect 140930 666300 141170 666540
rect 141260 666300 141500 666540
rect 141610 666300 141850 666540
rect 141940 666300 142180 666540
rect 142270 666300 142510 666540
rect 142600 666300 142840 666540
rect 142950 666300 143190 666540
rect 143280 666300 143520 666540
rect 143610 666300 143850 666540
rect 143940 666300 144180 666540
rect 144290 666300 144530 666540
rect 133570 665950 133810 666190
rect 133900 665950 134140 666190
rect 134230 665950 134470 666190
rect 134560 665950 134800 666190
rect 134910 665950 135150 666190
rect 135240 665950 135480 666190
rect 135570 665950 135810 666190
rect 135900 665950 136140 666190
rect 136250 665950 136490 666190
rect 136580 665950 136820 666190
rect 136910 665950 137150 666190
rect 137240 665950 137480 666190
rect 137590 665950 137830 666190
rect 137920 665950 138160 666190
rect 138250 665950 138490 666190
rect 138580 665950 138820 666190
rect 138930 665950 139170 666190
rect 139260 665950 139500 666190
rect 139590 665950 139830 666190
rect 139920 665950 140160 666190
rect 140270 665950 140510 666190
rect 140600 665950 140840 666190
rect 140930 665950 141170 666190
rect 141260 665950 141500 666190
rect 141610 665950 141850 666190
rect 141940 665950 142180 666190
rect 142270 665950 142510 666190
rect 142600 665950 142840 666190
rect 142950 665950 143190 666190
rect 143280 665950 143520 666190
rect 143610 665950 143850 666190
rect 143940 665950 144180 666190
rect 144290 665950 144530 666190
rect 133570 665620 133810 665860
rect 133900 665620 134140 665860
rect 134230 665620 134470 665860
rect 134560 665620 134800 665860
rect 134910 665620 135150 665860
rect 135240 665620 135480 665860
rect 135570 665620 135810 665860
rect 135900 665620 136140 665860
rect 136250 665620 136490 665860
rect 136580 665620 136820 665860
rect 136910 665620 137150 665860
rect 137240 665620 137480 665860
rect 137590 665620 137830 665860
rect 137920 665620 138160 665860
rect 138250 665620 138490 665860
rect 138580 665620 138820 665860
rect 138930 665620 139170 665860
rect 139260 665620 139500 665860
rect 139590 665620 139830 665860
rect 139920 665620 140160 665860
rect 140270 665620 140510 665860
rect 140600 665620 140840 665860
rect 140930 665620 141170 665860
rect 141260 665620 141500 665860
rect 141610 665620 141850 665860
rect 141940 665620 142180 665860
rect 142270 665620 142510 665860
rect 142600 665620 142840 665860
rect 142950 665620 143190 665860
rect 143280 665620 143520 665860
rect 143610 665620 143850 665860
rect 143940 665620 144180 665860
rect 144290 665620 144530 665860
rect 133570 665290 133810 665530
rect 133900 665290 134140 665530
rect 134230 665290 134470 665530
rect 134560 665290 134800 665530
rect 134910 665290 135150 665530
rect 135240 665290 135480 665530
rect 135570 665290 135810 665530
rect 135900 665290 136140 665530
rect 136250 665290 136490 665530
rect 136580 665290 136820 665530
rect 136910 665290 137150 665530
rect 137240 665290 137480 665530
rect 137590 665290 137830 665530
rect 137920 665290 138160 665530
rect 138250 665290 138490 665530
rect 138580 665290 138820 665530
rect 138930 665290 139170 665530
rect 139260 665290 139500 665530
rect 139590 665290 139830 665530
rect 139920 665290 140160 665530
rect 140270 665290 140510 665530
rect 140600 665290 140840 665530
rect 140930 665290 141170 665530
rect 141260 665290 141500 665530
rect 141610 665290 141850 665530
rect 141940 665290 142180 665530
rect 142270 665290 142510 665530
rect 142600 665290 142840 665530
rect 142950 665290 143190 665530
rect 143280 665290 143520 665530
rect 143610 665290 143850 665530
rect 143940 665290 144180 665530
rect 144290 665290 144530 665530
rect 133570 664960 133810 665200
rect 133900 664960 134140 665200
rect 134230 664960 134470 665200
rect 134560 664960 134800 665200
rect 134910 664960 135150 665200
rect 135240 664960 135480 665200
rect 135570 664960 135810 665200
rect 135900 664960 136140 665200
rect 136250 664960 136490 665200
rect 136580 664960 136820 665200
rect 136910 664960 137150 665200
rect 137240 664960 137480 665200
rect 137590 664960 137830 665200
rect 137920 664960 138160 665200
rect 138250 664960 138490 665200
rect 138580 664960 138820 665200
rect 138930 664960 139170 665200
rect 139260 664960 139500 665200
rect 139590 664960 139830 665200
rect 139920 664960 140160 665200
rect 140270 664960 140510 665200
rect 140600 664960 140840 665200
rect 140930 664960 141170 665200
rect 141260 664960 141500 665200
rect 141610 664960 141850 665200
rect 141940 664960 142180 665200
rect 142270 664960 142510 665200
rect 142600 664960 142840 665200
rect 142950 664960 143190 665200
rect 143280 664960 143520 665200
rect 143610 664960 143850 665200
rect 143940 664960 144180 665200
rect 144290 664960 144530 665200
rect 133570 664610 133810 664850
rect 133900 664610 134140 664850
rect 134230 664610 134470 664850
rect 134560 664610 134800 664850
rect 134910 664610 135150 664850
rect 135240 664610 135480 664850
rect 135570 664610 135810 664850
rect 135900 664610 136140 664850
rect 136250 664610 136490 664850
rect 136580 664610 136820 664850
rect 136910 664610 137150 664850
rect 137240 664610 137480 664850
rect 137590 664610 137830 664850
rect 137920 664610 138160 664850
rect 138250 664610 138490 664850
rect 138580 664610 138820 664850
rect 138930 664610 139170 664850
rect 139260 664610 139500 664850
rect 139590 664610 139830 664850
rect 139920 664610 140160 664850
rect 140270 664610 140510 664850
rect 140600 664610 140840 664850
rect 140930 664610 141170 664850
rect 141260 664610 141500 664850
rect 141610 664610 141850 664850
rect 141940 664610 142180 664850
rect 142270 664610 142510 664850
rect 142600 664610 142840 664850
rect 142950 664610 143190 664850
rect 143280 664610 143520 664850
rect 143610 664610 143850 664850
rect 143940 664610 144180 664850
rect 144290 664610 144530 664850
rect 133570 664280 133810 664520
rect 133900 664280 134140 664520
rect 134230 664280 134470 664520
rect 134560 664280 134800 664520
rect 134910 664280 135150 664520
rect 135240 664280 135480 664520
rect 135570 664280 135810 664520
rect 135900 664280 136140 664520
rect 136250 664280 136490 664520
rect 136580 664280 136820 664520
rect 136910 664280 137150 664520
rect 137240 664280 137480 664520
rect 137590 664280 137830 664520
rect 137920 664280 138160 664520
rect 138250 664280 138490 664520
rect 138580 664280 138820 664520
rect 138930 664280 139170 664520
rect 139260 664280 139500 664520
rect 139590 664280 139830 664520
rect 139920 664280 140160 664520
rect 140270 664280 140510 664520
rect 140600 664280 140840 664520
rect 140930 664280 141170 664520
rect 141260 664280 141500 664520
rect 141610 664280 141850 664520
rect 141940 664280 142180 664520
rect 142270 664280 142510 664520
rect 142600 664280 142840 664520
rect 142950 664280 143190 664520
rect 143280 664280 143520 664520
rect 143610 664280 143850 664520
rect 143940 664280 144180 664520
rect 144290 664280 144530 664520
rect 133570 663950 133810 664190
rect 133900 663950 134140 664190
rect 134230 663950 134470 664190
rect 134560 663950 134800 664190
rect 134910 663950 135150 664190
rect 135240 663950 135480 664190
rect 135570 663950 135810 664190
rect 135900 663950 136140 664190
rect 136250 663950 136490 664190
rect 136580 663950 136820 664190
rect 136910 663950 137150 664190
rect 137240 663950 137480 664190
rect 137590 663950 137830 664190
rect 137920 663950 138160 664190
rect 138250 663950 138490 664190
rect 138580 663950 138820 664190
rect 138930 663950 139170 664190
rect 139260 663950 139500 664190
rect 139590 663950 139830 664190
rect 139920 663950 140160 664190
rect 140270 663950 140510 664190
rect 140600 663950 140840 664190
rect 140930 663950 141170 664190
rect 141260 663950 141500 664190
rect 141610 663950 141850 664190
rect 141940 663950 142180 664190
rect 142270 663950 142510 664190
rect 142600 663950 142840 664190
rect 142950 663950 143190 664190
rect 143280 663950 143520 664190
rect 143610 663950 143850 664190
rect 143940 663950 144180 664190
rect 144290 663950 144530 664190
rect 133570 663620 133810 663860
rect 133900 663620 134140 663860
rect 134230 663620 134470 663860
rect 134560 663620 134800 663860
rect 134910 663620 135150 663860
rect 135240 663620 135480 663860
rect 135570 663620 135810 663860
rect 135900 663620 136140 663860
rect 136250 663620 136490 663860
rect 136580 663620 136820 663860
rect 136910 663620 137150 663860
rect 137240 663620 137480 663860
rect 137590 663620 137830 663860
rect 137920 663620 138160 663860
rect 138250 663620 138490 663860
rect 138580 663620 138820 663860
rect 138930 663620 139170 663860
rect 139260 663620 139500 663860
rect 139590 663620 139830 663860
rect 139920 663620 140160 663860
rect 140270 663620 140510 663860
rect 140600 663620 140840 663860
rect 140930 663620 141170 663860
rect 141260 663620 141500 663860
rect 141610 663620 141850 663860
rect 141940 663620 142180 663860
rect 142270 663620 142510 663860
rect 142600 663620 142840 663860
rect 142950 663620 143190 663860
rect 143280 663620 143520 663860
rect 143610 663620 143850 663860
rect 143940 663620 144180 663860
rect 144290 663620 144530 663860
rect 133570 663270 133810 663510
rect 133900 663270 134140 663510
rect 134230 663270 134470 663510
rect 134560 663270 134800 663510
rect 134910 663270 135150 663510
rect 135240 663270 135480 663510
rect 135570 663270 135810 663510
rect 135900 663270 136140 663510
rect 136250 663270 136490 663510
rect 136580 663270 136820 663510
rect 136910 663270 137150 663510
rect 137240 663270 137480 663510
rect 137590 663270 137830 663510
rect 137920 663270 138160 663510
rect 138250 663270 138490 663510
rect 138580 663270 138820 663510
rect 138930 663270 139170 663510
rect 139260 663270 139500 663510
rect 139590 663270 139830 663510
rect 139920 663270 140160 663510
rect 140270 663270 140510 663510
rect 140600 663270 140840 663510
rect 140930 663270 141170 663510
rect 141260 663270 141500 663510
rect 141610 663270 141850 663510
rect 141940 663270 142180 663510
rect 142270 663270 142510 663510
rect 142600 663270 142840 663510
rect 142950 663270 143190 663510
rect 143280 663270 143520 663510
rect 143610 663270 143850 663510
rect 143940 663270 144180 663510
rect 144290 663270 144530 663510
rect 133570 662940 133810 663180
rect 133900 662940 134140 663180
rect 134230 662940 134470 663180
rect 134560 662940 134800 663180
rect 134910 662940 135150 663180
rect 135240 662940 135480 663180
rect 135570 662940 135810 663180
rect 135900 662940 136140 663180
rect 136250 662940 136490 663180
rect 136580 662940 136820 663180
rect 136910 662940 137150 663180
rect 137240 662940 137480 663180
rect 137590 662940 137830 663180
rect 137920 662940 138160 663180
rect 138250 662940 138490 663180
rect 138580 662940 138820 663180
rect 138930 662940 139170 663180
rect 139260 662940 139500 663180
rect 139590 662940 139830 663180
rect 139920 662940 140160 663180
rect 140270 662940 140510 663180
rect 140600 662940 140840 663180
rect 140930 662940 141170 663180
rect 141260 662940 141500 663180
rect 141610 662940 141850 663180
rect 141940 662940 142180 663180
rect 142270 662940 142510 663180
rect 142600 662940 142840 663180
rect 142950 662940 143190 663180
rect 143280 662940 143520 663180
rect 143610 662940 143850 663180
rect 143940 662940 144180 663180
rect 144290 662940 144530 663180
rect 133570 662610 133810 662850
rect 133900 662610 134140 662850
rect 134230 662610 134470 662850
rect 134560 662610 134800 662850
rect 134910 662610 135150 662850
rect 135240 662610 135480 662850
rect 135570 662610 135810 662850
rect 135900 662610 136140 662850
rect 136250 662610 136490 662850
rect 136580 662610 136820 662850
rect 136910 662610 137150 662850
rect 137240 662610 137480 662850
rect 137590 662610 137830 662850
rect 137920 662610 138160 662850
rect 138250 662610 138490 662850
rect 138580 662610 138820 662850
rect 138930 662610 139170 662850
rect 139260 662610 139500 662850
rect 139590 662610 139830 662850
rect 139920 662610 140160 662850
rect 140270 662610 140510 662850
rect 140600 662610 140840 662850
rect 140930 662610 141170 662850
rect 141260 662610 141500 662850
rect 141610 662610 141850 662850
rect 141940 662610 142180 662850
rect 142270 662610 142510 662850
rect 142600 662610 142840 662850
rect 142950 662610 143190 662850
rect 143280 662610 143520 662850
rect 143610 662610 143850 662850
rect 143940 662610 144180 662850
rect 144290 662610 144530 662850
rect 133570 662280 133810 662520
rect 133900 662280 134140 662520
rect 134230 662280 134470 662520
rect 134560 662280 134800 662520
rect 134910 662280 135150 662520
rect 135240 662280 135480 662520
rect 135570 662280 135810 662520
rect 135900 662280 136140 662520
rect 136250 662280 136490 662520
rect 136580 662280 136820 662520
rect 136910 662280 137150 662520
rect 137240 662280 137480 662520
rect 137590 662280 137830 662520
rect 137920 662280 138160 662520
rect 138250 662280 138490 662520
rect 138580 662280 138820 662520
rect 138930 662280 139170 662520
rect 139260 662280 139500 662520
rect 139590 662280 139830 662520
rect 139920 662280 140160 662520
rect 140270 662280 140510 662520
rect 140600 662280 140840 662520
rect 140930 662280 141170 662520
rect 141260 662280 141500 662520
rect 141610 662280 141850 662520
rect 141940 662280 142180 662520
rect 142270 662280 142510 662520
rect 142600 662280 142840 662520
rect 142950 662280 143190 662520
rect 143280 662280 143520 662520
rect 143610 662280 143850 662520
rect 143940 662280 144180 662520
rect 144290 662280 144530 662520
rect 133570 661930 133810 662170
rect 133900 661930 134140 662170
rect 134230 661930 134470 662170
rect 134560 661930 134800 662170
rect 134910 661930 135150 662170
rect 135240 661930 135480 662170
rect 135570 661930 135810 662170
rect 135900 661930 136140 662170
rect 136250 661930 136490 662170
rect 136580 661930 136820 662170
rect 136910 661930 137150 662170
rect 137240 661930 137480 662170
rect 137590 661930 137830 662170
rect 137920 661930 138160 662170
rect 138250 661930 138490 662170
rect 138580 661930 138820 662170
rect 138930 661930 139170 662170
rect 139260 661930 139500 662170
rect 139590 661930 139830 662170
rect 139920 661930 140160 662170
rect 140270 661930 140510 662170
rect 140600 661930 140840 662170
rect 140930 661930 141170 662170
rect 141260 661930 141500 662170
rect 141610 661930 141850 662170
rect 141940 661930 142180 662170
rect 142270 661930 142510 662170
rect 142600 661930 142840 662170
rect 142950 661930 143190 662170
rect 143280 661930 143520 662170
rect 143610 661930 143850 662170
rect 143940 661930 144180 662170
rect 144290 661930 144530 662170
rect 133570 661600 133810 661840
rect 133900 661600 134140 661840
rect 134230 661600 134470 661840
rect 134560 661600 134800 661840
rect 134910 661600 135150 661840
rect 135240 661600 135480 661840
rect 135570 661600 135810 661840
rect 135900 661600 136140 661840
rect 136250 661600 136490 661840
rect 136580 661600 136820 661840
rect 136910 661600 137150 661840
rect 137240 661600 137480 661840
rect 137590 661600 137830 661840
rect 137920 661600 138160 661840
rect 138250 661600 138490 661840
rect 138580 661600 138820 661840
rect 138930 661600 139170 661840
rect 139260 661600 139500 661840
rect 139590 661600 139830 661840
rect 139920 661600 140160 661840
rect 140270 661600 140510 661840
rect 140600 661600 140840 661840
rect 140930 661600 141170 661840
rect 141260 661600 141500 661840
rect 141610 661600 141850 661840
rect 141940 661600 142180 661840
rect 142270 661600 142510 661840
rect 142600 661600 142840 661840
rect 142950 661600 143190 661840
rect 143280 661600 143520 661840
rect 143610 661600 143850 661840
rect 143940 661600 144180 661840
rect 144290 661600 144530 661840
rect 133570 661270 133810 661510
rect 133900 661270 134140 661510
rect 134230 661270 134470 661510
rect 134560 661270 134800 661510
rect 134910 661270 135150 661510
rect 135240 661270 135480 661510
rect 135570 661270 135810 661510
rect 135900 661270 136140 661510
rect 136250 661270 136490 661510
rect 136580 661270 136820 661510
rect 136910 661270 137150 661510
rect 137240 661270 137480 661510
rect 137590 661270 137830 661510
rect 137920 661270 138160 661510
rect 138250 661270 138490 661510
rect 138580 661270 138820 661510
rect 138930 661270 139170 661510
rect 139260 661270 139500 661510
rect 139590 661270 139830 661510
rect 139920 661270 140160 661510
rect 140270 661270 140510 661510
rect 140600 661270 140840 661510
rect 140930 661270 141170 661510
rect 141260 661270 141500 661510
rect 141610 661270 141850 661510
rect 141940 661270 142180 661510
rect 142270 661270 142510 661510
rect 142600 661270 142840 661510
rect 142950 661270 143190 661510
rect 143280 661270 143520 661510
rect 143610 661270 143850 661510
rect 143940 661270 144180 661510
rect 144290 661270 144530 661510
rect 133570 660940 133810 661180
rect 133900 660940 134140 661180
rect 134230 660940 134470 661180
rect 134560 660940 134800 661180
rect 134910 660940 135150 661180
rect 135240 660940 135480 661180
rect 135570 660940 135810 661180
rect 135900 660940 136140 661180
rect 136250 660940 136490 661180
rect 136580 660940 136820 661180
rect 136910 660940 137150 661180
rect 137240 660940 137480 661180
rect 137590 660940 137830 661180
rect 137920 660940 138160 661180
rect 138250 660940 138490 661180
rect 138580 660940 138820 661180
rect 138930 660940 139170 661180
rect 139260 660940 139500 661180
rect 139590 660940 139830 661180
rect 139920 660940 140160 661180
rect 140270 660940 140510 661180
rect 140600 660940 140840 661180
rect 140930 660940 141170 661180
rect 141260 660940 141500 661180
rect 141610 660940 141850 661180
rect 141940 660940 142180 661180
rect 142270 660940 142510 661180
rect 142600 660940 142840 661180
rect 142950 660940 143190 661180
rect 143280 660940 143520 661180
rect 143610 660940 143850 661180
rect 143940 660940 144180 661180
rect 144290 660940 144530 661180
rect 144950 671660 145190 671900
rect 145280 671660 145520 671900
rect 145610 671660 145850 671900
rect 145940 671660 146180 671900
rect 146290 671660 146530 671900
rect 146620 671660 146860 671900
rect 146950 671660 147190 671900
rect 147280 671660 147520 671900
rect 147630 671660 147870 671900
rect 147960 671660 148200 671900
rect 148290 671660 148530 671900
rect 148620 671660 148860 671900
rect 148970 671660 149210 671900
rect 149300 671660 149540 671900
rect 149630 671660 149870 671900
rect 149960 671660 150200 671900
rect 150310 671660 150550 671900
rect 150640 671660 150880 671900
rect 150970 671660 151210 671900
rect 151300 671660 151540 671900
rect 151650 671660 151890 671900
rect 151980 671660 152220 671900
rect 152310 671660 152550 671900
rect 152640 671660 152880 671900
rect 152990 671660 153230 671900
rect 153320 671660 153560 671900
rect 153650 671660 153890 671900
rect 153980 671660 154220 671900
rect 154330 671660 154570 671900
rect 154660 671660 154900 671900
rect 154990 671660 155230 671900
rect 155320 671660 155560 671900
rect 155670 671660 155910 671900
rect 144950 671310 145190 671550
rect 145280 671310 145520 671550
rect 145610 671310 145850 671550
rect 145940 671310 146180 671550
rect 146290 671310 146530 671550
rect 146620 671310 146860 671550
rect 146950 671310 147190 671550
rect 147280 671310 147520 671550
rect 147630 671310 147870 671550
rect 147960 671310 148200 671550
rect 148290 671310 148530 671550
rect 148620 671310 148860 671550
rect 148970 671310 149210 671550
rect 149300 671310 149540 671550
rect 149630 671310 149870 671550
rect 149960 671310 150200 671550
rect 150310 671310 150550 671550
rect 150640 671310 150880 671550
rect 150970 671310 151210 671550
rect 151300 671310 151540 671550
rect 151650 671310 151890 671550
rect 151980 671310 152220 671550
rect 152310 671310 152550 671550
rect 152640 671310 152880 671550
rect 152990 671310 153230 671550
rect 153320 671310 153560 671550
rect 153650 671310 153890 671550
rect 153980 671310 154220 671550
rect 154330 671310 154570 671550
rect 154660 671310 154900 671550
rect 154990 671310 155230 671550
rect 155320 671310 155560 671550
rect 155670 671310 155910 671550
rect 144950 670980 145190 671220
rect 145280 670980 145520 671220
rect 145610 670980 145850 671220
rect 145940 670980 146180 671220
rect 146290 670980 146530 671220
rect 146620 670980 146860 671220
rect 146950 670980 147190 671220
rect 147280 670980 147520 671220
rect 147630 670980 147870 671220
rect 147960 670980 148200 671220
rect 148290 670980 148530 671220
rect 148620 670980 148860 671220
rect 148970 670980 149210 671220
rect 149300 670980 149540 671220
rect 149630 670980 149870 671220
rect 149960 670980 150200 671220
rect 150310 670980 150550 671220
rect 150640 670980 150880 671220
rect 150970 670980 151210 671220
rect 151300 670980 151540 671220
rect 151650 670980 151890 671220
rect 151980 670980 152220 671220
rect 152310 670980 152550 671220
rect 152640 670980 152880 671220
rect 152990 670980 153230 671220
rect 153320 670980 153560 671220
rect 153650 670980 153890 671220
rect 153980 670980 154220 671220
rect 154330 670980 154570 671220
rect 154660 670980 154900 671220
rect 154990 670980 155230 671220
rect 155320 670980 155560 671220
rect 155670 670980 155910 671220
rect 144950 670650 145190 670890
rect 145280 670650 145520 670890
rect 145610 670650 145850 670890
rect 145940 670650 146180 670890
rect 146290 670650 146530 670890
rect 146620 670650 146860 670890
rect 146950 670650 147190 670890
rect 147280 670650 147520 670890
rect 147630 670650 147870 670890
rect 147960 670650 148200 670890
rect 148290 670650 148530 670890
rect 148620 670650 148860 670890
rect 148970 670650 149210 670890
rect 149300 670650 149540 670890
rect 149630 670650 149870 670890
rect 149960 670650 150200 670890
rect 150310 670650 150550 670890
rect 150640 670650 150880 670890
rect 150970 670650 151210 670890
rect 151300 670650 151540 670890
rect 151650 670650 151890 670890
rect 151980 670650 152220 670890
rect 152310 670650 152550 670890
rect 152640 670650 152880 670890
rect 152990 670650 153230 670890
rect 153320 670650 153560 670890
rect 153650 670650 153890 670890
rect 153980 670650 154220 670890
rect 154330 670650 154570 670890
rect 154660 670650 154900 670890
rect 154990 670650 155230 670890
rect 155320 670650 155560 670890
rect 155670 670650 155910 670890
rect 144950 670320 145190 670560
rect 145280 670320 145520 670560
rect 145610 670320 145850 670560
rect 145940 670320 146180 670560
rect 146290 670320 146530 670560
rect 146620 670320 146860 670560
rect 146950 670320 147190 670560
rect 147280 670320 147520 670560
rect 147630 670320 147870 670560
rect 147960 670320 148200 670560
rect 148290 670320 148530 670560
rect 148620 670320 148860 670560
rect 148970 670320 149210 670560
rect 149300 670320 149540 670560
rect 149630 670320 149870 670560
rect 149960 670320 150200 670560
rect 150310 670320 150550 670560
rect 150640 670320 150880 670560
rect 150970 670320 151210 670560
rect 151300 670320 151540 670560
rect 151650 670320 151890 670560
rect 151980 670320 152220 670560
rect 152310 670320 152550 670560
rect 152640 670320 152880 670560
rect 152990 670320 153230 670560
rect 153320 670320 153560 670560
rect 153650 670320 153890 670560
rect 153980 670320 154220 670560
rect 154330 670320 154570 670560
rect 154660 670320 154900 670560
rect 154990 670320 155230 670560
rect 155320 670320 155560 670560
rect 155670 670320 155910 670560
rect 144950 669970 145190 670210
rect 145280 669970 145520 670210
rect 145610 669970 145850 670210
rect 145940 669970 146180 670210
rect 146290 669970 146530 670210
rect 146620 669970 146860 670210
rect 146950 669970 147190 670210
rect 147280 669970 147520 670210
rect 147630 669970 147870 670210
rect 147960 669970 148200 670210
rect 148290 669970 148530 670210
rect 148620 669970 148860 670210
rect 148970 669970 149210 670210
rect 149300 669970 149540 670210
rect 149630 669970 149870 670210
rect 149960 669970 150200 670210
rect 150310 669970 150550 670210
rect 150640 669970 150880 670210
rect 150970 669970 151210 670210
rect 151300 669970 151540 670210
rect 151650 669970 151890 670210
rect 151980 669970 152220 670210
rect 152310 669970 152550 670210
rect 152640 669970 152880 670210
rect 152990 669970 153230 670210
rect 153320 669970 153560 670210
rect 153650 669970 153890 670210
rect 153980 669970 154220 670210
rect 154330 669970 154570 670210
rect 154660 669970 154900 670210
rect 154990 669970 155230 670210
rect 155320 669970 155560 670210
rect 155670 669970 155910 670210
rect 144950 669640 145190 669880
rect 145280 669640 145520 669880
rect 145610 669640 145850 669880
rect 145940 669640 146180 669880
rect 146290 669640 146530 669880
rect 146620 669640 146860 669880
rect 146950 669640 147190 669880
rect 147280 669640 147520 669880
rect 147630 669640 147870 669880
rect 147960 669640 148200 669880
rect 148290 669640 148530 669880
rect 148620 669640 148860 669880
rect 148970 669640 149210 669880
rect 149300 669640 149540 669880
rect 149630 669640 149870 669880
rect 149960 669640 150200 669880
rect 150310 669640 150550 669880
rect 150640 669640 150880 669880
rect 150970 669640 151210 669880
rect 151300 669640 151540 669880
rect 151650 669640 151890 669880
rect 151980 669640 152220 669880
rect 152310 669640 152550 669880
rect 152640 669640 152880 669880
rect 152990 669640 153230 669880
rect 153320 669640 153560 669880
rect 153650 669640 153890 669880
rect 153980 669640 154220 669880
rect 154330 669640 154570 669880
rect 154660 669640 154900 669880
rect 154990 669640 155230 669880
rect 155320 669640 155560 669880
rect 155670 669640 155910 669880
rect 144950 669310 145190 669550
rect 145280 669310 145520 669550
rect 145610 669310 145850 669550
rect 145940 669310 146180 669550
rect 146290 669310 146530 669550
rect 146620 669310 146860 669550
rect 146950 669310 147190 669550
rect 147280 669310 147520 669550
rect 147630 669310 147870 669550
rect 147960 669310 148200 669550
rect 148290 669310 148530 669550
rect 148620 669310 148860 669550
rect 148970 669310 149210 669550
rect 149300 669310 149540 669550
rect 149630 669310 149870 669550
rect 149960 669310 150200 669550
rect 150310 669310 150550 669550
rect 150640 669310 150880 669550
rect 150970 669310 151210 669550
rect 151300 669310 151540 669550
rect 151650 669310 151890 669550
rect 151980 669310 152220 669550
rect 152310 669310 152550 669550
rect 152640 669310 152880 669550
rect 152990 669310 153230 669550
rect 153320 669310 153560 669550
rect 153650 669310 153890 669550
rect 153980 669310 154220 669550
rect 154330 669310 154570 669550
rect 154660 669310 154900 669550
rect 154990 669310 155230 669550
rect 155320 669310 155560 669550
rect 155670 669310 155910 669550
rect 144950 668980 145190 669220
rect 145280 668980 145520 669220
rect 145610 668980 145850 669220
rect 145940 668980 146180 669220
rect 146290 668980 146530 669220
rect 146620 668980 146860 669220
rect 146950 668980 147190 669220
rect 147280 668980 147520 669220
rect 147630 668980 147870 669220
rect 147960 668980 148200 669220
rect 148290 668980 148530 669220
rect 148620 668980 148860 669220
rect 148970 668980 149210 669220
rect 149300 668980 149540 669220
rect 149630 668980 149870 669220
rect 149960 668980 150200 669220
rect 150310 668980 150550 669220
rect 150640 668980 150880 669220
rect 150970 668980 151210 669220
rect 151300 668980 151540 669220
rect 151650 668980 151890 669220
rect 151980 668980 152220 669220
rect 152310 668980 152550 669220
rect 152640 668980 152880 669220
rect 152990 668980 153230 669220
rect 153320 668980 153560 669220
rect 153650 668980 153890 669220
rect 153980 668980 154220 669220
rect 154330 668980 154570 669220
rect 154660 668980 154900 669220
rect 154990 668980 155230 669220
rect 155320 668980 155560 669220
rect 155670 668980 155910 669220
rect 144950 668630 145190 668870
rect 145280 668630 145520 668870
rect 145610 668630 145850 668870
rect 145940 668630 146180 668870
rect 146290 668630 146530 668870
rect 146620 668630 146860 668870
rect 146950 668630 147190 668870
rect 147280 668630 147520 668870
rect 147630 668630 147870 668870
rect 147960 668630 148200 668870
rect 148290 668630 148530 668870
rect 148620 668630 148860 668870
rect 148970 668630 149210 668870
rect 149300 668630 149540 668870
rect 149630 668630 149870 668870
rect 149960 668630 150200 668870
rect 150310 668630 150550 668870
rect 150640 668630 150880 668870
rect 150970 668630 151210 668870
rect 151300 668630 151540 668870
rect 151650 668630 151890 668870
rect 151980 668630 152220 668870
rect 152310 668630 152550 668870
rect 152640 668630 152880 668870
rect 152990 668630 153230 668870
rect 153320 668630 153560 668870
rect 153650 668630 153890 668870
rect 153980 668630 154220 668870
rect 154330 668630 154570 668870
rect 154660 668630 154900 668870
rect 154990 668630 155230 668870
rect 155320 668630 155560 668870
rect 155670 668630 155910 668870
rect 144950 668300 145190 668540
rect 145280 668300 145520 668540
rect 145610 668300 145850 668540
rect 145940 668300 146180 668540
rect 146290 668300 146530 668540
rect 146620 668300 146860 668540
rect 146950 668300 147190 668540
rect 147280 668300 147520 668540
rect 147630 668300 147870 668540
rect 147960 668300 148200 668540
rect 148290 668300 148530 668540
rect 148620 668300 148860 668540
rect 148970 668300 149210 668540
rect 149300 668300 149540 668540
rect 149630 668300 149870 668540
rect 149960 668300 150200 668540
rect 150310 668300 150550 668540
rect 150640 668300 150880 668540
rect 150970 668300 151210 668540
rect 151300 668300 151540 668540
rect 151650 668300 151890 668540
rect 151980 668300 152220 668540
rect 152310 668300 152550 668540
rect 152640 668300 152880 668540
rect 152990 668300 153230 668540
rect 153320 668300 153560 668540
rect 153650 668300 153890 668540
rect 153980 668300 154220 668540
rect 154330 668300 154570 668540
rect 154660 668300 154900 668540
rect 154990 668300 155230 668540
rect 155320 668300 155560 668540
rect 155670 668300 155910 668540
rect 144950 667970 145190 668210
rect 145280 667970 145520 668210
rect 145610 667970 145850 668210
rect 145940 667970 146180 668210
rect 146290 667970 146530 668210
rect 146620 667970 146860 668210
rect 146950 667970 147190 668210
rect 147280 667970 147520 668210
rect 147630 667970 147870 668210
rect 147960 667970 148200 668210
rect 148290 667970 148530 668210
rect 148620 667970 148860 668210
rect 148970 667970 149210 668210
rect 149300 667970 149540 668210
rect 149630 667970 149870 668210
rect 149960 667970 150200 668210
rect 150310 667970 150550 668210
rect 150640 667970 150880 668210
rect 150970 667970 151210 668210
rect 151300 667970 151540 668210
rect 151650 667970 151890 668210
rect 151980 667970 152220 668210
rect 152310 667970 152550 668210
rect 152640 667970 152880 668210
rect 152990 667970 153230 668210
rect 153320 667970 153560 668210
rect 153650 667970 153890 668210
rect 153980 667970 154220 668210
rect 154330 667970 154570 668210
rect 154660 667970 154900 668210
rect 154990 667970 155230 668210
rect 155320 667970 155560 668210
rect 155670 667970 155910 668210
rect 144950 667640 145190 667880
rect 145280 667640 145520 667880
rect 145610 667640 145850 667880
rect 145940 667640 146180 667880
rect 146290 667640 146530 667880
rect 146620 667640 146860 667880
rect 146950 667640 147190 667880
rect 147280 667640 147520 667880
rect 147630 667640 147870 667880
rect 147960 667640 148200 667880
rect 148290 667640 148530 667880
rect 148620 667640 148860 667880
rect 148970 667640 149210 667880
rect 149300 667640 149540 667880
rect 149630 667640 149870 667880
rect 149960 667640 150200 667880
rect 150310 667640 150550 667880
rect 150640 667640 150880 667880
rect 150970 667640 151210 667880
rect 151300 667640 151540 667880
rect 151650 667640 151890 667880
rect 151980 667640 152220 667880
rect 152310 667640 152550 667880
rect 152640 667640 152880 667880
rect 152990 667640 153230 667880
rect 153320 667640 153560 667880
rect 153650 667640 153890 667880
rect 153980 667640 154220 667880
rect 154330 667640 154570 667880
rect 154660 667640 154900 667880
rect 154990 667640 155230 667880
rect 155320 667640 155560 667880
rect 155670 667640 155910 667880
rect 144950 667290 145190 667530
rect 145280 667290 145520 667530
rect 145610 667290 145850 667530
rect 145940 667290 146180 667530
rect 146290 667290 146530 667530
rect 146620 667290 146860 667530
rect 146950 667290 147190 667530
rect 147280 667290 147520 667530
rect 147630 667290 147870 667530
rect 147960 667290 148200 667530
rect 148290 667290 148530 667530
rect 148620 667290 148860 667530
rect 148970 667290 149210 667530
rect 149300 667290 149540 667530
rect 149630 667290 149870 667530
rect 149960 667290 150200 667530
rect 150310 667290 150550 667530
rect 150640 667290 150880 667530
rect 150970 667290 151210 667530
rect 151300 667290 151540 667530
rect 151650 667290 151890 667530
rect 151980 667290 152220 667530
rect 152310 667290 152550 667530
rect 152640 667290 152880 667530
rect 152990 667290 153230 667530
rect 153320 667290 153560 667530
rect 153650 667290 153890 667530
rect 153980 667290 154220 667530
rect 154330 667290 154570 667530
rect 154660 667290 154900 667530
rect 154990 667290 155230 667530
rect 155320 667290 155560 667530
rect 155670 667290 155910 667530
rect 144950 666960 145190 667200
rect 145280 666960 145520 667200
rect 145610 666960 145850 667200
rect 145940 666960 146180 667200
rect 146290 666960 146530 667200
rect 146620 666960 146860 667200
rect 146950 666960 147190 667200
rect 147280 666960 147520 667200
rect 147630 666960 147870 667200
rect 147960 666960 148200 667200
rect 148290 666960 148530 667200
rect 148620 666960 148860 667200
rect 148970 666960 149210 667200
rect 149300 666960 149540 667200
rect 149630 666960 149870 667200
rect 149960 666960 150200 667200
rect 150310 666960 150550 667200
rect 150640 666960 150880 667200
rect 150970 666960 151210 667200
rect 151300 666960 151540 667200
rect 151650 666960 151890 667200
rect 151980 666960 152220 667200
rect 152310 666960 152550 667200
rect 152640 666960 152880 667200
rect 152990 666960 153230 667200
rect 153320 666960 153560 667200
rect 153650 666960 153890 667200
rect 153980 666960 154220 667200
rect 154330 666960 154570 667200
rect 154660 666960 154900 667200
rect 154990 666960 155230 667200
rect 155320 666960 155560 667200
rect 155670 666960 155910 667200
rect 144950 666630 145190 666870
rect 145280 666630 145520 666870
rect 145610 666630 145850 666870
rect 145940 666630 146180 666870
rect 146290 666630 146530 666870
rect 146620 666630 146860 666870
rect 146950 666630 147190 666870
rect 147280 666630 147520 666870
rect 147630 666630 147870 666870
rect 147960 666630 148200 666870
rect 148290 666630 148530 666870
rect 148620 666630 148860 666870
rect 148970 666630 149210 666870
rect 149300 666630 149540 666870
rect 149630 666630 149870 666870
rect 149960 666630 150200 666870
rect 150310 666630 150550 666870
rect 150640 666630 150880 666870
rect 150970 666630 151210 666870
rect 151300 666630 151540 666870
rect 151650 666630 151890 666870
rect 151980 666630 152220 666870
rect 152310 666630 152550 666870
rect 152640 666630 152880 666870
rect 152990 666630 153230 666870
rect 153320 666630 153560 666870
rect 153650 666630 153890 666870
rect 153980 666630 154220 666870
rect 154330 666630 154570 666870
rect 154660 666630 154900 666870
rect 154990 666630 155230 666870
rect 155320 666630 155560 666870
rect 155670 666630 155910 666870
rect 144950 666300 145190 666540
rect 145280 666300 145520 666540
rect 145610 666300 145850 666540
rect 145940 666300 146180 666540
rect 146290 666300 146530 666540
rect 146620 666300 146860 666540
rect 146950 666300 147190 666540
rect 147280 666300 147520 666540
rect 147630 666300 147870 666540
rect 147960 666300 148200 666540
rect 148290 666300 148530 666540
rect 148620 666300 148860 666540
rect 148970 666300 149210 666540
rect 149300 666300 149540 666540
rect 149630 666300 149870 666540
rect 149960 666300 150200 666540
rect 150310 666300 150550 666540
rect 150640 666300 150880 666540
rect 150970 666300 151210 666540
rect 151300 666300 151540 666540
rect 151650 666300 151890 666540
rect 151980 666300 152220 666540
rect 152310 666300 152550 666540
rect 152640 666300 152880 666540
rect 152990 666300 153230 666540
rect 153320 666300 153560 666540
rect 153650 666300 153890 666540
rect 153980 666300 154220 666540
rect 154330 666300 154570 666540
rect 154660 666300 154900 666540
rect 154990 666300 155230 666540
rect 155320 666300 155560 666540
rect 155670 666300 155910 666540
rect 144950 665950 145190 666190
rect 145280 665950 145520 666190
rect 145610 665950 145850 666190
rect 145940 665950 146180 666190
rect 146290 665950 146530 666190
rect 146620 665950 146860 666190
rect 146950 665950 147190 666190
rect 147280 665950 147520 666190
rect 147630 665950 147870 666190
rect 147960 665950 148200 666190
rect 148290 665950 148530 666190
rect 148620 665950 148860 666190
rect 148970 665950 149210 666190
rect 149300 665950 149540 666190
rect 149630 665950 149870 666190
rect 149960 665950 150200 666190
rect 150310 665950 150550 666190
rect 150640 665950 150880 666190
rect 150970 665950 151210 666190
rect 151300 665950 151540 666190
rect 151650 665950 151890 666190
rect 151980 665950 152220 666190
rect 152310 665950 152550 666190
rect 152640 665950 152880 666190
rect 152990 665950 153230 666190
rect 153320 665950 153560 666190
rect 153650 665950 153890 666190
rect 153980 665950 154220 666190
rect 154330 665950 154570 666190
rect 154660 665950 154900 666190
rect 154990 665950 155230 666190
rect 155320 665950 155560 666190
rect 155670 665950 155910 666190
rect 144950 665620 145190 665860
rect 145280 665620 145520 665860
rect 145610 665620 145850 665860
rect 145940 665620 146180 665860
rect 146290 665620 146530 665860
rect 146620 665620 146860 665860
rect 146950 665620 147190 665860
rect 147280 665620 147520 665860
rect 147630 665620 147870 665860
rect 147960 665620 148200 665860
rect 148290 665620 148530 665860
rect 148620 665620 148860 665860
rect 148970 665620 149210 665860
rect 149300 665620 149540 665860
rect 149630 665620 149870 665860
rect 149960 665620 150200 665860
rect 150310 665620 150550 665860
rect 150640 665620 150880 665860
rect 150970 665620 151210 665860
rect 151300 665620 151540 665860
rect 151650 665620 151890 665860
rect 151980 665620 152220 665860
rect 152310 665620 152550 665860
rect 152640 665620 152880 665860
rect 152990 665620 153230 665860
rect 153320 665620 153560 665860
rect 153650 665620 153890 665860
rect 153980 665620 154220 665860
rect 154330 665620 154570 665860
rect 154660 665620 154900 665860
rect 154990 665620 155230 665860
rect 155320 665620 155560 665860
rect 155670 665620 155910 665860
rect 144950 665290 145190 665530
rect 145280 665290 145520 665530
rect 145610 665290 145850 665530
rect 145940 665290 146180 665530
rect 146290 665290 146530 665530
rect 146620 665290 146860 665530
rect 146950 665290 147190 665530
rect 147280 665290 147520 665530
rect 147630 665290 147870 665530
rect 147960 665290 148200 665530
rect 148290 665290 148530 665530
rect 148620 665290 148860 665530
rect 148970 665290 149210 665530
rect 149300 665290 149540 665530
rect 149630 665290 149870 665530
rect 149960 665290 150200 665530
rect 150310 665290 150550 665530
rect 150640 665290 150880 665530
rect 150970 665290 151210 665530
rect 151300 665290 151540 665530
rect 151650 665290 151890 665530
rect 151980 665290 152220 665530
rect 152310 665290 152550 665530
rect 152640 665290 152880 665530
rect 152990 665290 153230 665530
rect 153320 665290 153560 665530
rect 153650 665290 153890 665530
rect 153980 665290 154220 665530
rect 154330 665290 154570 665530
rect 154660 665290 154900 665530
rect 154990 665290 155230 665530
rect 155320 665290 155560 665530
rect 155670 665290 155910 665530
rect 144950 664960 145190 665200
rect 145280 664960 145520 665200
rect 145610 664960 145850 665200
rect 145940 664960 146180 665200
rect 146290 664960 146530 665200
rect 146620 664960 146860 665200
rect 146950 664960 147190 665200
rect 147280 664960 147520 665200
rect 147630 664960 147870 665200
rect 147960 664960 148200 665200
rect 148290 664960 148530 665200
rect 148620 664960 148860 665200
rect 148970 664960 149210 665200
rect 149300 664960 149540 665200
rect 149630 664960 149870 665200
rect 149960 664960 150200 665200
rect 150310 664960 150550 665200
rect 150640 664960 150880 665200
rect 150970 664960 151210 665200
rect 151300 664960 151540 665200
rect 151650 664960 151890 665200
rect 151980 664960 152220 665200
rect 152310 664960 152550 665200
rect 152640 664960 152880 665200
rect 152990 664960 153230 665200
rect 153320 664960 153560 665200
rect 153650 664960 153890 665200
rect 153980 664960 154220 665200
rect 154330 664960 154570 665200
rect 154660 664960 154900 665200
rect 154990 664960 155230 665200
rect 155320 664960 155560 665200
rect 155670 664960 155910 665200
rect 144950 664610 145190 664850
rect 145280 664610 145520 664850
rect 145610 664610 145850 664850
rect 145940 664610 146180 664850
rect 146290 664610 146530 664850
rect 146620 664610 146860 664850
rect 146950 664610 147190 664850
rect 147280 664610 147520 664850
rect 147630 664610 147870 664850
rect 147960 664610 148200 664850
rect 148290 664610 148530 664850
rect 148620 664610 148860 664850
rect 148970 664610 149210 664850
rect 149300 664610 149540 664850
rect 149630 664610 149870 664850
rect 149960 664610 150200 664850
rect 150310 664610 150550 664850
rect 150640 664610 150880 664850
rect 150970 664610 151210 664850
rect 151300 664610 151540 664850
rect 151650 664610 151890 664850
rect 151980 664610 152220 664850
rect 152310 664610 152550 664850
rect 152640 664610 152880 664850
rect 152990 664610 153230 664850
rect 153320 664610 153560 664850
rect 153650 664610 153890 664850
rect 153980 664610 154220 664850
rect 154330 664610 154570 664850
rect 154660 664610 154900 664850
rect 154990 664610 155230 664850
rect 155320 664610 155560 664850
rect 155670 664610 155910 664850
rect 144950 664280 145190 664520
rect 145280 664280 145520 664520
rect 145610 664280 145850 664520
rect 145940 664280 146180 664520
rect 146290 664280 146530 664520
rect 146620 664280 146860 664520
rect 146950 664280 147190 664520
rect 147280 664280 147520 664520
rect 147630 664280 147870 664520
rect 147960 664280 148200 664520
rect 148290 664280 148530 664520
rect 148620 664280 148860 664520
rect 148970 664280 149210 664520
rect 149300 664280 149540 664520
rect 149630 664280 149870 664520
rect 149960 664280 150200 664520
rect 150310 664280 150550 664520
rect 150640 664280 150880 664520
rect 150970 664280 151210 664520
rect 151300 664280 151540 664520
rect 151650 664280 151890 664520
rect 151980 664280 152220 664520
rect 152310 664280 152550 664520
rect 152640 664280 152880 664520
rect 152990 664280 153230 664520
rect 153320 664280 153560 664520
rect 153650 664280 153890 664520
rect 153980 664280 154220 664520
rect 154330 664280 154570 664520
rect 154660 664280 154900 664520
rect 154990 664280 155230 664520
rect 155320 664280 155560 664520
rect 155670 664280 155910 664520
rect 144950 663950 145190 664190
rect 145280 663950 145520 664190
rect 145610 663950 145850 664190
rect 145940 663950 146180 664190
rect 146290 663950 146530 664190
rect 146620 663950 146860 664190
rect 146950 663950 147190 664190
rect 147280 663950 147520 664190
rect 147630 663950 147870 664190
rect 147960 663950 148200 664190
rect 148290 663950 148530 664190
rect 148620 663950 148860 664190
rect 148970 663950 149210 664190
rect 149300 663950 149540 664190
rect 149630 663950 149870 664190
rect 149960 663950 150200 664190
rect 150310 663950 150550 664190
rect 150640 663950 150880 664190
rect 150970 663950 151210 664190
rect 151300 663950 151540 664190
rect 151650 663950 151890 664190
rect 151980 663950 152220 664190
rect 152310 663950 152550 664190
rect 152640 663950 152880 664190
rect 152990 663950 153230 664190
rect 153320 663950 153560 664190
rect 153650 663950 153890 664190
rect 153980 663950 154220 664190
rect 154330 663950 154570 664190
rect 154660 663950 154900 664190
rect 154990 663950 155230 664190
rect 155320 663950 155560 664190
rect 155670 663950 155910 664190
rect 144950 663620 145190 663860
rect 145280 663620 145520 663860
rect 145610 663620 145850 663860
rect 145940 663620 146180 663860
rect 146290 663620 146530 663860
rect 146620 663620 146860 663860
rect 146950 663620 147190 663860
rect 147280 663620 147520 663860
rect 147630 663620 147870 663860
rect 147960 663620 148200 663860
rect 148290 663620 148530 663860
rect 148620 663620 148860 663860
rect 148970 663620 149210 663860
rect 149300 663620 149540 663860
rect 149630 663620 149870 663860
rect 149960 663620 150200 663860
rect 150310 663620 150550 663860
rect 150640 663620 150880 663860
rect 150970 663620 151210 663860
rect 151300 663620 151540 663860
rect 151650 663620 151890 663860
rect 151980 663620 152220 663860
rect 152310 663620 152550 663860
rect 152640 663620 152880 663860
rect 152990 663620 153230 663860
rect 153320 663620 153560 663860
rect 153650 663620 153890 663860
rect 153980 663620 154220 663860
rect 154330 663620 154570 663860
rect 154660 663620 154900 663860
rect 154990 663620 155230 663860
rect 155320 663620 155560 663860
rect 155670 663620 155910 663860
rect 144950 663270 145190 663510
rect 145280 663270 145520 663510
rect 145610 663270 145850 663510
rect 145940 663270 146180 663510
rect 146290 663270 146530 663510
rect 146620 663270 146860 663510
rect 146950 663270 147190 663510
rect 147280 663270 147520 663510
rect 147630 663270 147870 663510
rect 147960 663270 148200 663510
rect 148290 663270 148530 663510
rect 148620 663270 148860 663510
rect 148970 663270 149210 663510
rect 149300 663270 149540 663510
rect 149630 663270 149870 663510
rect 149960 663270 150200 663510
rect 150310 663270 150550 663510
rect 150640 663270 150880 663510
rect 150970 663270 151210 663510
rect 151300 663270 151540 663510
rect 151650 663270 151890 663510
rect 151980 663270 152220 663510
rect 152310 663270 152550 663510
rect 152640 663270 152880 663510
rect 152990 663270 153230 663510
rect 153320 663270 153560 663510
rect 153650 663270 153890 663510
rect 153980 663270 154220 663510
rect 154330 663270 154570 663510
rect 154660 663270 154900 663510
rect 154990 663270 155230 663510
rect 155320 663270 155560 663510
rect 155670 663270 155910 663510
rect 144950 662940 145190 663180
rect 145280 662940 145520 663180
rect 145610 662940 145850 663180
rect 145940 662940 146180 663180
rect 146290 662940 146530 663180
rect 146620 662940 146860 663180
rect 146950 662940 147190 663180
rect 147280 662940 147520 663180
rect 147630 662940 147870 663180
rect 147960 662940 148200 663180
rect 148290 662940 148530 663180
rect 148620 662940 148860 663180
rect 148970 662940 149210 663180
rect 149300 662940 149540 663180
rect 149630 662940 149870 663180
rect 149960 662940 150200 663180
rect 150310 662940 150550 663180
rect 150640 662940 150880 663180
rect 150970 662940 151210 663180
rect 151300 662940 151540 663180
rect 151650 662940 151890 663180
rect 151980 662940 152220 663180
rect 152310 662940 152550 663180
rect 152640 662940 152880 663180
rect 152990 662940 153230 663180
rect 153320 662940 153560 663180
rect 153650 662940 153890 663180
rect 153980 662940 154220 663180
rect 154330 662940 154570 663180
rect 154660 662940 154900 663180
rect 154990 662940 155230 663180
rect 155320 662940 155560 663180
rect 155670 662940 155910 663180
rect 144950 662610 145190 662850
rect 145280 662610 145520 662850
rect 145610 662610 145850 662850
rect 145940 662610 146180 662850
rect 146290 662610 146530 662850
rect 146620 662610 146860 662850
rect 146950 662610 147190 662850
rect 147280 662610 147520 662850
rect 147630 662610 147870 662850
rect 147960 662610 148200 662850
rect 148290 662610 148530 662850
rect 148620 662610 148860 662850
rect 148970 662610 149210 662850
rect 149300 662610 149540 662850
rect 149630 662610 149870 662850
rect 149960 662610 150200 662850
rect 150310 662610 150550 662850
rect 150640 662610 150880 662850
rect 150970 662610 151210 662850
rect 151300 662610 151540 662850
rect 151650 662610 151890 662850
rect 151980 662610 152220 662850
rect 152310 662610 152550 662850
rect 152640 662610 152880 662850
rect 152990 662610 153230 662850
rect 153320 662610 153560 662850
rect 153650 662610 153890 662850
rect 153980 662610 154220 662850
rect 154330 662610 154570 662850
rect 154660 662610 154900 662850
rect 154990 662610 155230 662850
rect 155320 662610 155560 662850
rect 155670 662610 155910 662850
rect 144950 662280 145190 662520
rect 145280 662280 145520 662520
rect 145610 662280 145850 662520
rect 145940 662280 146180 662520
rect 146290 662280 146530 662520
rect 146620 662280 146860 662520
rect 146950 662280 147190 662520
rect 147280 662280 147520 662520
rect 147630 662280 147870 662520
rect 147960 662280 148200 662520
rect 148290 662280 148530 662520
rect 148620 662280 148860 662520
rect 148970 662280 149210 662520
rect 149300 662280 149540 662520
rect 149630 662280 149870 662520
rect 149960 662280 150200 662520
rect 150310 662280 150550 662520
rect 150640 662280 150880 662520
rect 150970 662280 151210 662520
rect 151300 662280 151540 662520
rect 151650 662280 151890 662520
rect 151980 662280 152220 662520
rect 152310 662280 152550 662520
rect 152640 662280 152880 662520
rect 152990 662280 153230 662520
rect 153320 662280 153560 662520
rect 153650 662280 153890 662520
rect 153980 662280 154220 662520
rect 154330 662280 154570 662520
rect 154660 662280 154900 662520
rect 154990 662280 155230 662520
rect 155320 662280 155560 662520
rect 155670 662280 155910 662520
rect 144950 661930 145190 662170
rect 145280 661930 145520 662170
rect 145610 661930 145850 662170
rect 145940 661930 146180 662170
rect 146290 661930 146530 662170
rect 146620 661930 146860 662170
rect 146950 661930 147190 662170
rect 147280 661930 147520 662170
rect 147630 661930 147870 662170
rect 147960 661930 148200 662170
rect 148290 661930 148530 662170
rect 148620 661930 148860 662170
rect 148970 661930 149210 662170
rect 149300 661930 149540 662170
rect 149630 661930 149870 662170
rect 149960 661930 150200 662170
rect 150310 661930 150550 662170
rect 150640 661930 150880 662170
rect 150970 661930 151210 662170
rect 151300 661930 151540 662170
rect 151650 661930 151890 662170
rect 151980 661930 152220 662170
rect 152310 661930 152550 662170
rect 152640 661930 152880 662170
rect 152990 661930 153230 662170
rect 153320 661930 153560 662170
rect 153650 661930 153890 662170
rect 153980 661930 154220 662170
rect 154330 661930 154570 662170
rect 154660 661930 154900 662170
rect 154990 661930 155230 662170
rect 155320 661930 155560 662170
rect 155670 661930 155910 662170
rect 144950 661600 145190 661840
rect 145280 661600 145520 661840
rect 145610 661600 145850 661840
rect 145940 661600 146180 661840
rect 146290 661600 146530 661840
rect 146620 661600 146860 661840
rect 146950 661600 147190 661840
rect 147280 661600 147520 661840
rect 147630 661600 147870 661840
rect 147960 661600 148200 661840
rect 148290 661600 148530 661840
rect 148620 661600 148860 661840
rect 148970 661600 149210 661840
rect 149300 661600 149540 661840
rect 149630 661600 149870 661840
rect 149960 661600 150200 661840
rect 150310 661600 150550 661840
rect 150640 661600 150880 661840
rect 150970 661600 151210 661840
rect 151300 661600 151540 661840
rect 151650 661600 151890 661840
rect 151980 661600 152220 661840
rect 152310 661600 152550 661840
rect 152640 661600 152880 661840
rect 152990 661600 153230 661840
rect 153320 661600 153560 661840
rect 153650 661600 153890 661840
rect 153980 661600 154220 661840
rect 154330 661600 154570 661840
rect 154660 661600 154900 661840
rect 154990 661600 155230 661840
rect 155320 661600 155560 661840
rect 155670 661600 155910 661840
rect 144950 661270 145190 661510
rect 145280 661270 145520 661510
rect 145610 661270 145850 661510
rect 145940 661270 146180 661510
rect 146290 661270 146530 661510
rect 146620 661270 146860 661510
rect 146950 661270 147190 661510
rect 147280 661270 147520 661510
rect 147630 661270 147870 661510
rect 147960 661270 148200 661510
rect 148290 661270 148530 661510
rect 148620 661270 148860 661510
rect 148970 661270 149210 661510
rect 149300 661270 149540 661510
rect 149630 661270 149870 661510
rect 149960 661270 150200 661510
rect 150310 661270 150550 661510
rect 150640 661270 150880 661510
rect 150970 661270 151210 661510
rect 151300 661270 151540 661510
rect 151650 661270 151890 661510
rect 151980 661270 152220 661510
rect 152310 661270 152550 661510
rect 152640 661270 152880 661510
rect 152990 661270 153230 661510
rect 153320 661270 153560 661510
rect 153650 661270 153890 661510
rect 153980 661270 154220 661510
rect 154330 661270 154570 661510
rect 154660 661270 154900 661510
rect 154990 661270 155230 661510
rect 155320 661270 155560 661510
rect 155670 661270 155910 661510
rect 144950 660940 145190 661180
rect 145280 660940 145520 661180
rect 145610 660940 145850 661180
rect 145940 660940 146180 661180
rect 146290 660940 146530 661180
rect 146620 660940 146860 661180
rect 146950 660940 147190 661180
rect 147280 660940 147520 661180
rect 147630 660940 147870 661180
rect 147960 660940 148200 661180
rect 148290 660940 148530 661180
rect 148620 660940 148860 661180
rect 148970 660940 149210 661180
rect 149300 660940 149540 661180
rect 149630 660940 149870 661180
rect 149960 660940 150200 661180
rect 150310 660940 150550 661180
rect 150640 660940 150880 661180
rect 150970 660940 151210 661180
rect 151300 660940 151540 661180
rect 151650 660940 151890 661180
rect 151980 660940 152220 661180
rect 152310 660940 152550 661180
rect 152640 660940 152880 661180
rect 152990 660940 153230 661180
rect 153320 660940 153560 661180
rect 153650 660940 153890 661180
rect 153980 660940 154220 661180
rect 154330 660940 154570 661180
rect 154660 660940 154900 661180
rect 154990 660940 155230 661180
rect 155320 660940 155560 661180
rect 155670 660940 155910 661180
rect 110810 660100 111050 660340
rect 111160 660100 111400 660340
rect 111490 660100 111730 660340
rect 111820 660100 112060 660340
rect 112150 660100 112390 660340
rect 112500 660100 112740 660340
rect 112830 660100 113070 660340
rect 113160 660100 113400 660340
rect 113490 660100 113730 660340
rect 113840 660100 114080 660340
rect 114170 660100 114410 660340
rect 114500 660100 114740 660340
rect 114830 660100 115070 660340
rect 115180 660100 115420 660340
rect 115510 660100 115750 660340
rect 115840 660100 116080 660340
rect 116170 660100 116410 660340
rect 116520 660100 116760 660340
rect 116850 660100 117090 660340
rect 117180 660100 117420 660340
rect 117510 660100 117750 660340
rect 117860 660100 118100 660340
rect 118190 660100 118430 660340
rect 118520 660100 118760 660340
rect 118850 660100 119090 660340
rect 119200 660100 119440 660340
rect 119530 660100 119770 660340
rect 119860 660100 120100 660340
rect 120190 660100 120430 660340
rect 120540 660100 120780 660340
rect 120870 660100 121110 660340
rect 121200 660100 121440 660340
rect 121530 660100 121770 660340
rect 110810 659770 111050 660010
rect 111160 659770 111400 660010
rect 111490 659770 111730 660010
rect 111820 659770 112060 660010
rect 112150 659770 112390 660010
rect 112500 659770 112740 660010
rect 112830 659770 113070 660010
rect 113160 659770 113400 660010
rect 113490 659770 113730 660010
rect 113840 659770 114080 660010
rect 114170 659770 114410 660010
rect 114500 659770 114740 660010
rect 114830 659770 115070 660010
rect 115180 659770 115420 660010
rect 115510 659770 115750 660010
rect 115840 659770 116080 660010
rect 116170 659770 116410 660010
rect 116520 659770 116760 660010
rect 116850 659770 117090 660010
rect 117180 659770 117420 660010
rect 117510 659770 117750 660010
rect 117860 659770 118100 660010
rect 118190 659770 118430 660010
rect 118520 659770 118760 660010
rect 118850 659770 119090 660010
rect 119200 659770 119440 660010
rect 119530 659770 119770 660010
rect 119860 659770 120100 660010
rect 120190 659770 120430 660010
rect 120540 659770 120780 660010
rect 120870 659770 121110 660010
rect 121200 659770 121440 660010
rect 121530 659770 121770 660010
rect 110810 659440 111050 659680
rect 111160 659440 111400 659680
rect 111490 659440 111730 659680
rect 111820 659440 112060 659680
rect 112150 659440 112390 659680
rect 112500 659440 112740 659680
rect 112830 659440 113070 659680
rect 113160 659440 113400 659680
rect 113490 659440 113730 659680
rect 113840 659440 114080 659680
rect 114170 659440 114410 659680
rect 114500 659440 114740 659680
rect 114830 659440 115070 659680
rect 115180 659440 115420 659680
rect 115510 659440 115750 659680
rect 115840 659440 116080 659680
rect 116170 659440 116410 659680
rect 116520 659440 116760 659680
rect 116850 659440 117090 659680
rect 117180 659440 117420 659680
rect 117510 659440 117750 659680
rect 117860 659440 118100 659680
rect 118190 659440 118430 659680
rect 118520 659440 118760 659680
rect 118850 659440 119090 659680
rect 119200 659440 119440 659680
rect 119530 659440 119770 659680
rect 119860 659440 120100 659680
rect 120190 659440 120430 659680
rect 120540 659440 120780 659680
rect 120870 659440 121110 659680
rect 121200 659440 121440 659680
rect 121530 659440 121770 659680
rect 110810 659110 111050 659350
rect 111160 659110 111400 659350
rect 111490 659110 111730 659350
rect 111820 659110 112060 659350
rect 112150 659110 112390 659350
rect 112500 659110 112740 659350
rect 112830 659110 113070 659350
rect 113160 659110 113400 659350
rect 113490 659110 113730 659350
rect 113840 659110 114080 659350
rect 114170 659110 114410 659350
rect 114500 659110 114740 659350
rect 114830 659110 115070 659350
rect 115180 659110 115420 659350
rect 115510 659110 115750 659350
rect 115840 659110 116080 659350
rect 116170 659110 116410 659350
rect 116520 659110 116760 659350
rect 116850 659110 117090 659350
rect 117180 659110 117420 659350
rect 117510 659110 117750 659350
rect 117860 659110 118100 659350
rect 118190 659110 118430 659350
rect 118520 659110 118760 659350
rect 118850 659110 119090 659350
rect 119200 659110 119440 659350
rect 119530 659110 119770 659350
rect 119860 659110 120100 659350
rect 120190 659110 120430 659350
rect 120540 659110 120780 659350
rect 120870 659110 121110 659350
rect 121200 659110 121440 659350
rect 121530 659110 121770 659350
rect 110810 658760 111050 659000
rect 111160 658760 111400 659000
rect 111490 658760 111730 659000
rect 111820 658760 112060 659000
rect 112150 658760 112390 659000
rect 112500 658760 112740 659000
rect 112830 658760 113070 659000
rect 113160 658760 113400 659000
rect 113490 658760 113730 659000
rect 113840 658760 114080 659000
rect 114170 658760 114410 659000
rect 114500 658760 114740 659000
rect 114830 658760 115070 659000
rect 115180 658760 115420 659000
rect 115510 658760 115750 659000
rect 115840 658760 116080 659000
rect 116170 658760 116410 659000
rect 116520 658760 116760 659000
rect 116850 658760 117090 659000
rect 117180 658760 117420 659000
rect 117510 658760 117750 659000
rect 117860 658760 118100 659000
rect 118190 658760 118430 659000
rect 118520 658760 118760 659000
rect 118850 658760 119090 659000
rect 119200 658760 119440 659000
rect 119530 658760 119770 659000
rect 119860 658760 120100 659000
rect 120190 658760 120430 659000
rect 120540 658760 120780 659000
rect 120870 658760 121110 659000
rect 121200 658760 121440 659000
rect 121530 658760 121770 659000
rect 110810 658430 111050 658670
rect 111160 658430 111400 658670
rect 111490 658430 111730 658670
rect 111820 658430 112060 658670
rect 112150 658430 112390 658670
rect 112500 658430 112740 658670
rect 112830 658430 113070 658670
rect 113160 658430 113400 658670
rect 113490 658430 113730 658670
rect 113840 658430 114080 658670
rect 114170 658430 114410 658670
rect 114500 658430 114740 658670
rect 114830 658430 115070 658670
rect 115180 658430 115420 658670
rect 115510 658430 115750 658670
rect 115840 658430 116080 658670
rect 116170 658430 116410 658670
rect 116520 658430 116760 658670
rect 116850 658430 117090 658670
rect 117180 658430 117420 658670
rect 117510 658430 117750 658670
rect 117860 658430 118100 658670
rect 118190 658430 118430 658670
rect 118520 658430 118760 658670
rect 118850 658430 119090 658670
rect 119200 658430 119440 658670
rect 119530 658430 119770 658670
rect 119860 658430 120100 658670
rect 120190 658430 120430 658670
rect 120540 658430 120780 658670
rect 120870 658430 121110 658670
rect 121200 658430 121440 658670
rect 121530 658430 121770 658670
rect 110810 658100 111050 658340
rect 111160 658100 111400 658340
rect 111490 658100 111730 658340
rect 111820 658100 112060 658340
rect 112150 658100 112390 658340
rect 112500 658100 112740 658340
rect 112830 658100 113070 658340
rect 113160 658100 113400 658340
rect 113490 658100 113730 658340
rect 113840 658100 114080 658340
rect 114170 658100 114410 658340
rect 114500 658100 114740 658340
rect 114830 658100 115070 658340
rect 115180 658100 115420 658340
rect 115510 658100 115750 658340
rect 115840 658100 116080 658340
rect 116170 658100 116410 658340
rect 116520 658100 116760 658340
rect 116850 658100 117090 658340
rect 117180 658100 117420 658340
rect 117510 658100 117750 658340
rect 117860 658100 118100 658340
rect 118190 658100 118430 658340
rect 118520 658100 118760 658340
rect 118850 658100 119090 658340
rect 119200 658100 119440 658340
rect 119530 658100 119770 658340
rect 119860 658100 120100 658340
rect 120190 658100 120430 658340
rect 120540 658100 120780 658340
rect 120870 658100 121110 658340
rect 121200 658100 121440 658340
rect 121530 658100 121770 658340
rect 110810 657770 111050 658010
rect 111160 657770 111400 658010
rect 111490 657770 111730 658010
rect 111820 657770 112060 658010
rect 112150 657770 112390 658010
rect 112500 657770 112740 658010
rect 112830 657770 113070 658010
rect 113160 657770 113400 658010
rect 113490 657770 113730 658010
rect 113840 657770 114080 658010
rect 114170 657770 114410 658010
rect 114500 657770 114740 658010
rect 114830 657770 115070 658010
rect 115180 657770 115420 658010
rect 115510 657770 115750 658010
rect 115840 657770 116080 658010
rect 116170 657770 116410 658010
rect 116520 657770 116760 658010
rect 116850 657770 117090 658010
rect 117180 657770 117420 658010
rect 117510 657770 117750 658010
rect 117860 657770 118100 658010
rect 118190 657770 118430 658010
rect 118520 657770 118760 658010
rect 118850 657770 119090 658010
rect 119200 657770 119440 658010
rect 119530 657770 119770 658010
rect 119860 657770 120100 658010
rect 120190 657770 120430 658010
rect 120540 657770 120780 658010
rect 120870 657770 121110 658010
rect 121200 657770 121440 658010
rect 121530 657770 121770 658010
rect 110810 657420 111050 657660
rect 111160 657420 111400 657660
rect 111490 657420 111730 657660
rect 111820 657420 112060 657660
rect 112150 657420 112390 657660
rect 112500 657420 112740 657660
rect 112830 657420 113070 657660
rect 113160 657420 113400 657660
rect 113490 657420 113730 657660
rect 113840 657420 114080 657660
rect 114170 657420 114410 657660
rect 114500 657420 114740 657660
rect 114830 657420 115070 657660
rect 115180 657420 115420 657660
rect 115510 657420 115750 657660
rect 115840 657420 116080 657660
rect 116170 657420 116410 657660
rect 116520 657420 116760 657660
rect 116850 657420 117090 657660
rect 117180 657420 117420 657660
rect 117510 657420 117750 657660
rect 117860 657420 118100 657660
rect 118190 657420 118430 657660
rect 118520 657420 118760 657660
rect 118850 657420 119090 657660
rect 119200 657420 119440 657660
rect 119530 657420 119770 657660
rect 119860 657420 120100 657660
rect 120190 657420 120430 657660
rect 120540 657420 120780 657660
rect 120870 657420 121110 657660
rect 121200 657420 121440 657660
rect 121530 657420 121770 657660
rect 110810 657090 111050 657330
rect 111160 657090 111400 657330
rect 111490 657090 111730 657330
rect 111820 657090 112060 657330
rect 112150 657090 112390 657330
rect 112500 657090 112740 657330
rect 112830 657090 113070 657330
rect 113160 657090 113400 657330
rect 113490 657090 113730 657330
rect 113840 657090 114080 657330
rect 114170 657090 114410 657330
rect 114500 657090 114740 657330
rect 114830 657090 115070 657330
rect 115180 657090 115420 657330
rect 115510 657090 115750 657330
rect 115840 657090 116080 657330
rect 116170 657090 116410 657330
rect 116520 657090 116760 657330
rect 116850 657090 117090 657330
rect 117180 657090 117420 657330
rect 117510 657090 117750 657330
rect 117860 657090 118100 657330
rect 118190 657090 118430 657330
rect 118520 657090 118760 657330
rect 118850 657090 119090 657330
rect 119200 657090 119440 657330
rect 119530 657090 119770 657330
rect 119860 657090 120100 657330
rect 120190 657090 120430 657330
rect 120540 657090 120780 657330
rect 120870 657090 121110 657330
rect 121200 657090 121440 657330
rect 121530 657090 121770 657330
rect 110810 656760 111050 657000
rect 111160 656760 111400 657000
rect 111490 656760 111730 657000
rect 111820 656760 112060 657000
rect 112150 656760 112390 657000
rect 112500 656760 112740 657000
rect 112830 656760 113070 657000
rect 113160 656760 113400 657000
rect 113490 656760 113730 657000
rect 113840 656760 114080 657000
rect 114170 656760 114410 657000
rect 114500 656760 114740 657000
rect 114830 656760 115070 657000
rect 115180 656760 115420 657000
rect 115510 656760 115750 657000
rect 115840 656760 116080 657000
rect 116170 656760 116410 657000
rect 116520 656760 116760 657000
rect 116850 656760 117090 657000
rect 117180 656760 117420 657000
rect 117510 656760 117750 657000
rect 117860 656760 118100 657000
rect 118190 656760 118430 657000
rect 118520 656760 118760 657000
rect 118850 656760 119090 657000
rect 119200 656760 119440 657000
rect 119530 656760 119770 657000
rect 119860 656760 120100 657000
rect 120190 656760 120430 657000
rect 120540 656760 120780 657000
rect 120870 656760 121110 657000
rect 121200 656760 121440 657000
rect 121530 656760 121770 657000
rect 110810 656430 111050 656670
rect 111160 656430 111400 656670
rect 111490 656430 111730 656670
rect 111820 656430 112060 656670
rect 112150 656430 112390 656670
rect 112500 656430 112740 656670
rect 112830 656430 113070 656670
rect 113160 656430 113400 656670
rect 113490 656430 113730 656670
rect 113840 656430 114080 656670
rect 114170 656430 114410 656670
rect 114500 656430 114740 656670
rect 114830 656430 115070 656670
rect 115180 656430 115420 656670
rect 115510 656430 115750 656670
rect 115840 656430 116080 656670
rect 116170 656430 116410 656670
rect 116520 656430 116760 656670
rect 116850 656430 117090 656670
rect 117180 656430 117420 656670
rect 117510 656430 117750 656670
rect 117860 656430 118100 656670
rect 118190 656430 118430 656670
rect 118520 656430 118760 656670
rect 118850 656430 119090 656670
rect 119200 656430 119440 656670
rect 119530 656430 119770 656670
rect 119860 656430 120100 656670
rect 120190 656430 120430 656670
rect 120540 656430 120780 656670
rect 120870 656430 121110 656670
rect 121200 656430 121440 656670
rect 121530 656430 121770 656670
rect 110810 656080 111050 656320
rect 111160 656080 111400 656320
rect 111490 656080 111730 656320
rect 111820 656080 112060 656320
rect 112150 656080 112390 656320
rect 112500 656080 112740 656320
rect 112830 656080 113070 656320
rect 113160 656080 113400 656320
rect 113490 656080 113730 656320
rect 113840 656080 114080 656320
rect 114170 656080 114410 656320
rect 114500 656080 114740 656320
rect 114830 656080 115070 656320
rect 115180 656080 115420 656320
rect 115510 656080 115750 656320
rect 115840 656080 116080 656320
rect 116170 656080 116410 656320
rect 116520 656080 116760 656320
rect 116850 656080 117090 656320
rect 117180 656080 117420 656320
rect 117510 656080 117750 656320
rect 117860 656080 118100 656320
rect 118190 656080 118430 656320
rect 118520 656080 118760 656320
rect 118850 656080 119090 656320
rect 119200 656080 119440 656320
rect 119530 656080 119770 656320
rect 119860 656080 120100 656320
rect 120190 656080 120430 656320
rect 120540 656080 120780 656320
rect 120870 656080 121110 656320
rect 121200 656080 121440 656320
rect 121530 656080 121770 656320
rect 110810 655750 111050 655990
rect 111160 655750 111400 655990
rect 111490 655750 111730 655990
rect 111820 655750 112060 655990
rect 112150 655750 112390 655990
rect 112500 655750 112740 655990
rect 112830 655750 113070 655990
rect 113160 655750 113400 655990
rect 113490 655750 113730 655990
rect 113840 655750 114080 655990
rect 114170 655750 114410 655990
rect 114500 655750 114740 655990
rect 114830 655750 115070 655990
rect 115180 655750 115420 655990
rect 115510 655750 115750 655990
rect 115840 655750 116080 655990
rect 116170 655750 116410 655990
rect 116520 655750 116760 655990
rect 116850 655750 117090 655990
rect 117180 655750 117420 655990
rect 117510 655750 117750 655990
rect 117860 655750 118100 655990
rect 118190 655750 118430 655990
rect 118520 655750 118760 655990
rect 118850 655750 119090 655990
rect 119200 655750 119440 655990
rect 119530 655750 119770 655990
rect 119860 655750 120100 655990
rect 120190 655750 120430 655990
rect 120540 655750 120780 655990
rect 120870 655750 121110 655990
rect 121200 655750 121440 655990
rect 121530 655750 121770 655990
rect 110810 655420 111050 655660
rect 111160 655420 111400 655660
rect 111490 655420 111730 655660
rect 111820 655420 112060 655660
rect 112150 655420 112390 655660
rect 112500 655420 112740 655660
rect 112830 655420 113070 655660
rect 113160 655420 113400 655660
rect 113490 655420 113730 655660
rect 113840 655420 114080 655660
rect 114170 655420 114410 655660
rect 114500 655420 114740 655660
rect 114830 655420 115070 655660
rect 115180 655420 115420 655660
rect 115510 655420 115750 655660
rect 115840 655420 116080 655660
rect 116170 655420 116410 655660
rect 116520 655420 116760 655660
rect 116850 655420 117090 655660
rect 117180 655420 117420 655660
rect 117510 655420 117750 655660
rect 117860 655420 118100 655660
rect 118190 655420 118430 655660
rect 118520 655420 118760 655660
rect 118850 655420 119090 655660
rect 119200 655420 119440 655660
rect 119530 655420 119770 655660
rect 119860 655420 120100 655660
rect 120190 655420 120430 655660
rect 120540 655420 120780 655660
rect 120870 655420 121110 655660
rect 121200 655420 121440 655660
rect 121530 655420 121770 655660
rect 110810 655090 111050 655330
rect 111160 655090 111400 655330
rect 111490 655090 111730 655330
rect 111820 655090 112060 655330
rect 112150 655090 112390 655330
rect 112500 655090 112740 655330
rect 112830 655090 113070 655330
rect 113160 655090 113400 655330
rect 113490 655090 113730 655330
rect 113840 655090 114080 655330
rect 114170 655090 114410 655330
rect 114500 655090 114740 655330
rect 114830 655090 115070 655330
rect 115180 655090 115420 655330
rect 115510 655090 115750 655330
rect 115840 655090 116080 655330
rect 116170 655090 116410 655330
rect 116520 655090 116760 655330
rect 116850 655090 117090 655330
rect 117180 655090 117420 655330
rect 117510 655090 117750 655330
rect 117860 655090 118100 655330
rect 118190 655090 118430 655330
rect 118520 655090 118760 655330
rect 118850 655090 119090 655330
rect 119200 655090 119440 655330
rect 119530 655090 119770 655330
rect 119860 655090 120100 655330
rect 120190 655090 120430 655330
rect 120540 655090 120780 655330
rect 120870 655090 121110 655330
rect 121200 655090 121440 655330
rect 121530 655090 121770 655330
rect 110810 654740 111050 654980
rect 111160 654740 111400 654980
rect 111490 654740 111730 654980
rect 111820 654740 112060 654980
rect 112150 654740 112390 654980
rect 112500 654740 112740 654980
rect 112830 654740 113070 654980
rect 113160 654740 113400 654980
rect 113490 654740 113730 654980
rect 113840 654740 114080 654980
rect 114170 654740 114410 654980
rect 114500 654740 114740 654980
rect 114830 654740 115070 654980
rect 115180 654740 115420 654980
rect 115510 654740 115750 654980
rect 115840 654740 116080 654980
rect 116170 654740 116410 654980
rect 116520 654740 116760 654980
rect 116850 654740 117090 654980
rect 117180 654740 117420 654980
rect 117510 654740 117750 654980
rect 117860 654740 118100 654980
rect 118190 654740 118430 654980
rect 118520 654740 118760 654980
rect 118850 654740 119090 654980
rect 119200 654740 119440 654980
rect 119530 654740 119770 654980
rect 119860 654740 120100 654980
rect 120190 654740 120430 654980
rect 120540 654740 120780 654980
rect 120870 654740 121110 654980
rect 121200 654740 121440 654980
rect 121530 654740 121770 654980
rect 110810 654410 111050 654650
rect 111160 654410 111400 654650
rect 111490 654410 111730 654650
rect 111820 654410 112060 654650
rect 112150 654410 112390 654650
rect 112500 654410 112740 654650
rect 112830 654410 113070 654650
rect 113160 654410 113400 654650
rect 113490 654410 113730 654650
rect 113840 654410 114080 654650
rect 114170 654410 114410 654650
rect 114500 654410 114740 654650
rect 114830 654410 115070 654650
rect 115180 654410 115420 654650
rect 115510 654410 115750 654650
rect 115840 654410 116080 654650
rect 116170 654410 116410 654650
rect 116520 654410 116760 654650
rect 116850 654410 117090 654650
rect 117180 654410 117420 654650
rect 117510 654410 117750 654650
rect 117860 654410 118100 654650
rect 118190 654410 118430 654650
rect 118520 654410 118760 654650
rect 118850 654410 119090 654650
rect 119200 654410 119440 654650
rect 119530 654410 119770 654650
rect 119860 654410 120100 654650
rect 120190 654410 120430 654650
rect 120540 654410 120780 654650
rect 120870 654410 121110 654650
rect 121200 654410 121440 654650
rect 121530 654410 121770 654650
rect 110810 654080 111050 654320
rect 111160 654080 111400 654320
rect 111490 654080 111730 654320
rect 111820 654080 112060 654320
rect 112150 654080 112390 654320
rect 112500 654080 112740 654320
rect 112830 654080 113070 654320
rect 113160 654080 113400 654320
rect 113490 654080 113730 654320
rect 113840 654080 114080 654320
rect 114170 654080 114410 654320
rect 114500 654080 114740 654320
rect 114830 654080 115070 654320
rect 115180 654080 115420 654320
rect 115510 654080 115750 654320
rect 115840 654080 116080 654320
rect 116170 654080 116410 654320
rect 116520 654080 116760 654320
rect 116850 654080 117090 654320
rect 117180 654080 117420 654320
rect 117510 654080 117750 654320
rect 117860 654080 118100 654320
rect 118190 654080 118430 654320
rect 118520 654080 118760 654320
rect 118850 654080 119090 654320
rect 119200 654080 119440 654320
rect 119530 654080 119770 654320
rect 119860 654080 120100 654320
rect 120190 654080 120430 654320
rect 120540 654080 120780 654320
rect 120870 654080 121110 654320
rect 121200 654080 121440 654320
rect 121530 654080 121770 654320
rect 110810 653750 111050 653990
rect 111160 653750 111400 653990
rect 111490 653750 111730 653990
rect 111820 653750 112060 653990
rect 112150 653750 112390 653990
rect 112500 653750 112740 653990
rect 112830 653750 113070 653990
rect 113160 653750 113400 653990
rect 113490 653750 113730 653990
rect 113840 653750 114080 653990
rect 114170 653750 114410 653990
rect 114500 653750 114740 653990
rect 114830 653750 115070 653990
rect 115180 653750 115420 653990
rect 115510 653750 115750 653990
rect 115840 653750 116080 653990
rect 116170 653750 116410 653990
rect 116520 653750 116760 653990
rect 116850 653750 117090 653990
rect 117180 653750 117420 653990
rect 117510 653750 117750 653990
rect 117860 653750 118100 653990
rect 118190 653750 118430 653990
rect 118520 653750 118760 653990
rect 118850 653750 119090 653990
rect 119200 653750 119440 653990
rect 119530 653750 119770 653990
rect 119860 653750 120100 653990
rect 120190 653750 120430 653990
rect 120540 653750 120780 653990
rect 120870 653750 121110 653990
rect 121200 653750 121440 653990
rect 121530 653750 121770 653990
rect 110810 653400 111050 653640
rect 111160 653400 111400 653640
rect 111490 653400 111730 653640
rect 111820 653400 112060 653640
rect 112150 653400 112390 653640
rect 112500 653400 112740 653640
rect 112830 653400 113070 653640
rect 113160 653400 113400 653640
rect 113490 653400 113730 653640
rect 113840 653400 114080 653640
rect 114170 653400 114410 653640
rect 114500 653400 114740 653640
rect 114830 653400 115070 653640
rect 115180 653400 115420 653640
rect 115510 653400 115750 653640
rect 115840 653400 116080 653640
rect 116170 653400 116410 653640
rect 116520 653400 116760 653640
rect 116850 653400 117090 653640
rect 117180 653400 117420 653640
rect 117510 653400 117750 653640
rect 117860 653400 118100 653640
rect 118190 653400 118430 653640
rect 118520 653400 118760 653640
rect 118850 653400 119090 653640
rect 119200 653400 119440 653640
rect 119530 653400 119770 653640
rect 119860 653400 120100 653640
rect 120190 653400 120430 653640
rect 120540 653400 120780 653640
rect 120870 653400 121110 653640
rect 121200 653400 121440 653640
rect 121530 653400 121770 653640
rect 110810 653070 111050 653310
rect 111160 653070 111400 653310
rect 111490 653070 111730 653310
rect 111820 653070 112060 653310
rect 112150 653070 112390 653310
rect 112500 653070 112740 653310
rect 112830 653070 113070 653310
rect 113160 653070 113400 653310
rect 113490 653070 113730 653310
rect 113840 653070 114080 653310
rect 114170 653070 114410 653310
rect 114500 653070 114740 653310
rect 114830 653070 115070 653310
rect 115180 653070 115420 653310
rect 115510 653070 115750 653310
rect 115840 653070 116080 653310
rect 116170 653070 116410 653310
rect 116520 653070 116760 653310
rect 116850 653070 117090 653310
rect 117180 653070 117420 653310
rect 117510 653070 117750 653310
rect 117860 653070 118100 653310
rect 118190 653070 118430 653310
rect 118520 653070 118760 653310
rect 118850 653070 119090 653310
rect 119200 653070 119440 653310
rect 119530 653070 119770 653310
rect 119860 653070 120100 653310
rect 120190 653070 120430 653310
rect 120540 653070 120780 653310
rect 120870 653070 121110 653310
rect 121200 653070 121440 653310
rect 121530 653070 121770 653310
rect 110810 652740 111050 652980
rect 111160 652740 111400 652980
rect 111490 652740 111730 652980
rect 111820 652740 112060 652980
rect 112150 652740 112390 652980
rect 112500 652740 112740 652980
rect 112830 652740 113070 652980
rect 113160 652740 113400 652980
rect 113490 652740 113730 652980
rect 113840 652740 114080 652980
rect 114170 652740 114410 652980
rect 114500 652740 114740 652980
rect 114830 652740 115070 652980
rect 115180 652740 115420 652980
rect 115510 652740 115750 652980
rect 115840 652740 116080 652980
rect 116170 652740 116410 652980
rect 116520 652740 116760 652980
rect 116850 652740 117090 652980
rect 117180 652740 117420 652980
rect 117510 652740 117750 652980
rect 117860 652740 118100 652980
rect 118190 652740 118430 652980
rect 118520 652740 118760 652980
rect 118850 652740 119090 652980
rect 119200 652740 119440 652980
rect 119530 652740 119770 652980
rect 119860 652740 120100 652980
rect 120190 652740 120430 652980
rect 120540 652740 120780 652980
rect 120870 652740 121110 652980
rect 121200 652740 121440 652980
rect 121530 652740 121770 652980
rect 110810 652410 111050 652650
rect 111160 652410 111400 652650
rect 111490 652410 111730 652650
rect 111820 652410 112060 652650
rect 112150 652410 112390 652650
rect 112500 652410 112740 652650
rect 112830 652410 113070 652650
rect 113160 652410 113400 652650
rect 113490 652410 113730 652650
rect 113840 652410 114080 652650
rect 114170 652410 114410 652650
rect 114500 652410 114740 652650
rect 114830 652410 115070 652650
rect 115180 652410 115420 652650
rect 115510 652410 115750 652650
rect 115840 652410 116080 652650
rect 116170 652410 116410 652650
rect 116520 652410 116760 652650
rect 116850 652410 117090 652650
rect 117180 652410 117420 652650
rect 117510 652410 117750 652650
rect 117860 652410 118100 652650
rect 118190 652410 118430 652650
rect 118520 652410 118760 652650
rect 118850 652410 119090 652650
rect 119200 652410 119440 652650
rect 119530 652410 119770 652650
rect 119860 652410 120100 652650
rect 120190 652410 120430 652650
rect 120540 652410 120780 652650
rect 120870 652410 121110 652650
rect 121200 652410 121440 652650
rect 121530 652410 121770 652650
rect 110810 652060 111050 652300
rect 111160 652060 111400 652300
rect 111490 652060 111730 652300
rect 111820 652060 112060 652300
rect 112150 652060 112390 652300
rect 112500 652060 112740 652300
rect 112830 652060 113070 652300
rect 113160 652060 113400 652300
rect 113490 652060 113730 652300
rect 113840 652060 114080 652300
rect 114170 652060 114410 652300
rect 114500 652060 114740 652300
rect 114830 652060 115070 652300
rect 115180 652060 115420 652300
rect 115510 652060 115750 652300
rect 115840 652060 116080 652300
rect 116170 652060 116410 652300
rect 116520 652060 116760 652300
rect 116850 652060 117090 652300
rect 117180 652060 117420 652300
rect 117510 652060 117750 652300
rect 117860 652060 118100 652300
rect 118190 652060 118430 652300
rect 118520 652060 118760 652300
rect 118850 652060 119090 652300
rect 119200 652060 119440 652300
rect 119530 652060 119770 652300
rect 119860 652060 120100 652300
rect 120190 652060 120430 652300
rect 120540 652060 120780 652300
rect 120870 652060 121110 652300
rect 121200 652060 121440 652300
rect 121530 652060 121770 652300
rect 110810 651730 111050 651970
rect 111160 651730 111400 651970
rect 111490 651730 111730 651970
rect 111820 651730 112060 651970
rect 112150 651730 112390 651970
rect 112500 651730 112740 651970
rect 112830 651730 113070 651970
rect 113160 651730 113400 651970
rect 113490 651730 113730 651970
rect 113840 651730 114080 651970
rect 114170 651730 114410 651970
rect 114500 651730 114740 651970
rect 114830 651730 115070 651970
rect 115180 651730 115420 651970
rect 115510 651730 115750 651970
rect 115840 651730 116080 651970
rect 116170 651730 116410 651970
rect 116520 651730 116760 651970
rect 116850 651730 117090 651970
rect 117180 651730 117420 651970
rect 117510 651730 117750 651970
rect 117860 651730 118100 651970
rect 118190 651730 118430 651970
rect 118520 651730 118760 651970
rect 118850 651730 119090 651970
rect 119200 651730 119440 651970
rect 119530 651730 119770 651970
rect 119860 651730 120100 651970
rect 120190 651730 120430 651970
rect 120540 651730 120780 651970
rect 120870 651730 121110 651970
rect 121200 651730 121440 651970
rect 121530 651730 121770 651970
rect 110810 651400 111050 651640
rect 111160 651400 111400 651640
rect 111490 651400 111730 651640
rect 111820 651400 112060 651640
rect 112150 651400 112390 651640
rect 112500 651400 112740 651640
rect 112830 651400 113070 651640
rect 113160 651400 113400 651640
rect 113490 651400 113730 651640
rect 113840 651400 114080 651640
rect 114170 651400 114410 651640
rect 114500 651400 114740 651640
rect 114830 651400 115070 651640
rect 115180 651400 115420 651640
rect 115510 651400 115750 651640
rect 115840 651400 116080 651640
rect 116170 651400 116410 651640
rect 116520 651400 116760 651640
rect 116850 651400 117090 651640
rect 117180 651400 117420 651640
rect 117510 651400 117750 651640
rect 117860 651400 118100 651640
rect 118190 651400 118430 651640
rect 118520 651400 118760 651640
rect 118850 651400 119090 651640
rect 119200 651400 119440 651640
rect 119530 651400 119770 651640
rect 119860 651400 120100 651640
rect 120190 651400 120430 651640
rect 120540 651400 120780 651640
rect 120870 651400 121110 651640
rect 121200 651400 121440 651640
rect 121530 651400 121770 651640
rect 110810 651070 111050 651310
rect 111160 651070 111400 651310
rect 111490 651070 111730 651310
rect 111820 651070 112060 651310
rect 112150 651070 112390 651310
rect 112500 651070 112740 651310
rect 112830 651070 113070 651310
rect 113160 651070 113400 651310
rect 113490 651070 113730 651310
rect 113840 651070 114080 651310
rect 114170 651070 114410 651310
rect 114500 651070 114740 651310
rect 114830 651070 115070 651310
rect 115180 651070 115420 651310
rect 115510 651070 115750 651310
rect 115840 651070 116080 651310
rect 116170 651070 116410 651310
rect 116520 651070 116760 651310
rect 116850 651070 117090 651310
rect 117180 651070 117420 651310
rect 117510 651070 117750 651310
rect 117860 651070 118100 651310
rect 118190 651070 118430 651310
rect 118520 651070 118760 651310
rect 118850 651070 119090 651310
rect 119200 651070 119440 651310
rect 119530 651070 119770 651310
rect 119860 651070 120100 651310
rect 120190 651070 120430 651310
rect 120540 651070 120780 651310
rect 120870 651070 121110 651310
rect 121200 651070 121440 651310
rect 121530 651070 121770 651310
rect 110810 650720 111050 650960
rect 111160 650720 111400 650960
rect 111490 650720 111730 650960
rect 111820 650720 112060 650960
rect 112150 650720 112390 650960
rect 112500 650720 112740 650960
rect 112830 650720 113070 650960
rect 113160 650720 113400 650960
rect 113490 650720 113730 650960
rect 113840 650720 114080 650960
rect 114170 650720 114410 650960
rect 114500 650720 114740 650960
rect 114830 650720 115070 650960
rect 115180 650720 115420 650960
rect 115510 650720 115750 650960
rect 115840 650720 116080 650960
rect 116170 650720 116410 650960
rect 116520 650720 116760 650960
rect 116850 650720 117090 650960
rect 117180 650720 117420 650960
rect 117510 650720 117750 650960
rect 117860 650720 118100 650960
rect 118190 650720 118430 650960
rect 118520 650720 118760 650960
rect 118850 650720 119090 650960
rect 119200 650720 119440 650960
rect 119530 650720 119770 650960
rect 119860 650720 120100 650960
rect 120190 650720 120430 650960
rect 120540 650720 120780 650960
rect 120870 650720 121110 650960
rect 121200 650720 121440 650960
rect 121530 650720 121770 650960
rect 110810 650390 111050 650630
rect 111160 650390 111400 650630
rect 111490 650390 111730 650630
rect 111820 650390 112060 650630
rect 112150 650390 112390 650630
rect 112500 650390 112740 650630
rect 112830 650390 113070 650630
rect 113160 650390 113400 650630
rect 113490 650390 113730 650630
rect 113840 650390 114080 650630
rect 114170 650390 114410 650630
rect 114500 650390 114740 650630
rect 114830 650390 115070 650630
rect 115180 650390 115420 650630
rect 115510 650390 115750 650630
rect 115840 650390 116080 650630
rect 116170 650390 116410 650630
rect 116520 650390 116760 650630
rect 116850 650390 117090 650630
rect 117180 650390 117420 650630
rect 117510 650390 117750 650630
rect 117860 650390 118100 650630
rect 118190 650390 118430 650630
rect 118520 650390 118760 650630
rect 118850 650390 119090 650630
rect 119200 650390 119440 650630
rect 119530 650390 119770 650630
rect 119860 650390 120100 650630
rect 120190 650390 120430 650630
rect 120540 650390 120780 650630
rect 120870 650390 121110 650630
rect 121200 650390 121440 650630
rect 121530 650390 121770 650630
rect 110810 650060 111050 650300
rect 111160 650060 111400 650300
rect 111490 650060 111730 650300
rect 111820 650060 112060 650300
rect 112150 650060 112390 650300
rect 112500 650060 112740 650300
rect 112830 650060 113070 650300
rect 113160 650060 113400 650300
rect 113490 650060 113730 650300
rect 113840 650060 114080 650300
rect 114170 650060 114410 650300
rect 114500 650060 114740 650300
rect 114830 650060 115070 650300
rect 115180 650060 115420 650300
rect 115510 650060 115750 650300
rect 115840 650060 116080 650300
rect 116170 650060 116410 650300
rect 116520 650060 116760 650300
rect 116850 650060 117090 650300
rect 117180 650060 117420 650300
rect 117510 650060 117750 650300
rect 117860 650060 118100 650300
rect 118190 650060 118430 650300
rect 118520 650060 118760 650300
rect 118850 650060 119090 650300
rect 119200 650060 119440 650300
rect 119530 650060 119770 650300
rect 119860 650060 120100 650300
rect 120190 650060 120430 650300
rect 120540 650060 120780 650300
rect 120870 650060 121110 650300
rect 121200 650060 121440 650300
rect 121530 650060 121770 650300
rect 110810 649730 111050 649970
rect 111160 649730 111400 649970
rect 111490 649730 111730 649970
rect 111820 649730 112060 649970
rect 112150 649730 112390 649970
rect 112500 649730 112740 649970
rect 112830 649730 113070 649970
rect 113160 649730 113400 649970
rect 113490 649730 113730 649970
rect 113840 649730 114080 649970
rect 114170 649730 114410 649970
rect 114500 649730 114740 649970
rect 114830 649730 115070 649970
rect 115180 649730 115420 649970
rect 115510 649730 115750 649970
rect 115840 649730 116080 649970
rect 116170 649730 116410 649970
rect 116520 649730 116760 649970
rect 116850 649730 117090 649970
rect 117180 649730 117420 649970
rect 117510 649730 117750 649970
rect 117860 649730 118100 649970
rect 118190 649730 118430 649970
rect 118520 649730 118760 649970
rect 118850 649730 119090 649970
rect 119200 649730 119440 649970
rect 119530 649730 119770 649970
rect 119860 649730 120100 649970
rect 120190 649730 120430 649970
rect 120540 649730 120780 649970
rect 120870 649730 121110 649970
rect 121200 649730 121440 649970
rect 121530 649730 121770 649970
rect 110810 649380 111050 649620
rect 111160 649380 111400 649620
rect 111490 649380 111730 649620
rect 111820 649380 112060 649620
rect 112150 649380 112390 649620
rect 112500 649380 112740 649620
rect 112830 649380 113070 649620
rect 113160 649380 113400 649620
rect 113490 649380 113730 649620
rect 113840 649380 114080 649620
rect 114170 649380 114410 649620
rect 114500 649380 114740 649620
rect 114830 649380 115070 649620
rect 115180 649380 115420 649620
rect 115510 649380 115750 649620
rect 115840 649380 116080 649620
rect 116170 649380 116410 649620
rect 116520 649380 116760 649620
rect 116850 649380 117090 649620
rect 117180 649380 117420 649620
rect 117510 649380 117750 649620
rect 117860 649380 118100 649620
rect 118190 649380 118430 649620
rect 118520 649380 118760 649620
rect 118850 649380 119090 649620
rect 119200 649380 119440 649620
rect 119530 649380 119770 649620
rect 119860 649380 120100 649620
rect 120190 649380 120430 649620
rect 120540 649380 120780 649620
rect 120870 649380 121110 649620
rect 121200 649380 121440 649620
rect 121530 649380 121770 649620
rect 122190 660100 122430 660340
rect 122540 660100 122780 660340
rect 122870 660100 123110 660340
rect 123200 660100 123440 660340
rect 123530 660100 123770 660340
rect 123880 660100 124120 660340
rect 124210 660100 124450 660340
rect 124540 660100 124780 660340
rect 124870 660100 125110 660340
rect 125220 660100 125460 660340
rect 125550 660100 125790 660340
rect 125880 660100 126120 660340
rect 126210 660100 126450 660340
rect 126560 660100 126800 660340
rect 126890 660100 127130 660340
rect 127220 660100 127460 660340
rect 127550 660100 127790 660340
rect 127900 660100 128140 660340
rect 128230 660100 128470 660340
rect 128560 660100 128800 660340
rect 128890 660100 129130 660340
rect 129240 660100 129480 660340
rect 129570 660100 129810 660340
rect 129900 660100 130140 660340
rect 130230 660100 130470 660340
rect 130580 660100 130820 660340
rect 130910 660100 131150 660340
rect 131240 660100 131480 660340
rect 131570 660100 131810 660340
rect 131920 660100 132160 660340
rect 132250 660100 132490 660340
rect 132580 660100 132820 660340
rect 132910 660100 133150 660340
rect 122190 659770 122430 660010
rect 122540 659770 122780 660010
rect 122870 659770 123110 660010
rect 123200 659770 123440 660010
rect 123530 659770 123770 660010
rect 123880 659770 124120 660010
rect 124210 659770 124450 660010
rect 124540 659770 124780 660010
rect 124870 659770 125110 660010
rect 125220 659770 125460 660010
rect 125550 659770 125790 660010
rect 125880 659770 126120 660010
rect 126210 659770 126450 660010
rect 126560 659770 126800 660010
rect 126890 659770 127130 660010
rect 127220 659770 127460 660010
rect 127550 659770 127790 660010
rect 127900 659770 128140 660010
rect 128230 659770 128470 660010
rect 128560 659770 128800 660010
rect 128890 659770 129130 660010
rect 129240 659770 129480 660010
rect 129570 659770 129810 660010
rect 129900 659770 130140 660010
rect 130230 659770 130470 660010
rect 130580 659770 130820 660010
rect 130910 659770 131150 660010
rect 131240 659770 131480 660010
rect 131570 659770 131810 660010
rect 131920 659770 132160 660010
rect 132250 659770 132490 660010
rect 132580 659770 132820 660010
rect 132910 659770 133150 660010
rect 122190 659440 122430 659680
rect 122540 659440 122780 659680
rect 122870 659440 123110 659680
rect 123200 659440 123440 659680
rect 123530 659440 123770 659680
rect 123880 659440 124120 659680
rect 124210 659440 124450 659680
rect 124540 659440 124780 659680
rect 124870 659440 125110 659680
rect 125220 659440 125460 659680
rect 125550 659440 125790 659680
rect 125880 659440 126120 659680
rect 126210 659440 126450 659680
rect 126560 659440 126800 659680
rect 126890 659440 127130 659680
rect 127220 659440 127460 659680
rect 127550 659440 127790 659680
rect 127900 659440 128140 659680
rect 128230 659440 128470 659680
rect 128560 659440 128800 659680
rect 128890 659440 129130 659680
rect 129240 659440 129480 659680
rect 129570 659440 129810 659680
rect 129900 659440 130140 659680
rect 130230 659440 130470 659680
rect 130580 659440 130820 659680
rect 130910 659440 131150 659680
rect 131240 659440 131480 659680
rect 131570 659440 131810 659680
rect 131920 659440 132160 659680
rect 132250 659440 132490 659680
rect 132580 659440 132820 659680
rect 132910 659440 133150 659680
rect 122190 659110 122430 659350
rect 122540 659110 122780 659350
rect 122870 659110 123110 659350
rect 123200 659110 123440 659350
rect 123530 659110 123770 659350
rect 123880 659110 124120 659350
rect 124210 659110 124450 659350
rect 124540 659110 124780 659350
rect 124870 659110 125110 659350
rect 125220 659110 125460 659350
rect 125550 659110 125790 659350
rect 125880 659110 126120 659350
rect 126210 659110 126450 659350
rect 126560 659110 126800 659350
rect 126890 659110 127130 659350
rect 127220 659110 127460 659350
rect 127550 659110 127790 659350
rect 127900 659110 128140 659350
rect 128230 659110 128470 659350
rect 128560 659110 128800 659350
rect 128890 659110 129130 659350
rect 129240 659110 129480 659350
rect 129570 659110 129810 659350
rect 129900 659110 130140 659350
rect 130230 659110 130470 659350
rect 130580 659110 130820 659350
rect 130910 659110 131150 659350
rect 131240 659110 131480 659350
rect 131570 659110 131810 659350
rect 131920 659110 132160 659350
rect 132250 659110 132490 659350
rect 132580 659110 132820 659350
rect 132910 659110 133150 659350
rect 122190 658760 122430 659000
rect 122540 658760 122780 659000
rect 122870 658760 123110 659000
rect 123200 658760 123440 659000
rect 123530 658760 123770 659000
rect 123880 658760 124120 659000
rect 124210 658760 124450 659000
rect 124540 658760 124780 659000
rect 124870 658760 125110 659000
rect 125220 658760 125460 659000
rect 125550 658760 125790 659000
rect 125880 658760 126120 659000
rect 126210 658760 126450 659000
rect 126560 658760 126800 659000
rect 126890 658760 127130 659000
rect 127220 658760 127460 659000
rect 127550 658760 127790 659000
rect 127900 658760 128140 659000
rect 128230 658760 128470 659000
rect 128560 658760 128800 659000
rect 128890 658760 129130 659000
rect 129240 658760 129480 659000
rect 129570 658760 129810 659000
rect 129900 658760 130140 659000
rect 130230 658760 130470 659000
rect 130580 658760 130820 659000
rect 130910 658760 131150 659000
rect 131240 658760 131480 659000
rect 131570 658760 131810 659000
rect 131920 658760 132160 659000
rect 132250 658760 132490 659000
rect 132580 658760 132820 659000
rect 132910 658760 133150 659000
rect 122190 658430 122430 658670
rect 122540 658430 122780 658670
rect 122870 658430 123110 658670
rect 123200 658430 123440 658670
rect 123530 658430 123770 658670
rect 123880 658430 124120 658670
rect 124210 658430 124450 658670
rect 124540 658430 124780 658670
rect 124870 658430 125110 658670
rect 125220 658430 125460 658670
rect 125550 658430 125790 658670
rect 125880 658430 126120 658670
rect 126210 658430 126450 658670
rect 126560 658430 126800 658670
rect 126890 658430 127130 658670
rect 127220 658430 127460 658670
rect 127550 658430 127790 658670
rect 127900 658430 128140 658670
rect 128230 658430 128470 658670
rect 128560 658430 128800 658670
rect 128890 658430 129130 658670
rect 129240 658430 129480 658670
rect 129570 658430 129810 658670
rect 129900 658430 130140 658670
rect 130230 658430 130470 658670
rect 130580 658430 130820 658670
rect 130910 658430 131150 658670
rect 131240 658430 131480 658670
rect 131570 658430 131810 658670
rect 131920 658430 132160 658670
rect 132250 658430 132490 658670
rect 132580 658430 132820 658670
rect 132910 658430 133150 658670
rect 122190 658100 122430 658340
rect 122540 658100 122780 658340
rect 122870 658100 123110 658340
rect 123200 658100 123440 658340
rect 123530 658100 123770 658340
rect 123880 658100 124120 658340
rect 124210 658100 124450 658340
rect 124540 658100 124780 658340
rect 124870 658100 125110 658340
rect 125220 658100 125460 658340
rect 125550 658100 125790 658340
rect 125880 658100 126120 658340
rect 126210 658100 126450 658340
rect 126560 658100 126800 658340
rect 126890 658100 127130 658340
rect 127220 658100 127460 658340
rect 127550 658100 127790 658340
rect 127900 658100 128140 658340
rect 128230 658100 128470 658340
rect 128560 658100 128800 658340
rect 128890 658100 129130 658340
rect 129240 658100 129480 658340
rect 129570 658100 129810 658340
rect 129900 658100 130140 658340
rect 130230 658100 130470 658340
rect 130580 658100 130820 658340
rect 130910 658100 131150 658340
rect 131240 658100 131480 658340
rect 131570 658100 131810 658340
rect 131920 658100 132160 658340
rect 132250 658100 132490 658340
rect 132580 658100 132820 658340
rect 132910 658100 133150 658340
rect 122190 657770 122430 658010
rect 122540 657770 122780 658010
rect 122870 657770 123110 658010
rect 123200 657770 123440 658010
rect 123530 657770 123770 658010
rect 123880 657770 124120 658010
rect 124210 657770 124450 658010
rect 124540 657770 124780 658010
rect 124870 657770 125110 658010
rect 125220 657770 125460 658010
rect 125550 657770 125790 658010
rect 125880 657770 126120 658010
rect 126210 657770 126450 658010
rect 126560 657770 126800 658010
rect 126890 657770 127130 658010
rect 127220 657770 127460 658010
rect 127550 657770 127790 658010
rect 127900 657770 128140 658010
rect 128230 657770 128470 658010
rect 128560 657770 128800 658010
rect 128890 657770 129130 658010
rect 129240 657770 129480 658010
rect 129570 657770 129810 658010
rect 129900 657770 130140 658010
rect 130230 657770 130470 658010
rect 130580 657770 130820 658010
rect 130910 657770 131150 658010
rect 131240 657770 131480 658010
rect 131570 657770 131810 658010
rect 131920 657770 132160 658010
rect 132250 657770 132490 658010
rect 132580 657770 132820 658010
rect 132910 657770 133150 658010
rect 122190 657420 122430 657660
rect 122540 657420 122780 657660
rect 122870 657420 123110 657660
rect 123200 657420 123440 657660
rect 123530 657420 123770 657660
rect 123880 657420 124120 657660
rect 124210 657420 124450 657660
rect 124540 657420 124780 657660
rect 124870 657420 125110 657660
rect 125220 657420 125460 657660
rect 125550 657420 125790 657660
rect 125880 657420 126120 657660
rect 126210 657420 126450 657660
rect 126560 657420 126800 657660
rect 126890 657420 127130 657660
rect 127220 657420 127460 657660
rect 127550 657420 127790 657660
rect 127900 657420 128140 657660
rect 128230 657420 128470 657660
rect 128560 657420 128800 657660
rect 128890 657420 129130 657660
rect 129240 657420 129480 657660
rect 129570 657420 129810 657660
rect 129900 657420 130140 657660
rect 130230 657420 130470 657660
rect 130580 657420 130820 657660
rect 130910 657420 131150 657660
rect 131240 657420 131480 657660
rect 131570 657420 131810 657660
rect 131920 657420 132160 657660
rect 132250 657420 132490 657660
rect 132580 657420 132820 657660
rect 132910 657420 133150 657660
rect 122190 657090 122430 657330
rect 122540 657090 122780 657330
rect 122870 657090 123110 657330
rect 123200 657090 123440 657330
rect 123530 657090 123770 657330
rect 123880 657090 124120 657330
rect 124210 657090 124450 657330
rect 124540 657090 124780 657330
rect 124870 657090 125110 657330
rect 125220 657090 125460 657330
rect 125550 657090 125790 657330
rect 125880 657090 126120 657330
rect 126210 657090 126450 657330
rect 126560 657090 126800 657330
rect 126890 657090 127130 657330
rect 127220 657090 127460 657330
rect 127550 657090 127790 657330
rect 127900 657090 128140 657330
rect 128230 657090 128470 657330
rect 128560 657090 128800 657330
rect 128890 657090 129130 657330
rect 129240 657090 129480 657330
rect 129570 657090 129810 657330
rect 129900 657090 130140 657330
rect 130230 657090 130470 657330
rect 130580 657090 130820 657330
rect 130910 657090 131150 657330
rect 131240 657090 131480 657330
rect 131570 657090 131810 657330
rect 131920 657090 132160 657330
rect 132250 657090 132490 657330
rect 132580 657090 132820 657330
rect 132910 657090 133150 657330
rect 122190 656760 122430 657000
rect 122540 656760 122780 657000
rect 122870 656760 123110 657000
rect 123200 656760 123440 657000
rect 123530 656760 123770 657000
rect 123880 656760 124120 657000
rect 124210 656760 124450 657000
rect 124540 656760 124780 657000
rect 124870 656760 125110 657000
rect 125220 656760 125460 657000
rect 125550 656760 125790 657000
rect 125880 656760 126120 657000
rect 126210 656760 126450 657000
rect 126560 656760 126800 657000
rect 126890 656760 127130 657000
rect 127220 656760 127460 657000
rect 127550 656760 127790 657000
rect 127900 656760 128140 657000
rect 128230 656760 128470 657000
rect 128560 656760 128800 657000
rect 128890 656760 129130 657000
rect 129240 656760 129480 657000
rect 129570 656760 129810 657000
rect 129900 656760 130140 657000
rect 130230 656760 130470 657000
rect 130580 656760 130820 657000
rect 130910 656760 131150 657000
rect 131240 656760 131480 657000
rect 131570 656760 131810 657000
rect 131920 656760 132160 657000
rect 132250 656760 132490 657000
rect 132580 656760 132820 657000
rect 132910 656760 133150 657000
rect 122190 656430 122430 656670
rect 122540 656430 122780 656670
rect 122870 656430 123110 656670
rect 123200 656430 123440 656670
rect 123530 656430 123770 656670
rect 123880 656430 124120 656670
rect 124210 656430 124450 656670
rect 124540 656430 124780 656670
rect 124870 656430 125110 656670
rect 125220 656430 125460 656670
rect 125550 656430 125790 656670
rect 125880 656430 126120 656670
rect 126210 656430 126450 656670
rect 126560 656430 126800 656670
rect 126890 656430 127130 656670
rect 127220 656430 127460 656670
rect 127550 656430 127790 656670
rect 127900 656430 128140 656670
rect 128230 656430 128470 656670
rect 128560 656430 128800 656670
rect 128890 656430 129130 656670
rect 129240 656430 129480 656670
rect 129570 656430 129810 656670
rect 129900 656430 130140 656670
rect 130230 656430 130470 656670
rect 130580 656430 130820 656670
rect 130910 656430 131150 656670
rect 131240 656430 131480 656670
rect 131570 656430 131810 656670
rect 131920 656430 132160 656670
rect 132250 656430 132490 656670
rect 132580 656430 132820 656670
rect 132910 656430 133150 656670
rect 122190 656080 122430 656320
rect 122540 656080 122780 656320
rect 122870 656080 123110 656320
rect 123200 656080 123440 656320
rect 123530 656080 123770 656320
rect 123880 656080 124120 656320
rect 124210 656080 124450 656320
rect 124540 656080 124780 656320
rect 124870 656080 125110 656320
rect 125220 656080 125460 656320
rect 125550 656080 125790 656320
rect 125880 656080 126120 656320
rect 126210 656080 126450 656320
rect 126560 656080 126800 656320
rect 126890 656080 127130 656320
rect 127220 656080 127460 656320
rect 127550 656080 127790 656320
rect 127900 656080 128140 656320
rect 128230 656080 128470 656320
rect 128560 656080 128800 656320
rect 128890 656080 129130 656320
rect 129240 656080 129480 656320
rect 129570 656080 129810 656320
rect 129900 656080 130140 656320
rect 130230 656080 130470 656320
rect 130580 656080 130820 656320
rect 130910 656080 131150 656320
rect 131240 656080 131480 656320
rect 131570 656080 131810 656320
rect 131920 656080 132160 656320
rect 132250 656080 132490 656320
rect 132580 656080 132820 656320
rect 132910 656080 133150 656320
rect 122190 655750 122430 655990
rect 122540 655750 122780 655990
rect 122870 655750 123110 655990
rect 123200 655750 123440 655990
rect 123530 655750 123770 655990
rect 123880 655750 124120 655990
rect 124210 655750 124450 655990
rect 124540 655750 124780 655990
rect 124870 655750 125110 655990
rect 125220 655750 125460 655990
rect 125550 655750 125790 655990
rect 125880 655750 126120 655990
rect 126210 655750 126450 655990
rect 126560 655750 126800 655990
rect 126890 655750 127130 655990
rect 127220 655750 127460 655990
rect 127550 655750 127790 655990
rect 127900 655750 128140 655990
rect 128230 655750 128470 655990
rect 128560 655750 128800 655990
rect 128890 655750 129130 655990
rect 129240 655750 129480 655990
rect 129570 655750 129810 655990
rect 129900 655750 130140 655990
rect 130230 655750 130470 655990
rect 130580 655750 130820 655990
rect 130910 655750 131150 655990
rect 131240 655750 131480 655990
rect 131570 655750 131810 655990
rect 131920 655750 132160 655990
rect 132250 655750 132490 655990
rect 132580 655750 132820 655990
rect 132910 655750 133150 655990
rect 122190 655420 122430 655660
rect 122540 655420 122780 655660
rect 122870 655420 123110 655660
rect 123200 655420 123440 655660
rect 123530 655420 123770 655660
rect 123880 655420 124120 655660
rect 124210 655420 124450 655660
rect 124540 655420 124780 655660
rect 124870 655420 125110 655660
rect 125220 655420 125460 655660
rect 125550 655420 125790 655660
rect 125880 655420 126120 655660
rect 126210 655420 126450 655660
rect 126560 655420 126800 655660
rect 126890 655420 127130 655660
rect 127220 655420 127460 655660
rect 127550 655420 127790 655660
rect 127900 655420 128140 655660
rect 128230 655420 128470 655660
rect 128560 655420 128800 655660
rect 128890 655420 129130 655660
rect 129240 655420 129480 655660
rect 129570 655420 129810 655660
rect 129900 655420 130140 655660
rect 130230 655420 130470 655660
rect 130580 655420 130820 655660
rect 130910 655420 131150 655660
rect 131240 655420 131480 655660
rect 131570 655420 131810 655660
rect 131920 655420 132160 655660
rect 132250 655420 132490 655660
rect 132580 655420 132820 655660
rect 132910 655420 133150 655660
rect 122190 655090 122430 655330
rect 122540 655090 122780 655330
rect 122870 655090 123110 655330
rect 123200 655090 123440 655330
rect 123530 655090 123770 655330
rect 123880 655090 124120 655330
rect 124210 655090 124450 655330
rect 124540 655090 124780 655330
rect 124870 655090 125110 655330
rect 125220 655090 125460 655330
rect 125550 655090 125790 655330
rect 125880 655090 126120 655330
rect 126210 655090 126450 655330
rect 126560 655090 126800 655330
rect 126890 655090 127130 655330
rect 127220 655090 127460 655330
rect 127550 655090 127790 655330
rect 127900 655090 128140 655330
rect 128230 655090 128470 655330
rect 128560 655090 128800 655330
rect 128890 655090 129130 655330
rect 129240 655090 129480 655330
rect 129570 655090 129810 655330
rect 129900 655090 130140 655330
rect 130230 655090 130470 655330
rect 130580 655090 130820 655330
rect 130910 655090 131150 655330
rect 131240 655090 131480 655330
rect 131570 655090 131810 655330
rect 131920 655090 132160 655330
rect 132250 655090 132490 655330
rect 132580 655090 132820 655330
rect 132910 655090 133150 655330
rect 122190 654740 122430 654980
rect 122540 654740 122780 654980
rect 122870 654740 123110 654980
rect 123200 654740 123440 654980
rect 123530 654740 123770 654980
rect 123880 654740 124120 654980
rect 124210 654740 124450 654980
rect 124540 654740 124780 654980
rect 124870 654740 125110 654980
rect 125220 654740 125460 654980
rect 125550 654740 125790 654980
rect 125880 654740 126120 654980
rect 126210 654740 126450 654980
rect 126560 654740 126800 654980
rect 126890 654740 127130 654980
rect 127220 654740 127460 654980
rect 127550 654740 127790 654980
rect 127900 654740 128140 654980
rect 128230 654740 128470 654980
rect 128560 654740 128800 654980
rect 128890 654740 129130 654980
rect 129240 654740 129480 654980
rect 129570 654740 129810 654980
rect 129900 654740 130140 654980
rect 130230 654740 130470 654980
rect 130580 654740 130820 654980
rect 130910 654740 131150 654980
rect 131240 654740 131480 654980
rect 131570 654740 131810 654980
rect 131920 654740 132160 654980
rect 132250 654740 132490 654980
rect 132580 654740 132820 654980
rect 132910 654740 133150 654980
rect 122190 654410 122430 654650
rect 122540 654410 122780 654650
rect 122870 654410 123110 654650
rect 123200 654410 123440 654650
rect 123530 654410 123770 654650
rect 123880 654410 124120 654650
rect 124210 654410 124450 654650
rect 124540 654410 124780 654650
rect 124870 654410 125110 654650
rect 125220 654410 125460 654650
rect 125550 654410 125790 654650
rect 125880 654410 126120 654650
rect 126210 654410 126450 654650
rect 126560 654410 126800 654650
rect 126890 654410 127130 654650
rect 127220 654410 127460 654650
rect 127550 654410 127790 654650
rect 127900 654410 128140 654650
rect 128230 654410 128470 654650
rect 128560 654410 128800 654650
rect 128890 654410 129130 654650
rect 129240 654410 129480 654650
rect 129570 654410 129810 654650
rect 129900 654410 130140 654650
rect 130230 654410 130470 654650
rect 130580 654410 130820 654650
rect 130910 654410 131150 654650
rect 131240 654410 131480 654650
rect 131570 654410 131810 654650
rect 131920 654410 132160 654650
rect 132250 654410 132490 654650
rect 132580 654410 132820 654650
rect 132910 654410 133150 654650
rect 122190 654080 122430 654320
rect 122540 654080 122780 654320
rect 122870 654080 123110 654320
rect 123200 654080 123440 654320
rect 123530 654080 123770 654320
rect 123880 654080 124120 654320
rect 124210 654080 124450 654320
rect 124540 654080 124780 654320
rect 124870 654080 125110 654320
rect 125220 654080 125460 654320
rect 125550 654080 125790 654320
rect 125880 654080 126120 654320
rect 126210 654080 126450 654320
rect 126560 654080 126800 654320
rect 126890 654080 127130 654320
rect 127220 654080 127460 654320
rect 127550 654080 127790 654320
rect 127900 654080 128140 654320
rect 128230 654080 128470 654320
rect 128560 654080 128800 654320
rect 128890 654080 129130 654320
rect 129240 654080 129480 654320
rect 129570 654080 129810 654320
rect 129900 654080 130140 654320
rect 130230 654080 130470 654320
rect 130580 654080 130820 654320
rect 130910 654080 131150 654320
rect 131240 654080 131480 654320
rect 131570 654080 131810 654320
rect 131920 654080 132160 654320
rect 132250 654080 132490 654320
rect 132580 654080 132820 654320
rect 132910 654080 133150 654320
rect 122190 653750 122430 653990
rect 122540 653750 122780 653990
rect 122870 653750 123110 653990
rect 123200 653750 123440 653990
rect 123530 653750 123770 653990
rect 123880 653750 124120 653990
rect 124210 653750 124450 653990
rect 124540 653750 124780 653990
rect 124870 653750 125110 653990
rect 125220 653750 125460 653990
rect 125550 653750 125790 653990
rect 125880 653750 126120 653990
rect 126210 653750 126450 653990
rect 126560 653750 126800 653990
rect 126890 653750 127130 653990
rect 127220 653750 127460 653990
rect 127550 653750 127790 653990
rect 127900 653750 128140 653990
rect 128230 653750 128470 653990
rect 128560 653750 128800 653990
rect 128890 653750 129130 653990
rect 129240 653750 129480 653990
rect 129570 653750 129810 653990
rect 129900 653750 130140 653990
rect 130230 653750 130470 653990
rect 130580 653750 130820 653990
rect 130910 653750 131150 653990
rect 131240 653750 131480 653990
rect 131570 653750 131810 653990
rect 131920 653750 132160 653990
rect 132250 653750 132490 653990
rect 132580 653750 132820 653990
rect 132910 653750 133150 653990
rect 122190 653400 122430 653640
rect 122540 653400 122780 653640
rect 122870 653400 123110 653640
rect 123200 653400 123440 653640
rect 123530 653400 123770 653640
rect 123880 653400 124120 653640
rect 124210 653400 124450 653640
rect 124540 653400 124780 653640
rect 124870 653400 125110 653640
rect 125220 653400 125460 653640
rect 125550 653400 125790 653640
rect 125880 653400 126120 653640
rect 126210 653400 126450 653640
rect 126560 653400 126800 653640
rect 126890 653400 127130 653640
rect 127220 653400 127460 653640
rect 127550 653400 127790 653640
rect 127900 653400 128140 653640
rect 128230 653400 128470 653640
rect 128560 653400 128800 653640
rect 128890 653400 129130 653640
rect 129240 653400 129480 653640
rect 129570 653400 129810 653640
rect 129900 653400 130140 653640
rect 130230 653400 130470 653640
rect 130580 653400 130820 653640
rect 130910 653400 131150 653640
rect 131240 653400 131480 653640
rect 131570 653400 131810 653640
rect 131920 653400 132160 653640
rect 132250 653400 132490 653640
rect 132580 653400 132820 653640
rect 132910 653400 133150 653640
rect 122190 653070 122430 653310
rect 122540 653070 122780 653310
rect 122870 653070 123110 653310
rect 123200 653070 123440 653310
rect 123530 653070 123770 653310
rect 123880 653070 124120 653310
rect 124210 653070 124450 653310
rect 124540 653070 124780 653310
rect 124870 653070 125110 653310
rect 125220 653070 125460 653310
rect 125550 653070 125790 653310
rect 125880 653070 126120 653310
rect 126210 653070 126450 653310
rect 126560 653070 126800 653310
rect 126890 653070 127130 653310
rect 127220 653070 127460 653310
rect 127550 653070 127790 653310
rect 127900 653070 128140 653310
rect 128230 653070 128470 653310
rect 128560 653070 128800 653310
rect 128890 653070 129130 653310
rect 129240 653070 129480 653310
rect 129570 653070 129810 653310
rect 129900 653070 130140 653310
rect 130230 653070 130470 653310
rect 130580 653070 130820 653310
rect 130910 653070 131150 653310
rect 131240 653070 131480 653310
rect 131570 653070 131810 653310
rect 131920 653070 132160 653310
rect 132250 653070 132490 653310
rect 132580 653070 132820 653310
rect 132910 653070 133150 653310
rect 122190 652740 122430 652980
rect 122540 652740 122780 652980
rect 122870 652740 123110 652980
rect 123200 652740 123440 652980
rect 123530 652740 123770 652980
rect 123880 652740 124120 652980
rect 124210 652740 124450 652980
rect 124540 652740 124780 652980
rect 124870 652740 125110 652980
rect 125220 652740 125460 652980
rect 125550 652740 125790 652980
rect 125880 652740 126120 652980
rect 126210 652740 126450 652980
rect 126560 652740 126800 652980
rect 126890 652740 127130 652980
rect 127220 652740 127460 652980
rect 127550 652740 127790 652980
rect 127900 652740 128140 652980
rect 128230 652740 128470 652980
rect 128560 652740 128800 652980
rect 128890 652740 129130 652980
rect 129240 652740 129480 652980
rect 129570 652740 129810 652980
rect 129900 652740 130140 652980
rect 130230 652740 130470 652980
rect 130580 652740 130820 652980
rect 130910 652740 131150 652980
rect 131240 652740 131480 652980
rect 131570 652740 131810 652980
rect 131920 652740 132160 652980
rect 132250 652740 132490 652980
rect 132580 652740 132820 652980
rect 132910 652740 133150 652980
rect 122190 652410 122430 652650
rect 122540 652410 122780 652650
rect 122870 652410 123110 652650
rect 123200 652410 123440 652650
rect 123530 652410 123770 652650
rect 123880 652410 124120 652650
rect 124210 652410 124450 652650
rect 124540 652410 124780 652650
rect 124870 652410 125110 652650
rect 125220 652410 125460 652650
rect 125550 652410 125790 652650
rect 125880 652410 126120 652650
rect 126210 652410 126450 652650
rect 126560 652410 126800 652650
rect 126890 652410 127130 652650
rect 127220 652410 127460 652650
rect 127550 652410 127790 652650
rect 127900 652410 128140 652650
rect 128230 652410 128470 652650
rect 128560 652410 128800 652650
rect 128890 652410 129130 652650
rect 129240 652410 129480 652650
rect 129570 652410 129810 652650
rect 129900 652410 130140 652650
rect 130230 652410 130470 652650
rect 130580 652410 130820 652650
rect 130910 652410 131150 652650
rect 131240 652410 131480 652650
rect 131570 652410 131810 652650
rect 131920 652410 132160 652650
rect 132250 652410 132490 652650
rect 132580 652410 132820 652650
rect 132910 652410 133150 652650
rect 122190 652060 122430 652300
rect 122540 652060 122780 652300
rect 122870 652060 123110 652300
rect 123200 652060 123440 652300
rect 123530 652060 123770 652300
rect 123880 652060 124120 652300
rect 124210 652060 124450 652300
rect 124540 652060 124780 652300
rect 124870 652060 125110 652300
rect 125220 652060 125460 652300
rect 125550 652060 125790 652300
rect 125880 652060 126120 652300
rect 126210 652060 126450 652300
rect 126560 652060 126800 652300
rect 126890 652060 127130 652300
rect 127220 652060 127460 652300
rect 127550 652060 127790 652300
rect 127900 652060 128140 652300
rect 128230 652060 128470 652300
rect 128560 652060 128800 652300
rect 128890 652060 129130 652300
rect 129240 652060 129480 652300
rect 129570 652060 129810 652300
rect 129900 652060 130140 652300
rect 130230 652060 130470 652300
rect 130580 652060 130820 652300
rect 130910 652060 131150 652300
rect 131240 652060 131480 652300
rect 131570 652060 131810 652300
rect 131920 652060 132160 652300
rect 132250 652060 132490 652300
rect 132580 652060 132820 652300
rect 132910 652060 133150 652300
rect 122190 651730 122430 651970
rect 122540 651730 122780 651970
rect 122870 651730 123110 651970
rect 123200 651730 123440 651970
rect 123530 651730 123770 651970
rect 123880 651730 124120 651970
rect 124210 651730 124450 651970
rect 124540 651730 124780 651970
rect 124870 651730 125110 651970
rect 125220 651730 125460 651970
rect 125550 651730 125790 651970
rect 125880 651730 126120 651970
rect 126210 651730 126450 651970
rect 126560 651730 126800 651970
rect 126890 651730 127130 651970
rect 127220 651730 127460 651970
rect 127550 651730 127790 651970
rect 127900 651730 128140 651970
rect 128230 651730 128470 651970
rect 128560 651730 128800 651970
rect 128890 651730 129130 651970
rect 129240 651730 129480 651970
rect 129570 651730 129810 651970
rect 129900 651730 130140 651970
rect 130230 651730 130470 651970
rect 130580 651730 130820 651970
rect 130910 651730 131150 651970
rect 131240 651730 131480 651970
rect 131570 651730 131810 651970
rect 131920 651730 132160 651970
rect 132250 651730 132490 651970
rect 132580 651730 132820 651970
rect 132910 651730 133150 651970
rect 122190 651400 122430 651640
rect 122540 651400 122780 651640
rect 122870 651400 123110 651640
rect 123200 651400 123440 651640
rect 123530 651400 123770 651640
rect 123880 651400 124120 651640
rect 124210 651400 124450 651640
rect 124540 651400 124780 651640
rect 124870 651400 125110 651640
rect 125220 651400 125460 651640
rect 125550 651400 125790 651640
rect 125880 651400 126120 651640
rect 126210 651400 126450 651640
rect 126560 651400 126800 651640
rect 126890 651400 127130 651640
rect 127220 651400 127460 651640
rect 127550 651400 127790 651640
rect 127900 651400 128140 651640
rect 128230 651400 128470 651640
rect 128560 651400 128800 651640
rect 128890 651400 129130 651640
rect 129240 651400 129480 651640
rect 129570 651400 129810 651640
rect 129900 651400 130140 651640
rect 130230 651400 130470 651640
rect 130580 651400 130820 651640
rect 130910 651400 131150 651640
rect 131240 651400 131480 651640
rect 131570 651400 131810 651640
rect 131920 651400 132160 651640
rect 132250 651400 132490 651640
rect 132580 651400 132820 651640
rect 132910 651400 133150 651640
rect 122190 651070 122430 651310
rect 122540 651070 122780 651310
rect 122870 651070 123110 651310
rect 123200 651070 123440 651310
rect 123530 651070 123770 651310
rect 123880 651070 124120 651310
rect 124210 651070 124450 651310
rect 124540 651070 124780 651310
rect 124870 651070 125110 651310
rect 125220 651070 125460 651310
rect 125550 651070 125790 651310
rect 125880 651070 126120 651310
rect 126210 651070 126450 651310
rect 126560 651070 126800 651310
rect 126890 651070 127130 651310
rect 127220 651070 127460 651310
rect 127550 651070 127790 651310
rect 127900 651070 128140 651310
rect 128230 651070 128470 651310
rect 128560 651070 128800 651310
rect 128890 651070 129130 651310
rect 129240 651070 129480 651310
rect 129570 651070 129810 651310
rect 129900 651070 130140 651310
rect 130230 651070 130470 651310
rect 130580 651070 130820 651310
rect 130910 651070 131150 651310
rect 131240 651070 131480 651310
rect 131570 651070 131810 651310
rect 131920 651070 132160 651310
rect 132250 651070 132490 651310
rect 132580 651070 132820 651310
rect 132910 651070 133150 651310
rect 122190 650720 122430 650960
rect 122540 650720 122780 650960
rect 122870 650720 123110 650960
rect 123200 650720 123440 650960
rect 123530 650720 123770 650960
rect 123880 650720 124120 650960
rect 124210 650720 124450 650960
rect 124540 650720 124780 650960
rect 124870 650720 125110 650960
rect 125220 650720 125460 650960
rect 125550 650720 125790 650960
rect 125880 650720 126120 650960
rect 126210 650720 126450 650960
rect 126560 650720 126800 650960
rect 126890 650720 127130 650960
rect 127220 650720 127460 650960
rect 127550 650720 127790 650960
rect 127900 650720 128140 650960
rect 128230 650720 128470 650960
rect 128560 650720 128800 650960
rect 128890 650720 129130 650960
rect 129240 650720 129480 650960
rect 129570 650720 129810 650960
rect 129900 650720 130140 650960
rect 130230 650720 130470 650960
rect 130580 650720 130820 650960
rect 130910 650720 131150 650960
rect 131240 650720 131480 650960
rect 131570 650720 131810 650960
rect 131920 650720 132160 650960
rect 132250 650720 132490 650960
rect 132580 650720 132820 650960
rect 132910 650720 133150 650960
rect 122190 650390 122430 650630
rect 122540 650390 122780 650630
rect 122870 650390 123110 650630
rect 123200 650390 123440 650630
rect 123530 650390 123770 650630
rect 123880 650390 124120 650630
rect 124210 650390 124450 650630
rect 124540 650390 124780 650630
rect 124870 650390 125110 650630
rect 125220 650390 125460 650630
rect 125550 650390 125790 650630
rect 125880 650390 126120 650630
rect 126210 650390 126450 650630
rect 126560 650390 126800 650630
rect 126890 650390 127130 650630
rect 127220 650390 127460 650630
rect 127550 650390 127790 650630
rect 127900 650390 128140 650630
rect 128230 650390 128470 650630
rect 128560 650390 128800 650630
rect 128890 650390 129130 650630
rect 129240 650390 129480 650630
rect 129570 650390 129810 650630
rect 129900 650390 130140 650630
rect 130230 650390 130470 650630
rect 130580 650390 130820 650630
rect 130910 650390 131150 650630
rect 131240 650390 131480 650630
rect 131570 650390 131810 650630
rect 131920 650390 132160 650630
rect 132250 650390 132490 650630
rect 132580 650390 132820 650630
rect 132910 650390 133150 650630
rect 122190 650060 122430 650300
rect 122540 650060 122780 650300
rect 122870 650060 123110 650300
rect 123200 650060 123440 650300
rect 123530 650060 123770 650300
rect 123880 650060 124120 650300
rect 124210 650060 124450 650300
rect 124540 650060 124780 650300
rect 124870 650060 125110 650300
rect 125220 650060 125460 650300
rect 125550 650060 125790 650300
rect 125880 650060 126120 650300
rect 126210 650060 126450 650300
rect 126560 650060 126800 650300
rect 126890 650060 127130 650300
rect 127220 650060 127460 650300
rect 127550 650060 127790 650300
rect 127900 650060 128140 650300
rect 128230 650060 128470 650300
rect 128560 650060 128800 650300
rect 128890 650060 129130 650300
rect 129240 650060 129480 650300
rect 129570 650060 129810 650300
rect 129900 650060 130140 650300
rect 130230 650060 130470 650300
rect 130580 650060 130820 650300
rect 130910 650060 131150 650300
rect 131240 650060 131480 650300
rect 131570 650060 131810 650300
rect 131920 650060 132160 650300
rect 132250 650060 132490 650300
rect 132580 650060 132820 650300
rect 132910 650060 133150 650300
rect 122190 649730 122430 649970
rect 122540 649730 122780 649970
rect 122870 649730 123110 649970
rect 123200 649730 123440 649970
rect 123530 649730 123770 649970
rect 123880 649730 124120 649970
rect 124210 649730 124450 649970
rect 124540 649730 124780 649970
rect 124870 649730 125110 649970
rect 125220 649730 125460 649970
rect 125550 649730 125790 649970
rect 125880 649730 126120 649970
rect 126210 649730 126450 649970
rect 126560 649730 126800 649970
rect 126890 649730 127130 649970
rect 127220 649730 127460 649970
rect 127550 649730 127790 649970
rect 127900 649730 128140 649970
rect 128230 649730 128470 649970
rect 128560 649730 128800 649970
rect 128890 649730 129130 649970
rect 129240 649730 129480 649970
rect 129570 649730 129810 649970
rect 129900 649730 130140 649970
rect 130230 649730 130470 649970
rect 130580 649730 130820 649970
rect 130910 649730 131150 649970
rect 131240 649730 131480 649970
rect 131570 649730 131810 649970
rect 131920 649730 132160 649970
rect 132250 649730 132490 649970
rect 132580 649730 132820 649970
rect 132910 649730 133150 649970
rect 122190 649380 122430 649620
rect 122540 649380 122780 649620
rect 122870 649380 123110 649620
rect 123200 649380 123440 649620
rect 123530 649380 123770 649620
rect 123880 649380 124120 649620
rect 124210 649380 124450 649620
rect 124540 649380 124780 649620
rect 124870 649380 125110 649620
rect 125220 649380 125460 649620
rect 125550 649380 125790 649620
rect 125880 649380 126120 649620
rect 126210 649380 126450 649620
rect 126560 649380 126800 649620
rect 126890 649380 127130 649620
rect 127220 649380 127460 649620
rect 127550 649380 127790 649620
rect 127900 649380 128140 649620
rect 128230 649380 128470 649620
rect 128560 649380 128800 649620
rect 128890 649380 129130 649620
rect 129240 649380 129480 649620
rect 129570 649380 129810 649620
rect 129900 649380 130140 649620
rect 130230 649380 130470 649620
rect 130580 649380 130820 649620
rect 130910 649380 131150 649620
rect 131240 649380 131480 649620
rect 131570 649380 131810 649620
rect 131920 649380 132160 649620
rect 132250 649380 132490 649620
rect 132580 649380 132820 649620
rect 132910 649380 133150 649620
rect 133570 660100 133810 660340
rect 133920 660100 134160 660340
rect 134250 660100 134490 660340
rect 134580 660100 134820 660340
rect 134910 660100 135150 660340
rect 135260 660100 135500 660340
rect 135590 660100 135830 660340
rect 135920 660100 136160 660340
rect 136250 660100 136490 660340
rect 136600 660100 136840 660340
rect 136930 660100 137170 660340
rect 137260 660100 137500 660340
rect 137590 660100 137830 660340
rect 137940 660100 138180 660340
rect 138270 660100 138510 660340
rect 138600 660100 138840 660340
rect 138930 660100 139170 660340
rect 139280 660100 139520 660340
rect 139610 660100 139850 660340
rect 139940 660100 140180 660340
rect 140270 660100 140510 660340
rect 140620 660100 140860 660340
rect 140950 660100 141190 660340
rect 141280 660100 141520 660340
rect 141610 660100 141850 660340
rect 141960 660100 142200 660340
rect 142290 660100 142530 660340
rect 142620 660100 142860 660340
rect 142950 660100 143190 660340
rect 143300 660100 143540 660340
rect 143630 660100 143870 660340
rect 143960 660100 144200 660340
rect 144290 660100 144530 660340
rect 133570 659770 133810 660010
rect 133920 659770 134160 660010
rect 134250 659770 134490 660010
rect 134580 659770 134820 660010
rect 134910 659770 135150 660010
rect 135260 659770 135500 660010
rect 135590 659770 135830 660010
rect 135920 659770 136160 660010
rect 136250 659770 136490 660010
rect 136600 659770 136840 660010
rect 136930 659770 137170 660010
rect 137260 659770 137500 660010
rect 137590 659770 137830 660010
rect 137940 659770 138180 660010
rect 138270 659770 138510 660010
rect 138600 659770 138840 660010
rect 138930 659770 139170 660010
rect 139280 659770 139520 660010
rect 139610 659770 139850 660010
rect 139940 659770 140180 660010
rect 140270 659770 140510 660010
rect 140620 659770 140860 660010
rect 140950 659770 141190 660010
rect 141280 659770 141520 660010
rect 141610 659770 141850 660010
rect 141960 659770 142200 660010
rect 142290 659770 142530 660010
rect 142620 659770 142860 660010
rect 142950 659770 143190 660010
rect 143300 659770 143540 660010
rect 143630 659770 143870 660010
rect 143960 659770 144200 660010
rect 144290 659770 144530 660010
rect 133570 659440 133810 659680
rect 133920 659440 134160 659680
rect 134250 659440 134490 659680
rect 134580 659440 134820 659680
rect 134910 659440 135150 659680
rect 135260 659440 135500 659680
rect 135590 659440 135830 659680
rect 135920 659440 136160 659680
rect 136250 659440 136490 659680
rect 136600 659440 136840 659680
rect 136930 659440 137170 659680
rect 137260 659440 137500 659680
rect 137590 659440 137830 659680
rect 137940 659440 138180 659680
rect 138270 659440 138510 659680
rect 138600 659440 138840 659680
rect 138930 659440 139170 659680
rect 139280 659440 139520 659680
rect 139610 659440 139850 659680
rect 139940 659440 140180 659680
rect 140270 659440 140510 659680
rect 140620 659440 140860 659680
rect 140950 659440 141190 659680
rect 141280 659440 141520 659680
rect 141610 659440 141850 659680
rect 141960 659440 142200 659680
rect 142290 659440 142530 659680
rect 142620 659440 142860 659680
rect 142950 659440 143190 659680
rect 143300 659440 143540 659680
rect 143630 659440 143870 659680
rect 143960 659440 144200 659680
rect 144290 659440 144530 659680
rect 133570 659110 133810 659350
rect 133920 659110 134160 659350
rect 134250 659110 134490 659350
rect 134580 659110 134820 659350
rect 134910 659110 135150 659350
rect 135260 659110 135500 659350
rect 135590 659110 135830 659350
rect 135920 659110 136160 659350
rect 136250 659110 136490 659350
rect 136600 659110 136840 659350
rect 136930 659110 137170 659350
rect 137260 659110 137500 659350
rect 137590 659110 137830 659350
rect 137940 659110 138180 659350
rect 138270 659110 138510 659350
rect 138600 659110 138840 659350
rect 138930 659110 139170 659350
rect 139280 659110 139520 659350
rect 139610 659110 139850 659350
rect 139940 659110 140180 659350
rect 140270 659110 140510 659350
rect 140620 659110 140860 659350
rect 140950 659110 141190 659350
rect 141280 659110 141520 659350
rect 141610 659110 141850 659350
rect 141960 659110 142200 659350
rect 142290 659110 142530 659350
rect 142620 659110 142860 659350
rect 142950 659110 143190 659350
rect 143300 659110 143540 659350
rect 143630 659110 143870 659350
rect 143960 659110 144200 659350
rect 144290 659110 144530 659350
rect 133570 658760 133810 659000
rect 133920 658760 134160 659000
rect 134250 658760 134490 659000
rect 134580 658760 134820 659000
rect 134910 658760 135150 659000
rect 135260 658760 135500 659000
rect 135590 658760 135830 659000
rect 135920 658760 136160 659000
rect 136250 658760 136490 659000
rect 136600 658760 136840 659000
rect 136930 658760 137170 659000
rect 137260 658760 137500 659000
rect 137590 658760 137830 659000
rect 137940 658760 138180 659000
rect 138270 658760 138510 659000
rect 138600 658760 138840 659000
rect 138930 658760 139170 659000
rect 139280 658760 139520 659000
rect 139610 658760 139850 659000
rect 139940 658760 140180 659000
rect 140270 658760 140510 659000
rect 140620 658760 140860 659000
rect 140950 658760 141190 659000
rect 141280 658760 141520 659000
rect 141610 658760 141850 659000
rect 141960 658760 142200 659000
rect 142290 658760 142530 659000
rect 142620 658760 142860 659000
rect 142950 658760 143190 659000
rect 143300 658760 143540 659000
rect 143630 658760 143870 659000
rect 143960 658760 144200 659000
rect 144290 658760 144530 659000
rect 133570 658430 133810 658670
rect 133920 658430 134160 658670
rect 134250 658430 134490 658670
rect 134580 658430 134820 658670
rect 134910 658430 135150 658670
rect 135260 658430 135500 658670
rect 135590 658430 135830 658670
rect 135920 658430 136160 658670
rect 136250 658430 136490 658670
rect 136600 658430 136840 658670
rect 136930 658430 137170 658670
rect 137260 658430 137500 658670
rect 137590 658430 137830 658670
rect 137940 658430 138180 658670
rect 138270 658430 138510 658670
rect 138600 658430 138840 658670
rect 138930 658430 139170 658670
rect 139280 658430 139520 658670
rect 139610 658430 139850 658670
rect 139940 658430 140180 658670
rect 140270 658430 140510 658670
rect 140620 658430 140860 658670
rect 140950 658430 141190 658670
rect 141280 658430 141520 658670
rect 141610 658430 141850 658670
rect 141960 658430 142200 658670
rect 142290 658430 142530 658670
rect 142620 658430 142860 658670
rect 142950 658430 143190 658670
rect 143300 658430 143540 658670
rect 143630 658430 143870 658670
rect 143960 658430 144200 658670
rect 144290 658430 144530 658670
rect 133570 658100 133810 658340
rect 133920 658100 134160 658340
rect 134250 658100 134490 658340
rect 134580 658100 134820 658340
rect 134910 658100 135150 658340
rect 135260 658100 135500 658340
rect 135590 658100 135830 658340
rect 135920 658100 136160 658340
rect 136250 658100 136490 658340
rect 136600 658100 136840 658340
rect 136930 658100 137170 658340
rect 137260 658100 137500 658340
rect 137590 658100 137830 658340
rect 137940 658100 138180 658340
rect 138270 658100 138510 658340
rect 138600 658100 138840 658340
rect 138930 658100 139170 658340
rect 139280 658100 139520 658340
rect 139610 658100 139850 658340
rect 139940 658100 140180 658340
rect 140270 658100 140510 658340
rect 140620 658100 140860 658340
rect 140950 658100 141190 658340
rect 141280 658100 141520 658340
rect 141610 658100 141850 658340
rect 141960 658100 142200 658340
rect 142290 658100 142530 658340
rect 142620 658100 142860 658340
rect 142950 658100 143190 658340
rect 143300 658100 143540 658340
rect 143630 658100 143870 658340
rect 143960 658100 144200 658340
rect 144290 658100 144530 658340
rect 133570 657770 133810 658010
rect 133920 657770 134160 658010
rect 134250 657770 134490 658010
rect 134580 657770 134820 658010
rect 134910 657770 135150 658010
rect 135260 657770 135500 658010
rect 135590 657770 135830 658010
rect 135920 657770 136160 658010
rect 136250 657770 136490 658010
rect 136600 657770 136840 658010
rect 136930 657770 137170 658010
rect 137260 657770 137500 658010
rect 137590 657770 137830 658010
rect 137940 657770 138180 658010
rect 138270 657770 138510 658010
rect 138600 657770 138840 658010
rect 138930 657770 139170 658010
rect 139280 657770 139520 658010
rect 139610 657770 139850 658010
rect 139940 657770 140180 658010
rect 140270 657770 140510 658010
rect 140620 657770 140860 658010
rect 140950 657770 141190 658010
rect 141280 657770 141520 658010
rect 141610 657770 141850 658010
rect 141960 657770 142200 658010
rect 142290 657770 142530 658010
rect 142620 657770 142860 658010
rect 142950 657770 143190 658010
rect 143300 657770 143540 658010
rect 143630 657770 143870 658010
rect 143960 657770 144200 658010
rect 144290 657770 144530 658010
rect 133570 657420 133810 657660
rect 133920 657420 134160 657660
rect 134250 657420 134490 657660
rect 134580 657420 134820 657660
rect 134910 657420 135150 657660
rect 135260 657420 135500 657660
rect 135590 657420 135830 657660
rect 135920 657420 136160 657660
rect 136250 657420 136490 657660
rect 136600 657420 136840 657660
rect 136930 657420 137170 657660
rect 137260 657420 137500 657660
rect 137590 657420 137830 657660
rect 137940 657420 138180 657660
rect 138270 657420 138510 657660
rect 138600 657420 138840 657660
rect 138930 657420 139170 657660
rect 139280 657420 139520 657660
rect 139610 657420 139850 657660
rect 139940 657420 140180 657660
rect 140270 657420 140510 657660
rect 140620 657420 140860 657660
rect 140950 657420 141190 657660
rect 141280 657420 141520 657660
rect 141610 657420 141850 657660
rect 141960 657420 142200 657660
rect 142290 657420 142530 657660
rect 142620 657420 142860 657660
rect 142950 657420 143190 657660
rect 143300 657420 143540 657660
rect 143630 657420 143870 657660
rect 143960 657420 144200 657660
rect 144290 657420 144530 657660
rect 133570 657090 133810 657330
rect 133920 657090 134160 657330
rect 134250 657090 134490 657330
rect 134580 657090 134820 657330
rect 134910 657090 135150 657330
rect 135260 657090 135500 657330
rect 135590 657090 135830 657330
rect 135920 657090 136160 657330
rect 136250 657090 136490 657330
rect 136600 657090 136840 657330
rect 136930 657090 137170 657330
rect 137260 657090 137500 657330
rect 137590 657090 137830 657330
rect 137940 657090 138180 657330
rect 138270 657090 138510 657330
rect 138600 657090 138840 657330
rect 138930 657090 139170 657330
rect 139280 657090 139520 657330
rect 139610 657090 139850 657330
rect 139940 657090 140180 657330
rect 140270 657090 140510 657330
rect 140620 657090 140860 657330
rect 140950 657090 141190 657330
rect 141280 657090 141520 657330
rect 141610 657090 141850 657330
rect 141960 657090 142200 657330
rect 142290 657090 142530 657330
rect 142620 657090 142860 657330
rect 142950 657090 143190 657330
rect 143300 657090 143540 657330
rect 143630 657090 143870 657330
rect 143960 657090 144200 657330
rect 144290 657090 144530 657330
rect 133570 656760 133810 657000
rect 133920 656760 134160 657000
rect 134250 656760 134490 657000
rect 134580 656760 134820 657000
rect 134910 656760 135150 657000
rect 135260 656760 135500 657000
rect 135590 656760 135830 657000
rect 135920 656760 136160 657000
rect 136250 656760 136490 657000
rect 136600 656760 136840 657000
rect 136930 656760 137170 657000
rect 137260 656760 137500 657000
rect 137590 656760 137830 657000
rect 137940 656760 138180 657000
rect 138270 656760 138510 657000
rect 138600 656760 138840 657000
rect 138930 656760 139170 657000
rect 139280 656760 139520 657000
rect 139610 656760 139850 657000
rect 139940 656760 140180 657000
rect 140270 656760 140510 657000
rect 140620 656760 140860 657000
rect 140950 656760 141190 657000
rect 141280 656760 141520 657000
rect 141610 656760 141850 657000
rect 141960 656760 142200 657000
rect 142290 656760 142530 657000
rect 142620 656760 142860 657000
rect 142950 656760 143190 657000
rect 143300 656760 143540 657000
rect 143630 656760 143870 657000
rect 143960 656760 144200 657000
rect 144290 656760 144530 657000
rect 133570 656430 133810 656670
rect 133920 656430 134160 656670
rect 134250 656430 134490 656670
rect 134580 656430 134820 656670
rect 134910 656430 135150 656670
rect 135260 656430 135500 656670
rect 135590 656430 135830 656670
rect 135920 656430 136160 656670
rect 136250 656430 136490 656670
rect 136600 656430 136840 656670
rect 136930 656430 137170 656670
rect 137260 656430 137500 656670
rect 137590 656430 137830 656670
rect 137940 656430 138180 656670
rect 138270 656430 138510 656670
rect 138600 656430 138840 656670
rect 138930 656430 139170 656670
rect 139280 656430 139520 656670
rect 139610 656430 139850 656670
rect 139940 656430 140180 656670
rect 140270 656430 140510 656670
rect 140620 656430 140860 656670
rect 140950 656430 141190 656670
rect 141280 656430 141520 656670
rect 141610 656430 141850 656670
rect 141960 656430 142200 656670
rect 142290 656430 142530 656670
rect 142620 656430 142860 656670
rect 142950 656430 143190 656670
rect 143300 656430 143540 656670
rect 143630 656430 143870 656670
rect 143960 656430 144200 656670
rect 144290 656430 144530 656670
rect 133570 656080 133810 656320
rect 133920 656080 134160 656320
rect 134250 656080 134490 656320
rect 134580 656080 134820 656320
rect 134910 656080 135150 656320
rect 135260 656080 135500 656320
rect 135590 656080 135830 656320
rect 135920 656080 136160 656320
rect 136250 656080 136490 656320
rect 136600 656080 136840 656320
rect 136930 656080 137170 656320
rect 137260 656080 137500 656320
rect 137590 656080 137830 656320
rect 137940 656080 138180 656320
rect 138270 656080 138510 656320
rect 138600 656080 138840 656320
rect 138930 656080 139170 656320
rect 139280 656080 139520 656320
rect 139610 656080 139850 656320
rect 139940 656080 140180 656320
rect 140270 656080 140510 656320
rect 140620 656080 140860 656320
rect 140950 656080 141190 656320
rect 141280 656080 141520 656320
rect 141610 656080 141850 656320
rect 141960 656080 142200 656320
rect 142290 656080 142530 656320
rect 142620 656080 142860 656320
rect 142950 656080 143190 656320
rect 143300 656080 143540 656320
rect 143630 656080 143870 656320
rect 143960 656080 144200 656320
rect 144290 656080 144530 656320
rect 133570 655750 133810 655990
rect 133920 655750 134160 655990
rect 134250 655750 134490 655990
rect 134580 655750 134820 655990
rect 134910 655750 135150 655990
rect 135260 655750 135500 655990
rect 135590 655750 135830 655990
rect 135920 655750 136160 655990
rect 136250 655750 136490 655990
rect 136600 655750 136840 655990
rect 136930 655750 137170 655990
rect 137260 655750 137500 655990
rect 137590 655750 137830 655990
rect 137940 655750 138180 655990
rect 138270 655750 138510 655990
rect 138600 655750 138840 655990
rect 138930 655750 139170 655990
rect 139280 655750 139520 655990
rect 139610 655750 139850 655990
rect 139940 655750 140180 655990
rect 140270 655750 140510 655990
rect 140620 655750 140860 655990
rect 140950 655750 141190 655990
rect 141280 655750 141520 655990
rect 141610 655750 141850 655990
rect 141960 655750 142200 655990
rect 142290 655750 142530 655990
rect 142620 655750 142860 655990
rect 142950 655750 143190 655990
rect 143300 655750 143540 655990
rect 143630 655750 143870 655990
rect 143960 655750 144200 655990
rect 144290 655750 144530 655990
rect 133570 655420 133810 655660
rect 133920 655420 134160 655660
rect 134250 655420 134490 655660
rect 134580 655420 134820 655660
rect 134910 655420 135150 655660
rect 135260 655420 135500 655660
rect 135590 655420 135830 655660
rect 135920 655420 136160 655660
rect 136250 655420 136490 655660
rect 136600 655420 136840 655660
rect 136930 655420 137170 655660
rect 137260 655420 137500 655660
rect 137590 655420 137830 655660
rect 137940 655420 138180 655660
rect 138270 655420 138510 655660
rect 138600 655420 138840 655660
rect 138930 655420 139170 655660
rect 139280 655420 139520 655660
rect 139610 655420 139850 655660
rect 139940 655420 140180 655660
rect 140270 655420 140510 655660
rect 140620 655420 140860 655660
rect 140950 655420 141190 655660
rect 141280 655420 141520 655660
rect 141610 655420 141850 655660
rect 141960 655420 142200 655660
rect 142290 655420 142530 655660
rect 142620 655420 142860 655660
rect 142950 655420 143190 655660
rect 143300 655420 143540 655660
rect 143630 655420 143870 655660
rect 143960 655420 144200 655660
rect 144290 655420 144530 655660
rect 133570 655090 133810 655330
rect 133920 655090 134160 655330
rect 134250 655090 134490 655330
rect 134580 655090 134820 655330
rect 134910 655090 135150 655330
rect 135260 655090 135500 655330
rect 135590 655090 135830 655330
rect 135920 655090 136160 655330
rect 136250 655090 136490 655330
rect 136600 655090 136840 655330
rect 136930 655090 137170 655330
rect 137260 655090 137500 655330
rect 137590 655090 137830 655330
rect 137940 655090 138180 655330
rect 138270 655090 138510 655330
rect 138600 655090 138840 655330
rect 138930 655090 139170 655330
rect 139280 655090 139520 655330
rect 139610 655090 139850 655330
rect 139940 655090 140180 655330
rect 140270 655090 140510 655330
rect 140620 655090 140860 655330
rect 140950 655090 141190 655330
rect 141280 655090 141520 655330
rect 141610 655090 141850 655330
rect 141960 655090 142200 655330
rect 142290 655090 142530 655330
rect 142620 655090 142860 655330
rect 142950 655090 143190 655330
rect 143300 655090 143540 655330
rect 143630 655090 143870 655330
rect 143960 655090 144200 655330
rect 144290 655090 144530 655330
rect 133570 654740 133810 654980
rect 133920 654740 134160 654980
rect 134250 654740 134490 654980
rect 134580 654740 134820 654980
rect 134910 654740 135150 654980
rect 135260 654740 135500 654980
rect 135590 654740 135830 654980
rect 135920 654740 136160 654980
rect 136250 654740 136490 654980
rect 136600 654740 136840 654980
rect 136930 654740 137170 654980
rect 137260 654740 137500 654980
rect 137590 654740 137830 654980
rect 137940 654740 138180 654980
rect 138270 654740 138510 654980
rect 138600 654740 138840 654980
rect 138930 654740 139170 654980
rect 139280 654740 139520 654980
rect 139610 654740 139850 654980
rect 139940 654740 140180 654980
rect 140270 654740 140510 654980
rect 140620 654740 140860 654980
rect 140950 654740 141190 654980
rect 141280 654740 141520 654980
rect 141610 654740 141850 654980
rect 141960 654740 142200 654980
rect 142290 654740 142530 654980
rect 142620 654740 142860 654980
rect 142950 654740 143190 654980
rect 143300 654740 143540 654980
rect 143630 654740 143870 654980
rect 143960 654740 144200 654980
rect 144290 654740 144530 654980
rect 133570 654410 133810 654650
rect 133920 654410 134160 654650
rect 134250 654410 134490 654650
rect 134580 654410 134820 654650
rect 134910 654410 135150 654650
rect 135260 654410 135500 654650
rect 135590 654410 135830 654650
rect 135920 654410 136160 654650
rect 136250 654410 136490 654650
rect 136600 654410 136840 654650
rect 136930 654410 137170 654650
rect 137260 654410 137500 654650
rect 137590 654410 137830 654650
rect 137940 654410 138180 654650
rect 138270 654410 138510 654650
rect 138600 654410 138840 654650
rect 138930 654410 139170 654650
rect 139280 654410 139520 654650
rect 139610 654410 139850 654650
rect 139940 654410 140180 654650
rect 140270 654410 140510 654650
rect 140620 654410 140860 654650
rect 140950 654410 141190 654650
rect 141280 654410 141520 654650
rect 141610 654410 141850 654650
rect 141960 654410 142200 654650
rect 142290 654410 142530 654650
rect 142620 654410 142860 654650
rect 142950 654410 143190 654650
rect 143300 654410 143540 654650
rect 143630 654410 143870 654650
rect 143960 654410 144200 654650
rect 144290 654410 144530 654650
rect 133570 654080 133810 654320
rect 133920 654080 134160 654320
rect 134250 654080 134490 654320
rect 134580 654080 134820 654320
rect 134910 654080 135150 654320
rect 135260 654080 135500 654320
rect 135590 654080 135830 654320
rect 135920 654080 136160 654320
rect 136250 654080 136490 654320
rect 136600 654080 136840 654320
rect 136930 654080 137170 654320
rect 137260 654080 137500 654320
rect 137590 654080 137830 654320
rect 137940 654080 138180 654320
rect 138270 654080 138510 654320
rect 138600 654080 138840 654320
rect 138930 654080 139170 654320
rect 139280 654080 139520 654320
rect 139610 654080 139850 654320
rect 139940 654080 140180 654320
rect 140270 654080 140510 654320
rect 140620 654080 140860 654320
rect 140950 654080 141190 654320
rect 141280 654080 141520 654320
rect 141610 654080 141850 654320
rect 141960 654080 142200 654320
rect 142290 654080 142530 654320
rect 142620 654080 142860 654320
rect 142950 654080 143190 654320
rect 143300 654080 143540 654320
rect 143630 654080 143870 654320
rect 143960 654080 144200 654320
rect 144290 654080 144530 654320
rect 133570 653750 133810 653990
rect 133920 653750 134160 653990
rect 134250 653750 134490 653990
rect 134580 653750 134820 653990
rect 134910 653750 135150 653990
rect 135260 653750 135500 653990
rect 135590 653750 135830 653990
rect 135920 653750 136160 653990
rect 136250 653750 136490 653990
rect 136600 653750 136840 653990
rect 136930 653750 137170 653990
rect 137260 653750 137500 653990
rect 137590 653750 137830 653990
rect 137940 653750 138180 653990
rect 138270 653750 138510 653990
rect 138600 653750 138840 653990
rect 138930 653750 139170 653990
rect 139280 653750 139520 653990
rect 139610 653750 139850 653990
rect 139940 653750 140180 653990
rect 140270 653750 140510 653990
rect 140620 653750 140860 653990
rect 140950 653750 141190 653990
rect 141280 653750 141520 653990
rect 141610 653750 141850 653990
rect 141960 653750 142200 653990
rect 142290 653750 142530 653990
rect 142620 653750 142860 653990
rect 142950 653750 143190 653990
rect 143300 653750 143540 653990
rect 143630 653750 143870 653990
rect 143960 653750 144200 653990
rect 144290 653750 144530 653990
rect 133570 653400 133810 653640
rect 133920 653400 134160 653640
rect 134250 653400 134490 653640
rect 134580 653400 134820 653640
rect 134910 653400 135150 653640
rect 135260 653400 135500 653640
rect 135590 653400 135830 653640
rect 135920 653400 136160 653640
rect 136250 653400 136490 653640
rect 136600 653400 136840 653640
rect 136930 653400 137170 653640
rect 137260 653400 137500 653640
rect 137590 653400 137830 653640
rect 137940 653400 138180 653640
rect 138270 653400 138510 653640
rect 138600 653400 138840 653640
rect 138930 653400 139170 653640
rect 139280 653400 139520 653640
rect 139610 653400 139850 653640
rect 139940 653400 140180 653640
rect 140270 653400 140510 653640
rect 140620 653400 140860 653640
rect 140950 653400 141190 653640
rect 141280 653400 141520 653640
rect 141610 653400 141850 653640
rect 141960 653400 142200 653640
rect 142290 653400 142530 653640
rect 142620 653400 142860 653640
rect 142950 653400 143190 653640
rect 143300 653400 143540 653640
rect 143630 653400 143870 653640
rect 143960 653400 144200 653640
rect 144290 653400 144530 653640
rect 133570 653070 133810 653310
rect 133920 653070 134160 653310
rect 134250 653070 134490 653310
rect 134580 653070 134820 653310
rect 134910 653070 135150 653310
rect 135260 653070 135500 653310
rect 135590 653070 135830 653310
rect 135920 653070 136160 653310
rect 136250 653070 136490 653310
rect 136600 653070 136840 653310
rect 136930 653070 137170 653310
rect 137260 653070 137500 653310
rect 137590 653070 137830 653310
rect 137940 653070 138180 653310
rect 138270 653070 138510 653310
rect 138600 653070 138840 653310
rect 138930 653070 139170 653310
rect 139280 653070 139520 653310
rect 139610 653070 139850 653310
rect 139940 653070 140180 653310
rect 140270 653070 140510 653310
rect 140620 653070 140860 653310
rect 140950 653070 141190 653310
rect 141280 653070 141520 653310
rect 141610 653070 141850 653310
rect 141960 653070 142200 653310
rect 142290 653070 142530 653310
rect 142620 653070 142860 653310
rect 142950 653070 143190 653310
rect 143300 653070 143540 653310
rect 143630 653070 143870 653310
rect 143960 653070 144200 653310
rect 144290 653070 144530 653310
rect 133570 652740 133810 652980
rect 133920 652740 134160 652980
rect 134250 652740 134490 652980
rect 134580 652740 134820 652980
rect 134910 652740 135150 652980
rect 135260 652740 135500 652980
rect 135590 652740 135830 652980
rect 135920 652740 136160 652980
rect 136250 652740 136490 652980
rect 136600 652740 136840 652980
rect 136930 652740 137170 652980
rect 137260 652740 137500 652980
rect 137590 652740 137830 652980
rect 137940 652740 138180 652980
rect 138270 652740 138510 652980
rect 138600 652740 138840 652980
rect 138930 652740 139170 652980
rect 139280 652740 139520 652980
rect 139610 652740 139850 652980
rect 139940 652740 140180 652980
rect 140270 652740 140510 652980
rect 140620 652740 140860 652980
rect 140950 652740 141190 652980
rect 141280 652740 141520 652980
rect 141610 652740 141850 652980
rect 141960 652740 142200 652980
rect 142290 652740 142530 652980
rect 142620 652740 142860 652980
rect 142950 652740 143190 652980
rect 143300 652740 143540 652980
rect 143630 652740 143870 652980
rect 143960 652740 144200 652980
rect 144290 652740 144530 652980
rect 133570 652410 133810 652650
rect 133920 652410 134160 652650
rect 134250 652410 134490 652650
rect 134580 652410 134820 652650
rect 134910 652410 135150 652650
rect 135260 652410 135500 652650
rect 135590 652410 135830 652650
rect 135920 652410 136160 652650
rect 136250 652410 136490 652650
rect 136600 652410 136840 652650
rect 136930 652410 137170 652650
rect 137260 652410 137500 652650
rect 137590 652410 137830 652650
rect 137940 652410 138180 652650
rect 138270 652410 138510 652650
rect 138600 652410 138840 652650
rect 138930 652410 139170 652650
rect 139280 652410 139520 652650
rect 139610 652410 139850 652650
rect 139940 652410 140180 652650
rect 140270 652410 140510 652650
rect 140620 652410 140860 652650
rect 140950 652410 141190 652650
rect 141280 652410 141520 652650
rect 141610 652410 141850 652650
rect 141960 652410 142200 652650
rect 142290 652410 142530 652650
rect 142620 652410 142860 652650
rect 142950 652410 143190 652650
rect 143300 652410 143540 652650
rect 143630 652410 143870 652650
rect 143960 652410 144200 652650
rect 144290 652410 144530 652650
rect 133570 652060 133810 652300
rect 133920 652060 134160 652300
rect 134250 652060 134490 652300
rect 134580 652060 134820 652300
rect 134910 652060 135150 652300
rect 135260 652060 135500 652300
rect 135590 652060 135830 652300
rect 135920 652060 136160 652300
rect 136250 652060 136490 652300
rect 136600 652060 136840 652300
rect 136930 652060 137170 652300
rect 137260 652060 137500 652300
rect 137590 652060 137830 652300
rect 137940 652060 138180 652300
rect 138270 652060 138510 652300
rect 138600 652060 138840 652300
rect 138930 652060 139170 652300
rect 139280 652060 139520 652300
rect 139610 652060 139850 652300
rect 139940 652060 140180 652300
rect 140270 652060 140510 652300
rect 140620 652060 140860 652300
rect 140950 652060 141190 652300
rect 141280 652060 141520 652300
rect 141610 652060 141850 652300
rect 141960 652060 142200 652300
rect 142290 652060 142530 652300
rect 142620 652060 142860 652300
rect 142950 652060 143190 652300
rect 143300 652060 143540 652300
rect 143630 652060 143870 652300
rect 143960 652060 144200 652300
rect 144290 652060 144530 652300
rect 133570 651730 133810 651970
rect 133920 651730 134160 651970
rect 134250 651730 134490 651970
rect 134580 651730 134820 651970
rect 134910 651730 135150 651970
rect 135260 651730 135500 651970
rect 135590 651730 135830 651970
rect 135920 651730 136160 651970
rect 136250 651730 136490 651970
rect 136600 651730 136840 651970
rect 136930 651730 137170 651970
rect 137260 651730 137500 651970
rect 137590 651730 137830 651970
rect 137940 651730 138180 651970
rect 138270 651730 138510 651970
rect 138600 651730 138840 651970
rect 138930 651730 139170 651970
rect 139280 651730 139520 651970
rect 139610 651730 139850 651970
rect 139940 651730 140180 651970
rect 140270 651730 140510 651970
rect 140620 651730 140860 651970
rect 140950 651730 141190 651970
rect 141280 651730 141520 651970
rect 141610 651730 141850 651970
rect 141960 651730 142200 651970
rect 142290 651730 142530 651970
rect 142620 651730 142860 651970
rect 142950 651730 143190 651970
rect 143300 651730 143540 651970
rect 143630 651730 143870 651970
rect 143960 651730 144200 651970
rect 144290 651730 144530 651970
rect 133570 651400 133810 651640
rect 133920 651400 134160 651640
rect 134250 651400 134490 651640
rect 134580 651400 134820 651640
rect 134910 651400 135150 651640
rect 135260 651400 135500 651640
rect 135590 651400 135830 651640
rect 135920 651400 136160 651640
rect 136250 651400 136490 651640
rect 136600 651400 136840 651640
rect 136930 651400 137170 651640
rect 137260 651400 137500 651640
rect 137590 651400 137830 651640
rect 137940 651400 138180 651640
rect 138270 651400 138510 651640
rect 138600 651400 138840 651640
rect 138930 651400 139170 651640
rect 139280 651400 139520 651640
rect 139610 651400 139850 651640
rect 139940 651400 140180 651640
rect 140270 651400 140510 651640
rect 140620 651400 140860 651640
rect 140950 651400 141190 651640
rect 141280 651400 141520 651640
rect 141610 651400 141850 651640
rect 141960 651400 142200 651640
rect 142290 651400 142530 651640
rect 142620 651400 142860 651640
rect 142950 651400 143190 651640
rect 143300 651400 143540 651640
rect 143630 651400 143870 651640
rect 143960 651400 144200 651640
rect 144290 651400 144530 651640
rect 133570 651070 133810 651310
rect 133920 651070 134160 651310
rect 134250 651070 134490 651310
rect 134580 651070 134820 651310
rect 134910 651070 135150 651310
rect 135260 651070 135500 651310
rect 135590 651070 135830 651310
rect 135920 651070 136160 651310
rect 136250 651070 136490 651310
rect 136600 651070 136840 651310
rect 136930 651070 137170 651310
rect 137260 651070 137500 651310
rect 137590 651070 137830 651310
rect 137940 651070 138180 651310
rect 138270 651070 138510 651310
rect 138600 651070 138840 651310
rect 138930 651070 139170 651310
rect 139280 651070 139520 651310
rect 139610 651070 139850 651310
rect 139940 651070 140180 651310
rect 140270 651070 140510 651310
rect 140620 651070 140860 651310
rect 140950 651070 141190 651310
rect 141280 651070 141520 651310
rect 141610 651070 141850 651310
rect 141960 651070 142200 651310
rect 142290 651070 142530 651310
rect 142620 651070 142860 651310
rect 142950 651070 143190 651310
rect 143300 651070 143540 651310
rect 143630 651070 143870 651310
rect 143960 651070 144200 651310
rect 144290 651070 144530 651310
rect 133570 650720 133810 650960
rect 133920 650720 134160 650960
rect 134250 650720 134490 650960
rect 134580 650720 134820 650960
rect 134910 650720 135150 650960
rect 135260 650720 135500 650960
rect 135590 650720 135830 650960
rect 135920 650720 136160 650960
rect 136250 650720 136490 650960
rect 136600 650720 136840 650960
rect 136930 650720 137170 650960
rect 137260 650720 137500 650960
rect 137590 650720 137830 650960
rect 137940 650720 138180 650960
rect 138270 650720 138510 650960
rect 138600 650720 138840 650960
rect 138930 650720 139170 650960
rect 139280 650720 139520 650960
rect 139610 650720 139850 650960
rect 139940 650720 140180 650960
rect 140270 650720 140510 650960
rect 140620 650720 140860 650960
rect 140950 650720 141190 650960
rect 141280 650720 141520 650960
rect 141610 650720 141850 650960
rect 141960 650720 142200 650960
rect 142290 650720 142530 650960
rect 142620 650720 142860 650960
rect 142950 650720 143190 650960
rect 143300 650720 143540 650960
rect 143630 650720 143870 650960
rect 143960 650720 144200 650960
rect 144290 650720 144530 650960
rect 133570 650390 133810 650630
rect 133920 650390 134160 650630
rect 134250 650390 134490 650630
rect 134580 650390 134820 650630
rect 134910 650390 135150 650630
rect 135260 650390 135500 650630
rect 135590 650390 135830 650630
rect 135920 650390 136160 650630
rect 136250 650390 136490 650630
rect 136600 650390 136840 650630
rect 136930 650390 137170 650630
rect 137260 650390 137500 650630
rect 137590 650390 137830 650630
rect 137940 650390 138180 650630
rect 138270 650390 138510 650630
rect 138600 650390 138840 650630
rect 138930 650390 139170 650630
rect 139280 650390 139520 650630
rect 139610 650390 139850 650630
rect 139940 650390 140180 650630
rect 140270 650390 140510 650630
rect 140620 650390 140860 650630
rect 140950 650390 141190 650630
rect 141280 650390 141520 650630
rect 141610 650390 141850 650630
rect 141960 650390 142200 650630
rect 142290 650390 142530 650630
rect 142620 650390 142860 650630
rect 142950 650390 143190 650630
rect 143300 650390 143540 650630
rect 143630 650390 143870 650630
rect 143960 650390 144200 650630
rect 144290 650390 144530 650630
rect 133570 650060 133810 650300
rect 133920 650060 134160 650300
rect 134250 650060 134490 650300
rect 134580 650060 134820 650300
rect 134910 650060 135150 650300
rect 135260 650060 135500 650300
rect 135590 650060 135830 650300
rect 135920 650060 136160 650300
rect 136250 650060 136490 650300
rect 136600 650060 136840 650300
rect 136930 650060 137170 650300
rect 137260 650060 137500 650300
rect 137590 650060 137830 650300
rect 137940 650060 138180 650300
rect 138270 650060 138510 650300
rect 138600 650060 138840 650300
rect 138930 650060 139170 650300
rect 139280 650060 139520 650300
rect 139610 650060 139850 650300
rect 139940 650060 140180 650300
rect 140270 650060 140510 650300
rect 140620 650060 140860 650300
rect 140950 650060 141190 650300
rect 141280 650060 141520 650300
rect 141610 650060 141850 650300
rect 141960 650060 142200 650300
rect 142290 650060 142530 650300
rect 142620 650060 142860 650300
rect 142950 650060 143190 650300
rect 143300 650060 143540 650300
rect 143630 650060 143870 650300
rect 143960 650060 144200 650300
rect 144290 650060 144530 650300
rect 133570 649730 133810 649970
rect 133920 649730 134160 649970
rect 134250 649730 134490 649970
rect 134580 649730 134820 649970
rect 134910 649730 135150 649970
rect 135260 649730 135500 649970
rect 135590 649730 135830 649970
rect 135920 649730 136160 649970
rect 136250 649730 136490 649970
rect 136600 649730 136840 649970
rect 136930 649730 137170 649970
rect 137260 649730 137500 649970
rect 137590 649730 137830 649970
rect 137940 649730 138180 649970
rect 138270 649730 138510 649970
rect 138600 649730 138840 649970
rect 138930 649730 139170 649970
rect 139280 649730 139520 649970
rect 139610 649730 139850 649970
rect 139940 649730 140180 649970
rect 140270 649730 140510 649970
rect 140620 649730 140860 649970
rect 140950 649730 141190 649970
rect 141280 649730 141520 649970
rect 141610 649730 141850 649970
rect 141960 649730 142200 649970
rect 142290 649730 142530 649970
rect 142620 649730 142860 649970
rect 142950 649730 143190 649970
rect 143300 649730 143540 649970
rect 143630 649730 143870 649970
rect 143960 649730 144200 649970
rect 144290 649730 144530 649970
rect 133570 649380 133810 649620
rect 133920 649380 134160 649620
rect 134250 649380 134490 649620
rect 134580 649380 134820 649620
rect 134910 649380 135150 649620
rect 135260 649380 135500 649620
rect 135590 649380 135830 649620
rect 135920 649380 136160 649620
rect 136250 649380 136490 649620
rect 136600 649380 136840 649620
rect 136930 649380 137170 649620
rect 137260 649380 137500 649620
rect 137590 649380 137830 649620
rect 137940 649380 138180 649620
rect 138270 649380 138510 649620
rect 138600 649380 138840 649620
rect 138930 649380 139170 649620
rect 139280 649380 139520 649620
rect 139610 649380 139850 649620
rect 139940 649380 140180 649620
rect 140270 649380 140510 649620
rect 140620 649380 140860 649620
rect 140950 649380 141190 649620
rect 141280 649380 141520 649620
rect 141610 649380 141850 649620
rect 141960 649380 142200 649620
rect 142290 649380 142530 649620
rect 142620 649380 142860 649620
rect 142950 649380 143190 649620
rect 143300 649380 143540 649620
rect 143630 649380 143870 649620
rect 143960 649380 144200 649620
rect 144290 649380 144530 649620
rect 144950 660100 145190 660340
rect 145300 660100 145540 660340
rect 145630 660100 145870 660340
rect 145960 660100 146200 660340
rect 146290 660100 146530 660340
rect 146640 660100 146880 660340
rect 146970 660100 147210 660340
rect 147300 660100 147540 660340
rect 147630 660100 147870 660340
rect 147980 660100 148220 660340
rect 148310 660100 148550 660340
rect 148640 660100 148880 660340
rect 148970 660100 149210 660340
rect 149320 660100 149560 660340
rect 149650 660100 149890 660340
rect 149980 660100 150220 660340
rect 150310 660100 150550 660340
rect 150660 660100 150900 660340
rect 150990 660100 151230 660340
rect 151320 660100 151560 660340
rect 151650 660100 151890 660340
rect 152000 660100 152240 660340
rect 152330 660100 152570 660340
rect 152660 660100 152900 660340
rect 152990 660100 153230 660340
rect 153340 660100 153580 660340
rect 153670 660100 153910 660340
rect 154000 660100 154240 660340
rect 154330 660100 154570 660340
rect 154680 660100 154920 660340
rect 155010 660100 155250 660340
rect 155340 660100 155580 660340
rect 155670 660100 155910 660340
rect 144950 659770 145190 660010
rect 145300 659770 145540 660010
rect 145630 659770 145870 660010
rect 145960 659770 146200 660010
rect 146290 659770 146530 660010
rect 146640 659770 146880 660010
rect 146970 659770 147210 660010
rect 147300 659770 147540 660010
rect 147630 659770 147870 660010
rect 147980 659770 148220 660010
rect 148310 659770 148550 660010
rect 148640 659770 148880 660010
rect 148970 659770 149210 660010
rect 149320 659770 149560 660010
rect 149650 659770 149890 660010
rect 149980 659770 150220 660010
rect 150310 659770 150550 660010
rect 150660 659770 150900 660010
rect 150990 659770 151230 660010
rect 151320 659770 151560 660010
rect 151650 659770 151890 660010
rect 152000 659770 152240 660010
rect 152330 659770 152570 660010
rect 152660 659770 152900 660010
rect 152990 659770 153230 660010
rect 153340 659770 153580 660010
rect 153670 659770 153910 660010
rect 154000 659770 154240 660010
rect 154330 659770 154570 660010
rect 154680 659770 154920 660010
rect 155010 659770 155250 660010
rect 155340 659770 155580 660010
rect 155670 659770 155910 660010
rect 144950 659440 145190 659680
rect 145300 659440 145540 659680
rect 145630 659440 145870 659680
rect 145960 659440 146200 659680
rect 146290 659440 146530 659680
rect 146640 659440 146880 659680
rect 146970 659440 147210 659680
rect 147300 659440 147540 659680
rect 147630 659440 147870 659680
rect 147980 659440 148220 659680
rect 148310 659440 148550 659680
rect 148640 659440 148880 659680
rect 148970 659440 149210 659680
rect 149320 659440 149560 659680
rect 149650 659440 149890 659680
rect 149980 659440 150220 659680
rect 150310 659440 150550 659680
rect 150660 659440 150900 659680
rect 150990 659440 151230 659680
rect 151320 659440 151560 659680
rect 151650 659440 151890 659680
rect 152000 659440 152240 659680
rect 152330 659440 152570 659680
rect 152660 659440 152900 659680
rect 152990 659440 153230 659680
rect 153340 659440 153580 659680
rect 153670 659440 153910 659680
rect 154000 659440 154240 659680
rect 154330 659440 154570 659680
rect 154680 659440 154920 659680
rect 155010 659440 155250 659680
rect 155340 659440 155580 659680
rect 155670 659440 155910 659680
rect 144950 659110 145190 659350
rect 145300 659110 145540 659350
rect 145630 659110 145870 659350
rect 145960 659110 146200 659350
rect 146290 659110 146530 659350
rect 146640 659110 146880 659350
rect 146970 659110 147210 659350
rect 147300 659110 147540 659350
rect 147630 659110 147870 659350
rect 147980 659110 148220 659350
rect 148310 659110 148550 659350
rect 148640 659110 148880 659350
rect 148970 659110 149210 659350
rect 149320 659110 149560 659350
rect 149650 659110 149890 659350
rect 149980 659110 150220 659350
rect 150310 659110 150550 659350
rect 150660 659110 150900 659350
rect 150990 659110 151230 659350
rect 151320 659110 151560 659350
rect 151650 659110 151890 659350
rect 152000 659110 152240 659350
rect 152330 659110 152570 659350
rect 152660 659110 152900 659350
rect 152990 659110 153230 659350
rect 153340 659110 153580 659350
rect 153670 659110 153910 659350
rect 154000 659110 154240 659350
rect 154330 659110 154570 659350
rect 154680 659110 154920 659350
rect 155010 659110 155250 659350
rect 155340 659110 155580 659350
rect 155670 659110 155910 659350
rect 144950 658760 145190 659000
rect 145300 658760 145540 659000
rect 145630 658760 145870 659000
rect 145960 658760 146200 659000
rect 146290 658760 146530 659000
rect 146640 658760 146880 659000
rect 146970 658760 147210 659000
rect 147300 658760 147540 659000
rect 147630 658760 147870 659000
rect 147980 658760 148220 659000
rect 148310 658760 148550 659000
rect 148640 658760 148880 659000
rect 148970 658760 149210 659000
rect 149320 658760 149560 659000
rect 149650 658760 149890 659000
rect 149980 658760 150220 659000
rect 150310 658760 150550 659000
rect 150660 658760 150900 659000
rect 150990 658760 151230 659000
rect 151320 658760 151560 659000
rect 151650 658760 151890 659000
rect 152000 658760 152240 659000
rect 152330 658760 152570 659000
rect 152660 658760 152900 659000
rect 152990 658760 153230 659000
rect 153340 658760 153580 659000
rect 153670 658760 153910 659000
rect 154000 658760 154240 659000
rect 154330 658760 154570 659000
rect 154680 658760 154920 659000
rect 155010 658760 155250 659000
rect 155340 658760 155580 659000
rect 155670 658760 155910 659000
rect 144950 658430 145190 658670
rect 145300 658430 145540 658670
rect 145630 658430 145870 658670
rect 145960 658430 146200 658670
rect 146290 658430 146530 658670
rect 146640 658430 146880 658670
rect 146970 658430 147210 658670
rect 147300 658430 147540 658670
rect 147630 658430 147870 658670
rect 147980 658430 148220 658670
rect 148310 658430 148550 658670
rect 148640 658430 148880 658670
rect 148970 658430 149210 658670
rect 149320 658430 149560 658670
rect 149650 658430 149890 658670
rect 149980 658430 150220 658670
rect 150310 658430 150550 658670
rect 150660 658430 150900 658670
rect 150990 658430 151230 658670
rect 151320 658430 151560 658670
rect 151650 658430 151890 658670
rect 152000 658430 152240 658670
rect 152330 658430 152570 658670
rect 152660 658430 152900 658670
rect 152990 658430 153230 658670
rect 153340 658430 153580 658670
rect 153670 658430 153910 658670
rect 154000 658430 154240 658670
rect 154330 658430 154570 658670
rect 154680 658430 154920 658670
rect 155010 658430 155250 658670
rect 155340 658430 155580 658670
rect 155670 658430 155910 658670
rect 144950 658100 145190 658340
rect 145300 658100 145540 658340
rect 145630 658100 145870 658340
rect 145960 658100 146200 658340
rect 146290 658100 146530 658340
rect 146640 658100 146880 658340
rect 146970 658100 147210 658340
rect 147300 658100 147540 658340
rect 147630 658100 147870 658340
rect 147980 658100 148220 658340
rect 148310 658100 148550 658340
rect 148640 658100 148880 658340
rect 148970 658100 149210 658340
rect 149320 658100 149560 658340
rect 149650 658100 149890 658340
rect 149980 658100 150220 658340
rect 150310 658100 150550 658340
rect 150660 658100 150900 658340
rect 150990 658100 151230 658340
rect 151320 658100 151560 658340
rect 151650 658100 151890 658340
rect 152000 658100 152240 658340
rect 152330 658100 152570 658340
rect 152660 658100 152900 658340
rect 152990 658100 153230 658340
rect 153340 658100 153580 658340
rect 153670 658100 153910 658340
rect 154000 658100 154240 658340
rect 154330 658100 154570 658340
rect 154680 658100 154920 658340
rect 155010 658100 155250 658340
rect 155340 658100 155580 658340
rect 155670 658100 155910 658340
rect 144950 657770 145190 658010
rect 145300 657770 145540 658010
rect 145630 657770 145870 658010
rect 145960 657770 146200 658010
rect 146290 657770 146530 658010
rect 146640 657770 146880 658010
rect 146970 657770 147210 658010
rect 147300 657770 147540 658010
rect 147630 657770 147870 658010
rect 147980 657770 148220 658010
rect 148310 657770 148550 658010
rect 148640 657770 148880 658010
rect 148970 657770 149210 658010
rect 149320 657770 149560 658010
rect 149650 657770 149890 658010
rect 149980 657770 150220 658010
rect 150310 657770 150550 658010
rect 150660 657770 150900 658010
rect 150990 657770 151230 658010
rect 151320 657770 151560 658010
rect 151650 657770 151890 658010
rect 152000 657770 152240 658010
rect 152330 657770 152570 658010
rect 152660 657770 152900 658010
rect 152990 657770 153230 658010
rect 153340 657770 153580 658010
rect 153670 657770 153910 658010
rect 154000 657770 154240 658010
rect 154330 657770 154570 658010
rect 154680 657770 154920 658010
rect 155010 657770 155250 658010
rect 155340 657770 155580 658010
rect 155670 657770 155910 658010
rect 144950 657420 145190 657660
rect 145300 657420 145540 657660
rect 145630 657420 145870 657660
rect 145960 657420 146200 657660
rect 146290 657420 146530 657660
rect 146640 657420 146880 657660
rect 146970 657420 147210 657660
rect 147300 657420 147540 657660
rect 147630 657420 147870 657660
rect 147980 657420 148220 657660
rect 148310 657420 148550 657660
rect 148640 657420 148880 657660
rect 148970 657420 149210 657660
rect 149320 657420 149560 657660
rect 149650 657420 149890 657660
rect 149980 657420 150220 657660
rect 150310 657420 150550 657660
rect 150660 657420 150900 657660
rect 150990 657420 151230 657660
rect 151320 657420 151560 657660
rect 151650 657420 151890 657660
rect 152000 657420 152240 657660
rect 152330 657420 152570 657660
rect 152660 657420 152900 657660
rect 152990 657420 153230 657660
rect 153340 657420 153580 657660
rect 153670 657420 153910 657660
rect 154000 657420 154240 657660
rect 154330 657420 154570 657660
rect 154680 657420 154920 657660
rect 155010 657420 155250 657660
rect 155340 657420 155580 657660
rect 155670 657420 155910 657660
rect 144950 657090 145190 657330
rect 145300 657090 145540 657330
rect 145630 657090 145870 657330
rect 145960 657090 146200 657330
rect 146290 657090 146530 657330
rect 146640 657090 146880 657330
rect 146970 657090 147210 657330
rect 147300 657090 147540 657330
rect 147630 657090 147870 657330
rect 147980 657090 148220 657330
rect 148310 657090 148550 657330
rect 148640 657090 148880 657330
rect 148970 657090 149210 657330
rect 149320 657090 149560 657330
rect 149650 657090 149890 657330
rect 149980 657090 150220 657330
rect 150310 657090 150550 657330
rect 150660 657090 150900 657330
rect 150990 657090 151230 657330
rect 151320 657090 151560 657330
rect 151650 657090 151890 657330
rect 152000 657090 152240 657330
rect 152330 657090 152570 657330
rect 152660 657090 152900 657330
rect 152990 657090 153230 657330
rect 153340 657090 153580 657330
rect 153670 657090 153910 657330
rect 154000 657090 154240 657330
rect 154330 657090 154570 657330
rect 154680 657090 154920 657330
rect 155010 657090 155250 657330
rect 155340 657090 155580 657330
rect 155670 657090 155910 657330
rect 144950 656760 145190 657000
rect 145300 656760 145540 657000
rect 145630 656760 145870 657000
rect 145960 656760 146200 657000
rect 146290 656760 146530 657000
rect 146640 656760 146880 657000
rect 146970 656760 147210 657000
rect 147300 656760 147540 657000
rect 147630 656760 147870 657000
rect 147980 656760 148220 657000
rect 148310 656760 148550 657000
rect 148640 656760 148880 657000
rect 148970 656760 149210 657000
rect 149320 656760 149560 657000
rect 149650 656760 149890 657000
rect 149980 656760 150220 657000
rect 150310 656760 150550 657000
rect 150660 656760 150900 657000
rect 150990 656760 151230 657000
rect 151320 656760 151560 657000
rect 151650 656760 151890 657000
rect 152000 656760 152240 657000
rect 152330 656760 152570 657000
rect 152660 656760 152900 657000
rect 152990 656760 153230 657000
rect 153340 656760 153580 657000
rect 153670 656760 153910 657000
rect 154000 656760 154240 657000
rect 154330 656760 154570 657000
rect 154680 656760 154920 657000
rect 155010 656760 155250 657000
rect 155340 656760 155580 657000
rect 155670 656760 155910 657000
rect 144950 656430 145190 656670
rect 145300 656430 145540 656670
rect 145630 656430 145870 656670
rect 145960 656430 146200 656670
rect 146290 656430 146530 656670
rect 146640 656430 146880 656670
rect 146970 656430 147210 656670
rect 147300 656430 147540 656670
rect 147630 656430 147870 656670
rect 147980 656430 148220 656670
rect 148310 656430 148550 656670
rect 148640 656430 148880 656670
rect 148970 656430 149210 656670
rect 149320 656430 149560 656670
rect 149650 656430 149890 656670
rect 149980 656430 150220 656670
rect 150310 656430 150550 656670
rect 150660 656430 150900 656670
rect 150990 656430 151230 656670
rect 151320 656430 151560 656670
rect 151650 656430 151890 656670
rect 152000 656430 152240 656670
rect 152330 656430 152570 656670
rect 152660 656430 152900 656670
rect 152990 656430 153230 656670
rect 153340 656430 153580 656670
rect 153670 656430 153910 656670
rect 154000 656430 154240 656670
rect 154330 656430 154570 656670
rect 154680 656430 154920 656670
rect 155010 656430 155250 656670
rect 155340 656430 155580 656670
rect 155670 656430 155910 656670
rect 144950 656080 145190 656320
rect 145300 656080 145540 656320
rect 145630 656080 145870 656320
rect 145960 656080 146200 656320
rect 146290 656080 146530 656320
rect 146640 656080 146880 656320
rect 146970 656080 147210 656320
rect 147300 656080 147540 656320
rect 147630 656080 147870 656320
rect 147980 656080 148220 656320
rect 148310 656080 148550 656320
rect 148640 656080 148880 656320
rect 148970 656080 149210 656320
rect 149320 656080 149560 656320
rect 149650 656080 149890 656320
rect 149980 656080 150220 656320
rect 150310 656080 150550 656320
rect 150660 656080 150900 656320
rect 150990 656080 151230 656320
rect 151320 656080 151560 656320
rect 151650 656080 151890 656320
rect 152000 656080 152240 656320
rect 152330 656080 152570 656320
rect 152660 656080 152900 656320
rect 152990 656080 153230 656320
rect 153340 656080 153580 656320
rect 153670 656080 153910 656320
rect 154000 656080 154240 656320
rect 154330 656080 154570 656320
rect 154680 656080 154920 656320
rect 155010 656080 155250 656320
rect 155340 656080 155580 656320
rect 155670 656080 155910 656320
rect 144950 655750 145190 655990
rect 145300 655750 145540 655990
rect 145630 655750 145870 655990
rect 145960 655750 146200 655990
rect 146290 655750 146530 655990
rect 146640 655750 146880 655990
rect 146970 655750 147210 655990
rect 147300 655750 147540 655990
rect 147630 655750 147870 655990
rect 147980 655750 148220 655990
rect 148310 655750 148550 655990
rect 148640 655750 148880 655990
rect 148970 655750 149210 655990
rect 149320 655750 149560 655990
rect 149650 655750 149890 655990
rect 149980 655750 150220 655990
rect 150310 655750 150550 655990
rect 150660 655750 150900 655990
rect 150990 655750 151230 655990
rect 151320 655750 151560 655990
rect 151650 655750 151890 655990
rect 152000 655750 152240 655990
rect 152330 655750 152570 655990
rect 152660 655750 152900 655990
rect 152990 655750 153230 655990
rect 153340 655750 153580 655990
rect 153670 655750 153910 655990
rect 154000 655750 154240 655990
rect 154330 655750 154570 655990
rect 154680 655750 154920 655990
rect 155010 655750 155250 655990
rect 155340 655750 155580 655990
rect 155670 655750 155910 655990
rect 144950 655420 145190 655660
rect 145300 655420 145540 655660
rect 145630 655420 145870 655660
rect 145960 655420 146200 655660
rect 146290 655420 146530 655660
rect 146640 655420 146880 655660
rect 146970 655420 147210 655660
rect 147300 655420 147540 655660
rect 147630 655420 147870 655660
rect 147980 655420 148220 655660
rect 148310 655420 148550 655660
rect 148640 655420 148880 655660
rect 148970 655420 149210 655660
rect 149320 655420 149560 655660
rect 149650 655420 149890 655660
rect 149980 655420 150220 655660
rect 150310 655420 150550 655660
rect 150660 655420 150900 655660
rect 150990 655420 151230 655660
rect 151320 655420 151560 655660
rect 151650 655420 151890 655660
rect 152000 655420 152240 655660
rect 152330 655420 152570 655660
rect 152660 655420 152900 655660
rect 152990 655420 153230 655660
rect 153340 655420 153580 655660
rect 153670 655420 153910 655660
rect 154000 655420 154240 655660
rect 154330 655420 154570 655660
rect 154680 655420 154920 655660
rect 155010 655420 155250 655660
rect 155340 655420 155580 655660
rect 155670 655420 155910 655660
rect 144950 655090 145190 655330
rect 145300 655090 145540 655330
rect 145630 655090 145870 655330
rect 145960 655090 146200 655330
rect 146290 655090 146530 655330
rect 146640 655090 146880 655330
rect 146970 655090 147210 655330
rect 147300 655090 147540 655330
rect 147630 655090 147870 655330
rect 147980 655090 148220 655330
rect 148310 655090 148550 655330
rect 148640 655090 148880 655330
rect 148970 655090 149210 655330
rect 149320 655090 149560 655330
rect 149650 655090 149890 655330
rect 149980 655090 150220 655330
rect 150310 655090 150550 655330
rect 150660 655090 150900 655330
rect 150990 655090 151230 655330
rect 151320 655090 151560 655330
rect 151650 655090 151890 655330
rect 152000 655090 152240 655330
rect 152330 655090 152570 655330
rect 152660 655090 152900 655330
rect 152990 655090 153230 655330
rect 153340 655090 153580 655330
rect 153670 655090 153910 655330
rect 154000 655090 154240 655330
rect 154330 655090 154570 655330
rect 154680 655090 154920 655330
rect 155010 655090 155250 655330
rect 155340 655090 155580 655330
rect 155670 655090 155910 655330
rect 144950 654740 145190 654980
rect 145300 654740 145540 654980
rect 145630 654740 145870 654980
rect 145960 654740 146200 654980
rect 146290 654740 146530 654980
rect 146640 654740 146880 654980
rect 146970 654740 147210 654980
rect 147300 654740 147540 654980
rect 147630 654740 147870 654980
rect 147980 654740 148220 654980
rect 148310 654740 148550 654980
rect 148640 654740 148880 654980
rect 148970 654740 149210 654980
rect 149320 654740 149560 654980
rect 149650 654740 149890 654980
rect 149980 654740 150220 654980
rect 150310 654740 150550 654980
rect 150660 654740 150900 654980
rect 150990 654740 151230 654980
rect 151320 654740 151560 654980
rect 151650 654740 151890 654980
rect 152000 654740 152240 654980
rect 152330 654740 152570 654980
rect 152660 654740 152900 654980
rect 152990 654740 153230 654980
rect 153340 654740 153580 654980
rect 153670 654740 153910 654980
rect 154000 654740 154240 654980
rect 154330 654740 154570 654980
rect 154680 654740 154920 654980
rect 155010 654740 155250 654980
rect 155340 654740 155580 654980
rect 155670 654740 155910 654980
rect 144950 654410 145190 654650
rect 145300 654410 145540 654650
rect 145630 654410 145870 654650
rect 145960 654410 146200 654650
rect 146290 654410 146530 654650
rect 146640 654410 146880 654650
rect 146970 654410 147210 654650
rect 147300 654410 147540 654650
rect 147630 654410 147870 654650
rect 147980 654410 148220 654650
rect 148310 654410 148550 654650
rect 148640 654410 148880 654650
rect 148970 654410 149210 654650
rect 149320 654410 149560 654650
rect 149650 654410 149890 654650
rect 149980 654410 150220 654650
rect 150310 654410 150550 654650
rect 150660 654410 150900 654650
rect 150990 654410 151230 654650
rect 151320 654410 151560 654650
rect 151650 654410 151890 654650
rect 152000 654410 152240 654650
rect 152330 654410 152570 654650
rect 152660 654410 152900 654650
rect 152990 654410 153230 654650
rect 153340 654410 153580 654650
rect 153670 654410 153910 654650
rect 154000 654410 154240 654650
rect 154330 654410 154570 654650
rect 154680 654410 154920 654650
rect 155010 654410 155250 654650
rect 155340 654410 155580 654650
rect 155670 654410 155910 654650
rect 144950 654080 145190 654320
rect 145300 654080 145540 654320
rect 145630 654080 145870 654320
rect 145960 654080 146200 654320
rect 146290 654080 146530 654320
rect 146640 654080 146880 654320
rect 146970 654080 147210 654320
rect 147300 654080 147540 654320
rect 147630 654080 147870 654320
rect 147980 654080 148220 654320
rect 148310 654080 148550 654320
rect 148640 654080 148880 654320
rect 148970 654080 149210 654320
rect 149320 654080 149560 654320
rect 149650 654080 149890 654320
rect 149980 654080 150220 654320
rect 150310 654080 150550 654320
rect 150660 654080 150900 654320
rect 150990 654080 151230 654320
rect 151320 654080 151560 654320
rect 151650 654080 151890 654320
rect 152000 654080 152240 654320
rect 152330 654080 152570 654320
rect 152660 654080 152900 654320
rect 152990 654080 153230 654320
rect 153340 654080 153580 654320
rect 153670 654080 153910 654320
rect 154000 654080 154240 654320
rect 154330 654080 154570 654320
rect 154680 654080 154920 654320
rect 155010 654080 155250 654320
rect 155340 654080 155580 654320
rect 155670 654080 155910 654320
rect 144950 653750 145190 653990
rect 145300 653750 145540 653990
rect 145630 653750 145870 653990
rect 145960 653750 146200 653990
rect 146290 653750 146530 653990
rect 146640 653750 146880 653990
rect 146970 653750 147210 653990
rect 147300 653750 147540 653990
rect 147630 653750 147870 653990
rect 147980 653750 148220 653990
rect 148310 653750 148550 653990
rect 148640 653750 148880 653990
rect 148970 653750 149210 653990
rect 149320 653750 149560 653990
rect 149650 653750 149890 653990
rect 149980 653750 150220 653990
rect 150310 653750 150550 653990
rect 150660 653750 150900 653990
rect 150990 653750 151230 653990
rect 151320 653750 151560 653990
rect 151650 653750 151890 653990
rect 152000 653750 152240 653990
rect 152330 653750 152570 653990
rect 152660 653750 152900 653990
rect 152990 653750 153230 653990
rect 153340 653750 153580 653990
rect 153670 653750 153910 653990
rect 154000 653750 154240 653990
rect 154330 653750 154570 653990
rect 154680 653750 154920 653990
rect 155010 653750 155250 653990
rect 155340 653750 155580 653990
rect 155670 653750 155910 653990
rect 144950 653400 145190 653640
rect 145300 653400 145540 653640
rect 145630 653400 145870 653640
rect 145960 653400 146200 653640
rect 146290 653400 146530 653640
rect 146640 653400 146880 653640
rect 146970 653400 147210 653640
rect 147300 653400 147540 653640
rect 147630 653400 147870 653640
rect 147980 653400 148220 653640
rect 148310 653400 148550 653640
rect 148640 653400 148880 653640
rect 148970 653400 149210 653640
rect 149320 653400 149560 653640
rect 149650 653400 149890 653640
rect 149980 653400 150220 653640
rect 150310 653400 150550 653640
rect 150660 653400 150900 653640
rect 150990 653400 151230 653640
rect 151320 653400 151560 653640
rect 151650 653400 151890 653640
rect 152000 653400 152240 653640
rect 152330 653400 152570 653640
rect 152660 653400 152900 653640
rect 152990 653400 153230 653640
rect 153340 653400 153580 653640
rect 153670 653400 153910 653640
rect 154000 653400 154240 653640
rect 154330 653400 154570 653640
rect 154680 653400 154920 653640
rect 155010 653400 155250 653640
rect 155340 653400 155580 653640
rect 155670 653400 155910 653640
rect 144950 653070 145190 653310
rect 145300 653070 145540 653310
rect 145630 653070 145870 653310
rect 145960 653070 146200 653310
rect 146290 653070 146530 653310
rect 146640 653070 146880 653310
rect 146970 653070 147210 653310
rect 147300 653070 147540 653310
rect 147630 653070 147870 653310
rect 147980 653070 148220 653310
rect 148310 653070 148550 653310
rect 148640 653070 148880 653310
rect 148970 653070 149210 653310
rect 149320 653070 149560 653310
rect 149650 653070 149890 653310
rect 149980 653070 150220 653310
rect 150310 653070 150550 653310
rect 150660 653070 150900 653310
rect 150990 653070 151230 653310
rect 151320 653070 151560 653310
rect 151650 653070 151890 653310
rect 152000 653070 152240 653310
rect 152330 653070 152570 653310
rect 152660 653070 152900 653310
rect 152990 653070 153230 653310
rect 153340 653070 153580 653310
rect 153670 653070 153910 653310
rect 154000 653070 154240 653310
rect 154330 653070 154570 653310
rect 154680 653070 154920 653310
rect 155010 653070 155250 653310
rect 155340 653070 155580 653310
rect 155670 653070 155910 653310
rect 144950 652740 145190 652980
rect 145300 652740 145540 652980
rect 145630 652740 145870 652980
rect 145960 652740 146200 652980
rect 146290 652740 146530 652980
rect 146640 652740 146880 652980
rect 146970 652740 147210 652980
rect 147300 652740 147540 652980
rect 147630 652740 147870 652980
rect 147980 652740 148220 652980
rect 148310 652740 148550 652980
rect 148640 652740 148880 652980
rect 148970 652740 149210 652980
rect 149320 652740 149560 652980
rect 149650 652740 149890 652980
rect 149980 652740 150220 652980
rect 150310 652740 150550 652980
rect 150660 652740 150900 652980
rect 150990 652740 151230 652980
rect 151320 652740 151560 652980
rect 151650 652740 151890 652980
rect 152000 652740 152240 652980
rect 152330 652740 152570 652980
rect 152660 652740 152900 652980
rect 152990 652740 153230 652980
rect 153340 652740 153580 652980
rect 153670 652740 153910 652980
rect 154000 652740 154240 652980
rect 154330 652740 154570 652980
rect 154680 652740 154920 652980
rect 155010 652740 155250 652980
rect 155340 652740 155580 652980
rect 155670 652740 155910 652980
rect 144950 652410 145190 652650
rect 145300 652410 145540 652650
rect 145630 652410 145870 652650
rect 145960 652410 146200 652650
rect 146290 652410 146530 652650
rect 146640 652410 146880 652650
rect 146970 652410 147210 652650
rect 147300 652410 147540 652650
rect 147630 652410 147870 652650
rect 147980 652410 148220 652650
rect 148310 652410 148550 652650
rect 148640 652410 148880 652650
rect 148970 652410 149210 652650
rect 149320 652410 149560 652650
rect 149650 652410 149890 652650
rect 149980 652410 150220 652650
rect 150310 652410 150550 652650
rect 150660 652410 150900 652650
rect 150990 652410 151230 652650
rect 151320 652410 151560 652650
rect 151650 652410 151890 652650
rect 152000 652410 152240 652650
rect 152330 652410 152570 652650
rect 152660 652410 152900 652650
rect 152990 652410 153230 652650
rect 153340 652410 153580 652650
rect 153670 652410 153910 652650
rect 154000 652410 154240 652650
rect 154330 652410 154570 652650
rect 154680 652410 154920 652650
rect 155010 652410 155250 652650
rect 155340 652410 155580 652650
rect 155670 652410 155910 652650
rect 144950 652060 145190 652300
rect 145300 652060 145540 652300
rect 145630 652060 145870 652300
rect 145960 652060 146200 652300
rect 146290 652060 146530 652300
rect 146640 652060 146880 652300
rect 146970 652060 147210 652300
rect 147300 652060 147540 652300
rect 147630 652060 147870 652300
rect 147980 652060 148220 652300
rect 148310 652060 148550 652300
rect 148640 652060 148880 652300
rect 148970 652060 149210 652300
rect 149320 652060 149560 652300
rect 149650 652060 149890 652300
rect 149980 652060 150220 652300
rect 150310 652060 150550 652300
rect 150660 652060 150900 652300
rect 150990 652060 151230 652300
rect 151320 652060 151560 652300
rect 151650 652060 151890 652300
rect 152000 652060 152240 652300
rect 152330 652060 152570 652300
rect 152660 652060 152900 652300
rect 152990 652060 153230 652300
rect 153340 652060 153580 652300
rect 153670 652060 153910 652300
rect 154000 652060 154240 652300
rect 154330 652060 154570 652300
rect 154680 652060 154920 652300
rect 155010 652060 155250 652300
rect 155340 652060 155580 652300
rect 155670 652060 155910 652300
rect 144950 651730 145190 651970
rect 145300 651730 145540 651970
rect 145630 651730 145870 651970
rect 145960 651730 146200 651970
rect 146290 651730 146530 651970
rect 146640 651730 146880 651970
rect 146970 651730 147210 651970
rect 147300 651730 147540 651970
rect 147630 651730 147870 651970
rect 147980 651730 148220 651970
rect 148310 651730 148550 651970
rect 148640 651730 148880 651970
rect 148970 651730 149210 651970
rect 149320 651730 149560 651970
rect 149650 651730 149890 651970
rect 149980 651730 150220 651970
rect 150310 651730 150550 651970
rect 150660 651730 150900 651970
rect 150990 651730 151230 651970
rect 151320 651730 151560 651970
rect 151650 651730 151890 651970
rect 152000 651730 152240 651970
rect 152330 651730 152570 651970
rect 152660 651730 152900 651970
rect 152990 651730 153230 651970
rect 153340 651730 153580 651970
rect 153670 651730 153910 651970
rect 154000 651730 154240 651970
rect 154330 651730 154570 651970
rect 154680 651730 154920 651970
rect 155010 651730 155250 651970
rect 155340 651730 155580 651970
rect 155670 651730 155910 651970
rect 144950 651400 145190 651640
rect 145300 651400 145540 651640
rect 145630 651400 145870 651640
rect 145960 651400 146200 651640
rect 146290 651400 146530 651640
rect 146640 651400 146880 651640
rect 146970 651400 147210 651640
rect 147300 651400 147540 651640
rect 147630 651400 147870 651640
rect 147980 651400 148220 651640
rect 148310 651400 148550 651640
rect 148640 651400 148880 651640
rect 148970 651400 149210 651640
rect 149320 651400 149560 651640
rect 149650 651400 149890 651640
rect 149980 651400 150220 651640
rect 150310 651400 150550 651640
rect 150660 651400 150900 651640
rect 150990 651400 151230 651640
rect 151320 651400 151560 651640
rect 151650 651400 151890 651640
rect 152000 651400 152240 651640
rect 152330 651400 152570 651640
rect 152660 651400 152900 651640
rect 152990 651400 153230 651640
rect 153340 651400 153580 651640
rect 153670 651400 153910 651640
rect 154000 651400 154240 651640
rect 154330 651400 154570 651640
rect 154680 651400 154920 651640
rect 155010 651400 155250 651640
rect 155340 651400 155580 651640
rect 155670 651400 155910 651640
rect 144950 651070 145190 651310
rect 145300 651070 145540 651310
rect 145630 651070 145870 651310
rect 145960 651070 146200 651310
rect 146290 651070 146530 651310
rect 146640 651070 146880 651310
rect 146970 651070 147210 651310
rect 147300 651070 147540 651310
rect 147630 651070 147870 651310
rect 147980 651070 148220 651310
rect 148310 651070 148550 651310
rect 148640 651070 148880 651310
rect 148970 651070 149210 651310
rect 149320 651070 149560 651310
rect 149650 651070 149890 651310
rect 149980 651070 150220 651310
rect 150310 651070 150550 651310
rect 150660 651070 150900 651310
rect 150990 651070 151230 651310
rect 151320 651070 151560 651310
rect 151650 651070 151890 651310
rect 152000 651070 152240 651310
rect 152330 651070 152570 651310
rect 152660 651070 152900 651310
rect 152990 651070 153230 651310
rect 153340 651070 153580 651310
rect 153670 651070 153910 651310
rect 154000 651070 154240 651310
rect 154330 651070 154570 651310
rect 154680 651070 154920 651310
rect 155010 651070 155250 651310
rect 155340 651070 155580 651310
rect 155670 651070 155910 651310
rect 144950 650720 145190 650960
rect 145300 650720 145540 650960
rect 145630 650720 145870 650960
rect 145960 650720 146200 650960
rect 146290 650720 146530 650960
rect 146640 650720 146880 650960
rect 146970 650720 147210 650960
rect 147300 650720 147540 650960
rect 147630 650720 147870 650960
rect 147980 650720 148220 650960
rect 148310 650720 148550 650960
rect 148640 650720 148880 650960
rect 148970 650720 149210 650960
rect 149320 650720 149560 650960
rect 149650 650720 149890 650960
rect 149980 650720 150220 650960
rect 150310 650720 150550 650960
rect 150660 650720 150900 650960
rect 150990 650720 151230 650960
rect 151320 650720 151560 650960
rect 151650 650720 151890 650960
rect 152000 650720 152240 650960
rect 152330 650720 152570 650960
rect 152660 650720 152900 650960
rect 152990 650720 153230 650960
rect 153340 650720 153580 650960
rect 153670 650720 153910 650960
rect 154000 650720 154240 650960
rect 154330 650720 154570 650960
rect 154680 650720 154920 650960
rect 155010 650720 155250 650960
rect 155340 650720 155580 650960
rect 155670 650720 155910 650960
rect 144950 650390 145190 650630
rect 145300 650390 145540 650630
rect 145630 650390 145870 650630
rect 145960 650390 146200 650630
rect 146290 650390 146530 650630
rect 146640 650390 146880 650630
rect 146970 650390 147210 650630
rect 147300 650390 147540 650630
rect 147630 650390 147870 650630
rect 147980 650390 148220 650630
rect 148310 650390 148550 650630
rect 148640 650390 148880 650630
rect 148970 650390 149210 650630
rect 149320 650390 149560 650630
rect 149650 650390 149890 650630
rect 149980 650390 150220 650630
rect 150310 650390 150550 650630
rect 150660 650390 150900 650630
rect 150990 650390 151230 650630
rect 151320 650390 151560 650630
rect 151650 650390 151890 650630
rect 152000 650390 152240 650630
rect 152330 650390 152570 650630
rect 152660 650390 152900 650630
rect 152990 650390 153230 650630
rect 153340 650390 153580 650630
rect 153670 650390 153910 650630
rect 154000 650390 154240 650630
rect 154330 650390 154570 650630
rect 154680 650390 154920 650630
rect 155010 650390 155250 650630
rect 155340 650390 155580 650630
rect 155670 650390 155910 650630
rect 144950 650060 145190 650300
rect 145300 650060 145540 650300
rect 145630 650060 145870 650300
rect 145960 650060 146200 650300
rect 146290 650060 146530 650300
rect 146640 650060 146880 650300
rect 146970 650060 147210 650300
rect 147300 650060 147540 650300
rect 147630 650060 147870 650300
rect 147980 650060 148220 650300
rect 148310 650060 148550 650300
rect 148640 650060 148880 650300
rect 148970 650060 149210 650300
rect 149320 650060 149560 650300
rect 149650 650060 149890 650300
rect 149980 650060 150220 650300
rect 150310 650060 150550 650300
rect 150660 650060 150900 650300
rect 150990 650060 151230 650300
rect 151320 650060 151560 650300
rect 151650 650060 151890 650300
rect 152000 650060 152240 650300
rect 152330 650060 152570 650300
rect 152660 650060 152900 650300
rect 152990 650060 153230 650300
rect 153340 650060 153580 650300
rect 153670 650060 153910 650300
rect 154000 650060 154240 650300
rect 154330 650060 154570 650300
rect 154680 650060 154920 650300
rect 155010 650060 155250 650300
rect 155340 650060 155580 650300
rect 155670 650060 155910 650300
rect 144950 649730 145190 649970
rect 145300 649730 145540 649970
rect 145630 649730 145870 649970
rect 145960 649730 146200 649970
rect 146290 649730 146530 649970
rect 146640 649730 146880 649970
rect 146970 649730 147210 649970
rect 147300 649730 147540 649970
rect 147630 649730 147870 649970
rect 147980 649730 148220 649970
rect 148310 649730 148550 649970
rect 148640 649730 148880 649970
rect 148970 649730 149210 649970
rect 149320 649730 149560 649970
rect 149650 649730 149890 649970
rect 149980 649730 150220 649970
rect 150310 649730 150550 649970
rect 150660 649730 150900 649970
rect 150990 649730 151230 649970
rect 151320 649730 151560 649970
rect 151650 649730 151890 649970
rect 152000 649730 152240 649970
rect 152330 649730 152570 649970
rect 152660 649730 152900 649970
rect 152990 649730 153230 649970
rect 153340 649730 153580 649970
rect 153670 649730 153910 649970
rect 154000 649730 154240 649970
rect 154330 649730 154570 649970
rect 154680 649730 154920 649970
rect 155010 649730 155250 649970
rect 155340 649730 155580 649970
rect 155670 649730 155910 649970
rect 144950 649380 145190 649620
rect 145300 649380 145540 649620
rect 145630 649380 145870 649620
rect 145960 649380 146200 649620
rect 146290 649380 146530 649620
rect 146640 649380 146880 649620
rect 146970 649380 147210 649620
rect 147300 649380 147540 649620
rect 147630 649380 147870 649620
rect 147980 649380 148220 649620
rect 148310 649380 148550 649620
rect 148640 649380 148880 649620
rect 148970 649380 149210 649620
rect 149320 649380 149560 649620
rect 149650 649380 149890 649620
rect 149980 649380 150220 649620
rect 150310 649380 150550 649620
rect 150660 649380 150900 649620
rect 150990 649380 151230 649620
rect 151320 649380 151560 649620
rect 151650 649380 151890 649620
rect 152000 649380 152240 649620
rect 152330 649380 152570 649620
rect 152660 649380 152900 649620
rect 152990 649380 153230 649620
rect 153340 649380 153580 649620
rect 153670 649380 153910 649620
rect 154000 649380 154240 649620
rect 154330 649380 154570 649620
rect 154680 649380 154920 649620
rect 155010 649380 155250 649620
rect 155340 649380 155580 649620
rect 155670 649380 155910 649620
<< metal4 >>
rect 16194 703800 21194 704000
rect 16194 703500 16352 703800
rect 16652 703500 16852 703800
rect 17152 703500 17352 703800
rect 17652 703500 17852 703800
rect 18152 703500 18352 703800
rect 18652 703500 18852 703800
rect 19152 703500 19352 703800
rect 19652 703500 19852 703800
rect 20152 703500 20352 703800
rect 20652 703500 20852 703800
rect 21152 703500 21194 703800
rect 16194 703300 21194 703500
rect 16194 703000 16352 703300
rect 16652 703000 16852 703300
rect 17152 703000 17352 703300
rect 17652 703000 17852 703300
rect 18152 703000 18352 703300
rect 18652 703000 18852 703300
rect 19152 703000 19352 703300
rect 19652 703000 19852 703300
rect 20152 703000 20352 703300
rect 20652 703000 20852 703300
rect 21152 703000 21194 703300
rect 16194 702800 21194 703000
rect 16194 702500 16352 702800
rect 16652 702500 16852 702800
rect 17152 702500 17352 702800
rect 17652 702500 17852 702800
rect 18152 702500 18352 702800
rect 18652 702500 18852 702800
rect 19152 702500 19352 702800
rect 19652 702500 19852 702800
rect 20152 702500 20352 702800
rect 20652 702500 20852 702800
rect 21152 702500 21194 702800
rect 16194 697044 21194 702500
rect 70217 703200 71237 703371
rect 70217 703000 70300 703200
rect 70500 703000 70600 703200
rect 70800 703000 70900 703200
rect 71100 703000 71237 703200
rect 70217 702900 71237 703000
rect 70217 702700 70300 702900
rect 70500 702700 70600 702900
rect 70800 702700 70900 702900
rect 71100 702700 71237 702900
rect 70217 702600 71237 702700
rect 70217 702400 70300 702600
rect 70500 702400 70600 702600
rect 70800 702400 70900 702600
rect 71100 702400 71237 702600
rect 70217 701358 71237 702400
rect 122042 703194 123062 703365
rect 122042 702994 122179 703194
rect 122379 702994 122479 703194
rect 122679 702994 122779 703194
rect 122979 702994 123062 703194
rect 122042 702894 123062 702994
rect 122042 702694 122179 702894
rect 122379 702694 122479 702894
rect 122679 702694 122779 702894
rect 122979 702694 123062 702894
rect 122042 702594 123062 702694
rect 122042 702394 122179 702594
rect 122379 702394 122479 702594
rect 122679 702394 122779 702594
rect 122979 702394 123062 702594
rect 70217 700338 95358 701358
rect 122042 701352 123062 702394
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 467200 703310 467520 703330
rect 467200 703240 467220 703310
rect 467290 703240 467320 703310
rect 467390 703240 467420 703310
rect 467490 703240 467520 703310
rect 467200 703220 467520 703240
rect 415740 703110 416220 703170
rect 415740 703040 415760 703110
rect 415830 703040 415850 703110
rect 415920 703040 415940 703110
rect 416010 703040 416030 703110
rect 416100 703040 416120 703110
rect 416190 703040 416220 703110
rect 415740 703020 416220 703040
rect 415740 702950 415760 703020
rect 415830 702950 415850 703020
rect 415920 702950 415940 703020
rect 416010 702950 416030 703020
rect 416100 702950 416120 703020
rect 416190 702950 416220 703020
rect 415740 702930 416220 702950
rect 415740 702860 415760 702930
rect 415830 702860 415850 702930
rect 415920 702860 415940 702930
rect 416010 702860 416030 702930
rect 416100 702860 416120 702930
rect 416190 702860 416220 702930
rect 415740 702840 416220 702860
rect 415740 702770 415760 702840
rect 415830 702770 415850 702840
rect 415920 702770 415940 702840
rect 416010 702770 416030 702840
rect 416100 702770 416120 702840
rect 416190 702770 416220 702840
rect 415740 702750 416220 702770
rect 415740 702680 415760 702750
rect 415830 702680 415850 702750
rect 415920 702680 415940 702750
rect 416010 702680 416030 702750
rect 416100 702680 416120 702750
rect 416190 702680 416220 702750
rect 0 685200 2500 685242
rect 0 684900 200 685200
rect 500 684900 700 685200
rect 1000 684900 1200 685200
rect 1500 684900 2500 685200
rect 0 684700 2500 684900
rect 0 684400 200 684700
rect 500 684400 700 684700
rect 1000 684400 1200 684700
rect 1500 684400 2500 684700
rect 0 684200 2500 684400
rect 0 683900 200 684200
rect 500 683900 700 684200
rect 1000 683900 1200 684200
rect 1500 683900 2500 684200
rect 0 683700 2500 683900
rect 0 683400 200 683700
rect 500 683400 700 683700
rect 1000 683400 1200 683700
rect 1500 683400 2500 683700
rect 0 683200 2500 683400
rect 0 682900 200 683200
rect 500 682900 700 683200
rect 1000 682900 1200 683200
rect 1500 682900 2500 683200
rect 0 682700 2500 682900
rect 0 682400 200 682700
rect 500 682400 700 682700
rect 1000 682400 1200 682700
rect 1500 682400 2500 682700
rect 0 682200 2500 682400
rect 0 681900 200 682200
rect 500 681900 700 682200
rect 1000 681900 1200 682200
rect 1500 681900 2500 682200
rect 0 681700 2500 681900
rect 0 681400 200 681700
rect 500 681400 700 681700
rect 1000 681400 1200 681700
rect 1500 681400 2500 681700
rect 0 681200 2500 681400
rect 0 680900 200 681200
rect 500 680900 700 681200
rect 1000 680900 1200 681200
rect 1500 680900 2500 681200
rect 0 680700 2500 680900
rect 0 680400 200 680700
rect 500 680400 700 680700
rect 1000 680400 1200 680700
rect 1500 680400 2500 680700
rect 0 680242 2500 680400
rect 94338 643561 95358 700338
rect 98509 700332 123062 701352
rect 98509 645944 99529 700332
rect 110760 694840 155960 694890
rect 110760 694600 110810 694840
rect 111050 694600 111140 694840
rect 111380 694600 111470 694840
rect 111710 694600 111800 694840
rect 112040 694600 112150 694840
rect 112390 694600 112480 694840
rect 112720 694600 112810 694840
rect 113050 694600 113140 694840
rect 113380 694600 113490 694840
rect 113730 694600 113820 694840
rect 114060 694600 114150 694840
rect 114390 694600 114480 694840
rect 114720 694600 114830 694840
rect 115070 694600 115160 694840
rect 115400 694600 115490 694840
rect 115730 694600 115820 694840
rect 116060 694600 116170 694840
rect 116410 694600 116500 694840
rect 116740 694600 116830 694840
rect 117070 694600 117160 694840
rect 117400 694600 117510 694840
rect 117750 694600 117840 694840
rect 118080 694600 118170 694840
rect 118410 694600 118500 694840
rect 118740 694600 118850 694840
rect 119090 694600 119180 694840
rect 119420 694600 119510 694840
rect 119750 694600 119840 694840
rect 120080 694600 120190 694840
rect 120430 694600 120520 694840
rect 120760 694600 120850 694840
rect 121090 694600 121180 694840
rect 121420 694600 121530 694840
rect 121770 694600 122190 694840
rect 122430 694600 122520 694840
rect 122760 694600 122850 694840
rect 123090 694600 123180 694840
rect 123420 694600 123530 694840
rect 123770 694600 123860 694840
rect 124100 694600 124190 694840
rect 124430 694600 124520 694840
rect 124760 694600 124870 694840
rect 125110 694600 125200 694840
rect 125440 694600 125530 694840
rect 125770 694600 125860 694840
rect 126100 694600 126210 694840
rect 126450 694600 126540 694840
rect 126780 694600 126870 694840
rect 127110 694600 127200 694840
rect 127440 694600 127550 694840
rect 127790 694600 127880 694840
rect 128120 694600 128210 694840
rect 128450 694600 128540 694840
rect 128780 694600 128890 694840
rect 129130 694600 129220 694840
rect 129460 694600 129550 694840
rect 129790 694600 129880 694840
rect 130120 694600 130230 694840
rect 130470 694600 130560 694840
rect 130800 694600 130890 694840
rect 131130 694600 131220 694840
rect 131460 694600 131570 694840
rect 131810 694600 131900 694840
rect 132140 694600 132230 694840
rect 132470 694600 132560 694840
rect 132800 694600 132910 694840
rect 133150 694600 133570 694840
rect 133810 694600 133900 694840
rect 134140 694600 134230 694840
rect 134470 694600 134560 694840
rect 134800 694600 134910 694840
rect 135150 694600 135240 694840
rect 135480 694600 135570 694840
rect 135810 694600 135900 694840
rect 136140 694600 136250 694840
rect 136490 694600 136580 694840
rect 136820 694600 136910 694840
rect 137150 694600 137240 694840
rect 137480 694600 137590 694840
rect 137830 694600 137920 694840
rect 138160 694600 138250 694840
rect 138490 694600 138580 694840
rect 138820 694600 138930 694840
rect 139170 694600 139260 694840
rect 139500 694600 139590 694840
rect 139830 694600 139920 694840
rect 140160 694600 140270 694840
rect 140510 694600 140600 694840
rect 140840 694600 140930 694840
rect 141170 694600 141260 694840
rect 141500 694600 141610 694840
rect 141850 694600 141940 694840
rect 142180 694600 142270 694840
rect 142510 694600 142600 694840
rect 142840 694600 142950 694840
rect 143190 694600 143280 694840
rect 143520 694600 143610 694840
rect 143850 694600 143940 694840
rect 144180 694600 144290 694840
rect 144530 694600 144950 694840
rect 145190 694600 145280 694840
rect 145520 694600 145610 694840
rect 145850 694600 145940 694840
rect 146180 694600 146290 694840
rect 146530 694600 146620 694840
rect 146860 694600 146950 694840
rect 147190 694600 147280 694840
rect 147520 694600 147630 694840
rect 147870 694600 147960 694840
rect 148200 694600 148290 694840
rect 148530 694600 148620 694840
rect 148860 694600 148970 694840
rect 149210 694600 149300 694840
rect 149540 694600 149630 694840
rect 149870 694600 149960 694840
rect 150200 694600 150310 694840
rect 150550 694600 150640 694840
rect 150880 694600 150970 694840
rect 151210 694600 151300 694840
rect 151540 694600 151650 694840
rect 151890 694600 151980 694840
rect 152220 694600 152310 694840
rect 152550 694600 152640 694840
rect 152880 694600 152990 694840
rect 153230 694600 153320 694840
rect 153560 694600 153650 694840
rect 153890 694600 153980 694840
rect 154220 694600 154330 694840
rect 154570 694600 154660 694840
rect 154900 694600 154990 694840
rect 155230 694600 155320 694840
rect 155560 694600 155670 694840
rect 155910 694600 155960 694840
rect 110760 694490 155960 694600
rect 110760 694250 110810 694490
rect 111050 694250 111140 694490
rect 111380 694250 111470 694490
rect 111710 694250 111800 694490
rect 112040 694250 112150 694490
rect 112390 694250 112480 694490
rect 112720 694250 112810 694490
rect 113050 694250 113140 694490
rect 113380 694250 113490 694490
rect 113730 694250 113820 694490
rect 114060 694250 114150 694490
rect 114390 694250 114480 694490
rect 114720 694250 114830 694490
rect 115070 694250 115160 694490
rect 115400 694250 115490 694490
rect 115730 694250 115820 694490
rect 116060 694250 116170 694490
rect 116410 694250 116500 694490
rect 116740 694250 116830 694490
rect 117070 694250 117160 694490
rect 117400 694250 117510 694490
rect 117750 694250 117840 694490
rect 118080 694250 118170 694490
rect 118410 694250 118500 694490
rect 118740 694250 118850 694490
rect 119090 694250 119180 694490
rect 119420 694250 119510 694490
rect 119750 694250 119840 694490
rect 120080 694250 120190 694490
rect 120430 694250 120520 694490
rect 120760 694250 120850 694490
rect 121090 694250 121180 694490
rect 121420 694250 121530 694490
rect 121770 694250 122190 694490
rect 122430 694250 122520 694490
rect 122760 694250 122850 694490
rect 123090 694250 123180 694490
rect 123420 694250 123530 694490
rect 123770 694250 123860 694490
rect 124100 694250 124190 694490
rect 124430 694250 124520 694490
rect 124760 694250 124870 694490
rect 125110 694250 125200 694490
rect 125440 694250 125530 694490
rect 125770 694250 125860 694490
rect 126100 694250 126210 694490
rect 126450 694250 126540 694490
rect 126780 694250 126870 694490
rect 127110 694250 127200 694490
rect 127440 694250 127550 694490
rect 127790 694250 127880 694490
rect 128120 694250 128210 694490
rect 128450 694250 128540 694490
rect 128780 694250 128890 694490
rect 129130 694250 129220 694490
rect 129460 694250 129550 694490
rect 129790 694250 129880 694490
rect 130120 694250 130230 694490
rect 130470 694250 130560 694490
rect 130800 694250 130890 694490
rect 131130 694250 131220 694490
rect 131460 694250 131570 694490
rect 131810 694250 131900 694490
rect 132140 694250 132230 694490
rect 132470 694250 132560 694490
rect 132800 694250 132910 694490
rect 133150 694250 133570 694490
rect 133810 694250 133900 694490
rect 134140 694250 134230 694490
rect 134470 694250 134560 694490
rect 134800 694250 134910 694490
rect 135150 694250 135240 694490
rect 135480 694250 135570 694490
rect 135810 694250 135900 694490
rect 136140 694250 136250 694490
rect 136490 694250 136580 694490
rect 136820 694250 136910 694490
rect 137150 694250 137240 694490
rect 137480 694250 137590 694490
rect 137830 694250 137920 694490
rect 138160 694250 138250 694490
rect 138490 694250 138580 694490
rect 138820 694250 138930 694490
rect 139170 694250 139260 694490
rect 139500 694250 139590 694490
rect 139830 694250 139920 694490
rect 140160 694250 140270 694490
rect 140510 694250 140600 694490
rect 140840 694250 140930 694490
rect 141170 694250 141260 694490
rect 141500 694250 141610 694490
rect 141850 694250 141940 694490
rect 142180 694250 142270 694490
rect 142510 694250 142600 694490
rect 142840 694250 142950 694490
rect 143190 694250 143280 694490
rect 143520 694250 143610 694490
rect 143850 694250 143940 694490
rect 144180 694250 144290 694490
rect 144530 694250 144950 694490
rect 145190 694250 145280 694490
rect 145520 694250 145610 694490
rect 145850 694250 145940 694490
rect 146180 694250 146290 694490
rect 146530 694250 146620 694490
rect 146860 694250 146950 694490
rect 147190 694250 147280 694490
rect 147520 694250 147630 694490
rect 147870 694250 147960 694490
rect 148200 694250 148290 694490
rect 148530 694250 148620 694490
rect 148860 694250 148970 694490
rect 149210 694250 149300 694490
rect 149540 694250 149630 694490
rect 149870 694250 149960 694490
rect 150200 694250 150310 694490
rect 150550 694250 150640 694490
rect 150880 694250 150970 694490
rect 151210 694250 151300 694490
rect 151540 694250 151650 694490
rect 151890 694250 151980 694490
rect 152220 694250 152310 694490
rect 152550 694250 152640 694490
rect 152880 694250 152990 694490
rect 153230 694250 153320 694490
rect 153560 694250 153650 694490
rect 153890 694250 153980 694490
rect 154220 694250 154330 694490
rect 154570 694250 154660 694490
rect 154900 694250 154990 694490
rect 155230 694250 155320 694490
rect 155560 694250 155670 694490
rect 155910 694250 155960 694490
rect 110760 694160 155960 694250
rect 110760 693920 110810 694160
rect 111050 693920 111140 694160
rect 111380 693920 111470 694160
rect 111710 693920 111800 694160
rect 112040 693920 112150 694160
rect 112390 693920 112480 694160
rect 112720 693920 112810 694160
rect 113050 693920 113140 694160
rect 113380 693920 113490 694160
rect 113730 693920 113820 694160
rect 114060 693920 114150 694160
rect 114390 693920 114480 694160
rect 114720 693920 114830 694160
rect 115070 693920 115160 694160
rect 115400 693920 115490 694160
rect 115730 693920 115820 694160
rect 116060 693920 116170 694160
rect 116410 693920 116500 694160
rect 116740 693920 116830 694160
rect 117070 693920 117160 694160
rect 117400 693920 117510 694160
rect 117750 693920 117840 694160
rect 118080 693920 118170 694160
rect 118410 693920 118500 694160
rect 118740 693920 118850 694160
rect 119090 693920 119180 694160
rect 119420 693920 119510 694160
rect 119750 693920 119840 694160
rect 120080 693920 120190 694160
rect 120430 693920 120520 694160
rect 120760 693920 120850 694160
rect 121090 693920 121180 694160
rect 121420 693920 121530 694160
rect 121770 693920 122190 694160
rect 122430 693920 122520 694160
rect 122760 693920 122850 694160
rect 123090 693920 123180 694160
rect 123420 693920 123530 694160
rect 123770 693920 123860 694160
rect 124100 693920 124190 694160
rect 124430 693920 124520 694160
rect 124760 693920 124870 694160
rect 125110 693920 125200 694160
rect 125440 693920 125530 694160
rect 125770 693920 125860 694160
rect 126100 693920 126210 694160
rect 126450 693920 126540 694160
rect 126780 693920 126870 694160
rect 127110 693920 127200 694160
rect 127440 693920 127550 694160
rect 127790 693920 127880 694160
rect 128120 693920 128210 694160
rect 128450 693920 128540 694160
rect 128780 693920 128890 694160
rect 129130 693920 129220 694160
rect 129460 693920 129550 694160
rect 129790 693920 129880 694160
rect 130120 693920 130230 694160
rect 130470 693920 130560 694160
rect 130800 693920 130890 694160
rect 131130 693920 131220 694160
rect 131460 693920 131570 694160
rect 131810 693920 131900 694160
rect 132140 693920 132230 694160
rect 132470 693920 132560 694160
rect 132800 693920 132910 694160
rect 133150 693920 133570 694160
rect 133810 693920 133900 694160
rect 134140 693920 134230 694160
rect 134470 693920 134560 694160
rect 134800 693920 134910 694160
rect 135150 693920 135240 694160
rect 135480 693920 135570 694160
rect 135810 693920 135900 694160
rect 136140 693920 136250 694160
rect 136490 693920 136580 694160
rect 136820 693920 136910 694160
rect 137150 693920 137240 694160
rect 137480 693920 137590 694160
rect 137830 693920 137920 694160
rect 138160 693920 138250 694160
rect 138490 693920 138580 694160
rect 138820 693920 138930 694160
rect 139170 693920 139260 694160
rect 139500 693920 139590 694160
rect 139830 693920 139920 694160
rect 140160 693920 140270 694160
rect 140510 693920 140600 694160
rect 140840 693920 140930 694160
rect 141170 693920 141260 694160
rect 141500 693920 141610 694160
rect 141850 693920 141940 694160
rect 142180 693920 142270 694160
rect 142510 693920 142600 694160
rect 142840 693920 142950 694160
rect 143190 693920 143280 694160
rect 143520 693920 143610 694160
rect 143850 693920 143940 694160
rect 144180 693920 144290 694160
rect 144530 693920 144950 694160
rect 145190 693920 145280 694160
rect 145520 693920 145610 694160
rect 145850 693920 145940 694160
rect 146180 693920 146290 694160
rect 146530 693920 146620 694160
rect 146860 693920 146950 694160
rect 147190 693920 147280 694160
rect 147520 693920 147630 694160
rect 147870 693920 147960 694160
rect 148200 693920 148290 694160
rect 148530 693920 148620 694160
rect 148860 693920 148970 694160
rect 149210 693920 149300 694160
rect 149540 693920 149630 694160
rect 149870 693920 149960 694160
rect 150200 693920 150310 694160
rect 150550 693920 150640 694160
rect 150880 693920 150970 694160
rect 151210 693920 151300 694160
rect 151540 693920 151650 694160
rect 151890 693920 151980 694160
rect 152220 693920 152310 694160
rect 152550 693920 152640 694160
rect 152880 693920 152990 694160
rect 153230 693920 153320 694160
rect 153560 693920 153650 694160
rect 153890 693920 153980 694160
rect 154220 693920 154330 694160
rect 154570 693920 154660 694160
rect 154900 693920 154990 694160
rect 155230 693920 155320 694160
rect 155560 693920 155670 694160
rect 155910 693920 155960 694160
rect 110760 693830 155960 693920
rect 110760 693590 110810 693830
rect 111050 693590 111140 693830
rect 111380 693590 111470 693830
rect 111710 693590 111800 693830
rect 112040 693590 112150 693830
rect 112390 693590 112480 693830
rect 112720 693590 112810 693830
rect 113050 693590 113140 693830
rect 113380 693590 113490 693830
rect 113730 693590 113820 693830
rect 114060 693590 114150 693830
rect 114390 693590 114480 693830
rect 114720 693590 114830 693830
rect 115070 693590 115160 693830
rect 115400 693590 115490 693830
rect 115730 693590 115820 693830
rect 116060 693590 116170 693830
rect 116410 693590 116500 693830
rect 116740 693590 116830 693830
rect 117070 693590 117160 693830
rect 117400 693590 117510 693830
rect 117750 693590 117840 693830
rect 118080 693590 118170 693830
rect 118410 693590 118500 693830
rect 118740 693590 118850 693830
rect 119090 693590 119180 693830
rect 119420 693590 119510 693830
rect 119750 693590 119840 693830
rect 120080 693590 120190 693830
rect 120430 693590 120520 693830
rect 120760 693590 120850 693830
rect 121090 693590 121180 693830
rect 121420 693590 121530 693830
rect 121770 693590 122190 693830
rect 122430 693590 122520 693830
rect 122760 693590 122850 693830
rect 123090 693590 123180 693830
rect 123420 693590 123530 693830
rect 123770 693590 123860 693830
rect 124100 693590 124190 693830
rect 124430 693590 124520 693830
rect 124760 693590 124870 693830
rect 125110 693590 125200 693830
rect 125440 693590 125530 693830
rect 125770 693590 125860 693830
rect 126100 693590 126210 693830
rect 126450 693590 126540 693830
rect 126780 693590 126870 693830
rect 127110 693590 127200 693830
rect 127440 693590 127550 693830
rect 127790 693590 127880 693830
rect 128120 693590 128210 693830
rect 128450 693590 128540 693830
rect 128780 693590 128890 693830
rect 129130 693590 129220 693830
rect 129460 693590 129550 693830
rect 129790 693590 129880 693830
rect 130120 693590 130230 693830
rect 130470 693590 130560 693830
rect 130800 693590 130890 693830
rect 131130 693590 131220 693830
rect 131460 693590 131570 693830
rect 131810 693590 131900 693830
rect 132140 693590 132230 693830
rect 132470 693590 132560 693830
rect 132800 693590 132910 693830
rect 133150 693590 133570 693830
rect 133810 693590 133900 693830
rect 134140 693590 134230 693830
rect 134470 693590 134560 693830
rect 134800 693590 134910 693830
rect 135150 693590 135240 693830
rect 135480 693590 135570 693830
rect 135810 693590 135900 693830
rect 136140 693590 136250 693830
rect 136490 693590 136580 693830
rect 136820 693590 136910 693830
rect 137150 693590 137240 693830
rect 137480 693590 137590 693830
rect 137830 693590 137920 693830
rect 138160 693590 138250 693830
rect 138490 693590 138580 693830
rect 138820 693590 138930 693830
rect 139170 693590 139260 693830
rect 139500 693590 139590 693830
rect 139830 693590 139920 693830
rect 140160 693590 140270 693830
rect 140510 693590 140600 693830
rect 140840 693590 140930 693830
rect 141170 693590 141260 693830
rect 141500 693590 141610 693830
rect 141850 693590 141940 693830
rect 142180 693590 142270 693830
rect 142510 693590 142600 693830
rect 142840 693590 142950 693830
rect 143190 693590 143280 693830
rect 143520 693590 143610 693830
rect 143850 693590 143940 693830
rect 144180 693590 144290 693830
rect 144530 693590 144950 693830
rect 145190 693590 145280 693830
rect 145520 693590 145610 693830
rect 145850 693590 145940 693830
rect 146180 693590 146290 693830
rect 146530 693590 146620 693830
rect 146860 693590 146950 693830
rect 147190 693590 147280 693830
rect 147520 693590 147630 693830
rect 147870 693590 147960 693830
rect 148200 693590 148290 693830
rect 148530 693590 148620 693830
rect 148860 693590 148970 693830
rect 149210 693590 149300 693830
rect 149540 693590 149630 693830
rect 149870 693590 149960 693830
rect 150200 693590 150310 693830
rect 150550 693590 150640 693830
rect 150880 693590 150970 693830
rect 151210 693590 151300 693830
rect 151540 693590 151650 693830
rect 151890 693590 151980 693830
rect 152220 693590 152310 693830
rect 152550 693590 152640 693830
rect 152880 693590 152990 693830
rect 153230 693590 153320 693830
rect 153560 693590 153650 693830
rect 153890 693590 153980 693830
rect 154220 693590 154330 693830
rect 154570 693590 154660 693830
rect 154900 693590 154990 693830
rect 155230 693590 155320 693830
rect 155560 693590 155670 693830
rect 155910 693590 155960 693830
rect 110760 693500 155960 693590
rect 110760 693260 110810 693500
rect 111050 693260 111140 693500
rect 111380 693260 111470 693500
rect 111710 693260 111800 693500
rect 112040 693260 112150 693500
rect 112390 693260 112480 693500
rect 112720 693260 112810 693500
rect 113050 693260 113140 693500
rect 113380 693260 113490 693500
rect 113730 693260 113820 693500
rect 114060 693260 114150 693500
rect 114390 693260 114480 693500
rect 114720 693260 114830 693500
rect 115070 693260 115160 693500
rect 115400 693260 115490 693500
rect 115730 693260 115820 693500
rect 116060 693260 116170 693500
rect 116410 693260 116500 693500
rect 116740 693260 116830 693500
rect 117070 693260 117160 693500
rect 117400 693260 117510 693500
rect 117750 693260 117840 693500
rect 118080 693260 118170 693500
rect 118410 693260 118500 693500
rect 118740 693260 118850 693500
rect 119090 693260 119180 693500
rect 119420 693260 119510 693500
rect 119750 693260 119840 693500
rect 120080 693260 120190 693500
rect 120430 693260 120520 693500
rect 120760 693260 120850 693500
rect 121090 693260 121180 693500
rect 121420 693260 121530 693500
rect 121770 693260 122190 693500
rect 122430 693260 122520 693500
rect 122760 693260 122850 693500
rect 123090 693260 123180 693500
rect 123420 693260 123530 693500
rect 123770 693260 123860 693500
rect 124100 693260 124190 693500
rect 124430 693260 124520 693500
rect 124760 693260 124870 693500
rect 125110 693260 125200 693500
rect 125440 693260 125530 693500
rect 125770 693260 125860 693500
rect 126100 693260 126210 693500
rect 126450 693260 126540 693500
rect 126780 693260 126870 693500
rect 127110 693260 127200 693500
rect 127440 693260 127550 693500
rect 127790 693260 127880 693500
rect 128120 693260 128210 693500
rect 128450 693260 128540 693500
rect 128780 693260 128890 693500
rect 129130 693260 129220 693500
rect 129460 693260 129550 693500
rect 129790 693260 129880 693500
rect 130120 693260 130230 693500
rect 130470 693260 130560 693500
rect 130800 693260 130890 693500
rect 131130 693260 131220 693500
rect 131460 693260 131570 693500
rect 131810 693260 131900 693500
rect 132140 693260 132230 693500
rect 132470 693260 132560 693500
rect 132800 693260 132910 693500
rect 133150 693260 133570 693500
rect 133810 693260 133900 693500
rect 134140 693260 134230 693500
rect 134470 693260 134560 693500
rect 134800 693260 134910 693500
rect 135150 693260 135240 693500
rect 135480 693260 135570 693500
rect 135810 693260 135900 693500
rect 136140 693260 136250 693500
rect 136490 693260 136580 693500
rect 136820 693260 136910 693500
rect 137150 693260 137240 693500
rect 137480 693260 137590 693500
rect 137830 693260 137920 693500
rect 138160 693260 138250 693500
rect 138490 693260 138580 693500
rect 138820 693260 138930 693500
rect 139170 693260 139260 693500
rect 139500 693260 139590 693500
rect 139830 693260 139920 693500
rect 140160 693260 140270 693500
rect 140510 693260 140600 693500
rect 140840 693260 140930 693500
rect 141170 693260 141260 693500
rect 141500 693260 141610 693500
rect 141850 693260 141940 693500
rect 142180 693260 142270 693500
rect 142510 693260 142600 693500
rect 142840 693260 142950 693500
rect 143190 693260 143280 693500
rect 143520 693260 143610 693500
rect 143850 693260 143940 693500
rect 144180 693260 144290 693500
rect 144530 693260 144950 693500
rect 145190 693260 145280 693500
rect 145520 693260 145610 693500
rect 145850 693260 145940 693500
rect 146180 693260 146290 693500
rect 146530 693260 146620 693500
rect 146860 693260 146950 693500
rect 147190 693260 147280 693500
rect 147520 693260 147630 693500
rect 147870 693260 147960 693500
rect 148200 693260 148290 693500
rect 148530 693260 148620 693500
rect 148860 693260 148970 693500
rect 149210 693260 149300 693500
rect 149540 693260 149630 693500
rect 149870 693260 149960 693500
rect 150200 693260 150310 693500
rect 150550 693260 150640 693500
rect 150880 693260 150970 693500
rect 151210 693260 151300 693500
rect 151540 693260 151650 693500
rect 151890 693260 151980 693500
rect 152220 693260 152310 693500
rect 152550 693260 152640 693500
rect 152880 693260 152990 693500
rect 153230 693260 153320 693500
rect 153560 693260 153650 693500
rect 153890 693260 153980 693500
rect 154220 693260 154330 693500
rect 154570 693260 154660 693500
rect 154900 693260 154990 693500
rect 155230 693260 155320 693500
rect 155560 693260 155670 693500
rect 155910 693260 155960 693500
rect 110760 693150 155960 693260
rect 110760 692910 110810 693150
rect 111050 692910 111140 693150
rect 111380 692910 111470 693150
rect 111710 692910 111800 693150
rect 112040 692910 112150 693150
rect 112390 692910 112480 693150
rect 112720 692910 112810 693150
rect 113050 692910 113140 693150
rect 113380 692910 113490 693150
rect 113730 692910 113820 693150
rect 114060 692910 114150 693150
rect 114390 692910 114480 693150
rect 114720 692910 114830 693150
rect 115070 692910 115160 693150
rect 115400 692910 115490 693150
rect 115730 692910 115820 693150
rect 116060 692910 116170 693150
rect 116410 692910 116500 693150
rect 116740 692910 116830 693150
rect 117070 692910 117160 693150
rect 117400 692910 117510 693150
rect 117750 692910 117840 693150
rect 118080 692910 118170 693150
rect 118410 692910 118500 693150
rect 118740 692910 118850 693150
rect 119090 692910 119180 693150
rect 119420 692910 119510 693150
rect 119750 692910 119840 693150
rect 120080 692910 120190 693150
rect 120430 692910 120520 693150
rect 120760 692910 120850 693150
rect 121090 692910 121180 693150
rect 121420 692910 121530 693150
rect 121770 692910 122190 693150
rect 122430 692910 122520 693150
rect 122760 692910 122850 693150
rect 123090 692910 123180 693150
rect 123420 692910 123530 693150
rect 123770 692910 123860 693150
rect 124100 692910 124190 693150
rect 124430 692910 124520 693150
rect 124760 692910 124870 693150
rect 125110 692910 125200 693150
rect 125440 692910 125530 693150
rect 125770 692910 125860 693150
rect 126100 692910 126210 693150
rect 126450 692910 126540 693150
rect 126780 692910 126870 693150
rect 127110 692910 127200 693150
rect 127440 692910 127550 693150
rect 127790 692910 127880 693150
rect 128120 692910 128210 693150
rect 128450 692910 128540 693150
rect 128780 692910 128890 693150
rect 129130 692910 129220 693150
rect 129460 692910 129550 693150
rect 129790 692910 129880 693150
rect 130120 692910 130230 693150
rect 130470 692910 130560 693150
rect 130800 692910 130890 693150
rect 131130 692910 131220 693150
rect 131460 692910 131570 693150
rect 131810 692910 131900 693150
rect 132140 692910 132230 693150
rect 132470 692910 132560 693150
rect 132800 692910 132910 693150
rect 133150 692910 133570 693150
rect 133810 692910 133900 693150
rect 134140 692910 134230 693150
rect 134470 692910 134560 693150
rect 134800 692910 134910 693150
rect 135150 692910 135240 693150
rect 135480 692910 135570 693150
rect 135810 692910 135900 693150
rect 136140 692910 136250 693150
rect 136490 692910 136580 693150
rect 136820 692910 136910 693150
rect 137150 692910 137240 693150
rect 137480 692910 137590 693150
rect 137830 692910 137920 693150
rect 138160 692910 138250 693150
rect 138490 692910 138580 693150
rect 138820 692910 138930 693150
rect 139170 692910 139260 693150
rect 139500 692910 139590 693150
rect 139830 692910 139920 693150
rect 140160 692910 140270 693150
rect 140510 692910 140600 693150
rect 140840 692910 140930 693150
rect 141170 692910 141260 693150
rect 141500 692910 141610 693150
rect 141850 692910 141940 693150
rect 142180 692910 142270 693150
rect 142510 692910 142600 693150
rect 142840 692910 142950 693150
rect 143190 692910 143280 693150
rect 143520 692910 143610 693150
rect 143850 692910 143940 693150
rect 144180 692910 144290 693150
rect 144530 692910 144950 693150
rect 145190 692910 145280 693150
rect 145520 692910 145610 693150
rect 145850 692910 145940 693150
rect 146180 692910 146290 693150
rect 146530 692910 146620 693150
rect 146860 692910 146950 693150
rect 147190 692910 147280 693150
rect 147520 692910 147630 693150
rect 147870 692910 147960 693150
rect 148200 692910 148290 693150
rect 148530 692910 148620 693150
rect 148860 692910 148970 693150
rect 149210 692910 149300 693150
rect 149540 692910 149630 693150
rect 149870 692910 149960 693150
rect 150200 692910 150310 693150
rect 150550 692910 150640 693150
rect 150880 692910 150970 693150
rect 151210 692910 151300 693150
rect 151540 692910 151650 693150
rect 151890 692910 151980 693150
rect 152220 692910 152310 693150
rect 152550 692910 152640 693150
rect 152880 692910 152990 693150
rect 153230 692910 153320 693150
rect 153560 692910 153650 693150
rect 153890 692910 153980 693150
rect 154220 692910 154330 693150
rect 154570 692910 154660 693150
rect 154900 692910 154990 693150
rect 155230 692910 155320 693150
rect 155560 692910 155670 693150
rect 155910 692910 155960 693150
rect 110760 692820 155960 692910
rect 110760 692580 110810 692820
rect 111050 692580 111140 692820
rect 111380 692580 111470 692820
rect 111710 692580 111800 692820
rect 112040 692580 112150 692820
rect 112390 692580 112480 692820
rect 112720 692580 112810 692820
rect 113050 692580 113140 692820
rect 113380 692580 113490 692820
rect 113730 692580 113820 692820
rect 114060 692580 114150 692820
rect 114390 692580 114480 692820
rect 114720 692580 114830 692820
rect 115070 692580 115160 692820
rect 115400 692580 115490 692820
rect 115730 692580 115820 692820
rect 116060 692580 116170 692820
rect 116410 692580 116500 692820
rect 116740 692580 116830 692820
rect 117070 692580 117160 692820
rect 117400 692580 117510 692820
rect 117750 692580 117840 692820
rect 118080 692580 118170 692820
rect 118410 692580 118500 692820
rect 118740 692580 118850 692820
rect 119090 692580 119180 692820
rect 119420 692580 119510 692820
rect 119750 692580 119840 692820
rect 120080 692580 120190 692820
rect 120430 692580 120520 692820
rect 120760 692580 120850 692820
rect 121090 692580 121180 692820
rect 121420 692580 121530 692820
rect 121770 692580 122190 692820
rect 122430 692580 122520 692820
rect 122760 692580 122850 692820
rect 123090 692580 123180 692820
rect 123420 692580 123530 692820
rect 123770 692580 123860 692820
rect 124100 692580 124190 692820
rect 124430 692580 124520 692820
rect 124760 692580 124870 692820
rect 125110 692580 125200 692820
rect 125440 692580 125530 692820
rect 125770 692580 125860 692820
rect 126100 692580 126210 692820
rect 126450 692580 126540 692820
rect 126780 692580 126870 692820
rect 127110 692580 127200 692820
rect 127440 692580 127550 692820
rect 127790 692580 127880 692820
rect 128120 692580 128210 692820
rect 128450 692580 128540 692820
rect 128780 692580 128890 692820
rect 129130 692580 129220 692820
rect 129460 692580 129550 692820
rect 129790 692580 129880 692820
rect 130120 692580 130230 692820
rect 130470 692580 130560 692820
rect 130800 692580 130890 692820
rect 131130 692580 131220 692820
rect 131460 692580 131570 692820
rect 131810 692580 131900 692820
rect 132140 692580 132230 692820
rect 132470 692580 132560 692820
rect 132800 692580 132910 692820
rect 133150 692580 133570 692820
rect 133810 692580 133900 692820
rect 134140 692580 134230 692820
rect 134470 692580 134560 692820
rect 134800 692580 134910 692820
rect 135150 692580 135240 692820
rect 135480 692580 135570 692820
rect 135810 692580 135900 692820
rect 136140 692580 136250 692820
rect 136490 692580 136580 692820
rect 136820 692580 136910 692820
rect 137150 692580 137240 692820
rect 137480 692580 137590 692820
rect 137830 692580 137920 692820
rect 138160 692580 138250 692820
rect 138490 692580 138580 692820
rect 138820 692580 138930 692820
rect 139170 692580 139260 692820
rect 139500 692580 139590 692820
rect 139830 692580 139920 692820
rect 140160 692580 140270 692820
rect 140510 692580 140600 692820
rect 140840 692580 140930 692820
rect 141170 692580 141260 692820
rect 141500 692580 141610 692820
rect 141850 692580 141940 692820
rect 142180 692580 142270 692820
rect 142510 692580 142600 692820
rect 142840 692580 142950 692820
rect 143190 692580 143280 692820
rect 143520 692580 143610 692820
rect 143850 692580 143940 692820
rect 144180 692580 144290 692820
rect 144530 692580 144950 692820
rect 145190 692580 145280 692820
rect 145520 692580 145610 692820
rect 145850 692580 145940 692820
rect 146180 692580 146290 692820
rect 146530 692580 146620 692820
rect 146860 692580 146950 692820
rect 147190 692580 147280 692820
rect 147520 692580 147630 692820
rect 147870 692580 147960 692820
rect 148200 692580 148290 692820
rect 148530 692580 148620 692820
rect 148860 692580 148970 692820
rect 149210 692580 149300 692820
rect 149540 692580 149630 692820
rect 149870 692580 149960 692820
rect 150200 692580 150310 692820
rect 150550 692580 150640 692820
rect 150880 692580 150970 692820
rect 151210 692580 151300 692820
rect 151540 692580 151650 692820
rect 151890 692580 151980 692820
rect 152220 692580 152310 692820
rect 152550 692580 152640 692820
rect 152880 692580 152990 692820
rect 153230 692580 153320 692820
rect 153560 692580 153650 692820
rect 153890 692580 153980 692820
rect 154220 692580 154330 692820
rect 154570 692580 154660 692820
rect 154900 692580 154990 692820
rect 155230 692580 155320 692820
rect 155560 692580 155670 692820
rect 155910 692580 155960 692820
rect 110760 692490 155960 692580
rect 110760 692250 110810 692490
rect 111050 692250 111140 692490
rect 111380 692250 111470 692490
rect 111710 692250 111800 692490
rect 112040 692250 112150 692490
rect 112390 692250 112480 692490
rect 112720 692250 112810 692490
rect 113050 692250 113140 692490
rect 113380 692250 113490 692490
rect 113730 692250 113820 692490
rect 114060 692250 114150 692490
rect 114390 692250 114480 692490
rect 114720 692250 114830 692490
rect 115070 692250 115160 692490
rect 115400 692250 115490 692490
rect 115730 692250 115820 692490
rect 116060 692250 116170 692490
rect 116410 692250 116500 692490
rect 116740 692250 116830 692490
rect 117070 692250 117160 692490
rect 117400 692250 117510 692490
rect 117750 692250 117840 692490
rect 118080 692250 118170 692490
rect 118410 692250 118500 692490
rect 118740 692250 118850 692490
rect 119090 692250 119180 692490
rect 119420 692250 119510 692490
rect 119750 692250 119840 692490
rect 120080 692250 120190 692490
rect 120430 692250 120520 692490
rect 120760 692250 120850 692490
rect 121090 692250 121180 692490
rect 121420 692250 121530 692490
rect 121770 692250 122190 692490
rect 122430 692250 122520 692490
rect 122760 692250 122850 692490
rect 123090 692250 123180 692490
rect 123420 692250 123530 692490
rect 123770 692250 123860 692490
rect 124100 692250 124190 692490
rect 124430 692250 124520 692490
rect 124760 692250 124870 692490
rect 125110 692250 125200 692490
rect 125440 692250 125530 692490
rect 125770 692250 125860 692490
rect 126100 692250 126210 692490
rect 126450 692250 126540 692490
rect 126780 692250 126870 692490
rect 127110 692250 127200 692490
rect 127440 692250 127550 692490
rect 127790 692250 127880 692490
rect 128120 692250 128210 692490
rect 128450 692250 128540 692490
rect 128780 692250 128890 692490
rect 129130 692250 129220 692490
rect 129460 692250 129550 692490
rect 129790 692250 129880 692490
rect 130120 692250 130230 692490
rect 130470 692250 130560 692490
rect 130800 692250 130890 692490
rect 131130 692250 131220 692490
rect 131460 692250 131570 692490
rect 131810 692250 131900 692490
rect 132140 692250 132230 692490
rect 132470 692250 132560 692490
rect 132800 692250 132910 692490
rect 133150 692250 133570 692490
rect 133810 692250 133900 692490
rect 134140 692250 134230 692490
rect 134470 692250 134560 692490
rect 134800 692250 134910 692490
rect 135150 692250 135240 692490
rect 135480 692250 135570 692490
rect 135810 692250 135900 692490
rect 136140 692250 136250 692490
rect 136490 692250 136580 692490
rect 136820 692250 136910 692490
rect 137150 692250 137240 692490
rect 137480 692250 137590 692490
rect 137830 692250 137920 692490
rect 138160 692250 138250 692490
rect 138490 692250 138580 692490
rect 138820 692250 138930 692490
rect 139170 692250 139260 692490
rect 139500 692250 139590 692490
rect 139830 692250 139920 692490
rect 140160 692250 140270 692490
rect 140510 692250 140600 692490
rect 140840 692250 140930 692490
rect 141170 692250 141260 692490
rect 141500 692250 141610 692490
rect 141850 692250 141940 692490
rect 142180 692250 142270 692490
rect 142510 692250 142600 692490
rect 142840 692250 142950 692490
rect 143190 692250 143280 692490
rect 143520 692250 143610 692490
rect 143850 692250 143940 692490
rect 144180 692250 144290 692490
rect 144530 692250 144950 692490
rect 145190 692250 145280 692490
rect 145520 692250 145610 692490
rect 145850 692250 145940 692490
rect 146180 692250 146290 692490
rect 146530 692250 146620 692490
rect 146860 692250 146950 692490
rect 147190 692250 147280 692490
rect 147520 692250 147630 692490
rect 147870 692250 147960 692490
rect 148200 692250 148290 692490
rect 148530 692250 148620 692490
rect 148860 692250 148970 692490
rect 149210 692250 149300 692490
rect 149540 692250 149630 692490
rect 149870 692250 149960 692490
rect 150200 692250 150310 692490
rect 150550 692250 150640 692490
rect 150880 692250 150970 692490
rect 151210 692250 151300 692490
rect 151540 692250 151650 692490
rect 151890 692250 151980 692490
rect 152220 692250 152310 692490
rect 152550 692250 152640 692490
rect 152880 692250 152990 692490
rect 153230 692250 153320 692490
rect 153560 692250 153650 692490
rect 153890 692250 153980 692490
rect 154220 692250 154330 692490
rect 154570 692250 154660 692490
rect 154900 692250 154990 692490
rect 155230 692250 155320 692490
rect 155560 692250 155670 692490
rect 155910 692250 155960 692490
rect 110760 692160 155960 692250
rect 110760 691920 110810 692160
rect 111050 691920 111140 692160
rect 111380 691920 111470 692160
rect 111710 691920 111800 692160
rect 112040 691920 112150 692160
rect 112390 691920 112480 692160
rect 112720 691920 112810 692160
rect 113050 691920 113140 692160
rect 113380 691920 113490 692160
rect 113730 691920 113820 692160
rect 114060 691920 114150 692160
rect 114390 691920 114480 692160
rect 114720 691920 114830 692160
rect 115070 691920 115160 692160
rect 115400 691920 115490 692160
rect 115730 691920 115820 692160
rect 116060 691920 116170 692160
rect 116410 691920 116500 692160
rect 116740 691920 116830 692160
rect 117070 691920 117160 692160
rect 117400 691920 117510 692160
rect 117750 691920 117840 692160
rect 118080 691920 118170 692160
rect 118410 691920 118500 692160
rect 118740 691920 118850 692160
rect 119090 691920 119180 692160
rect 119420 691920 119510 692160
rect 119750 691920 119840 692160
rect 120080 691920 120190 692160
rect 120430 691920 120520 692160
rect 120760 691920 120850 692160
rect 121090 691920 121180 692160
rect 121420 691920 121530 692160
rect 121770 691920 122190 692160
rect 122430 691920 122520 692160
rect 122760 691920 122850 692160
rect 123090 691920 123180 692160
rect 123420 691920 123530 692160
rect 123770 691920 123860 692160
rect 124100 691920 124190 692160
rect 124430 691920 124520 692160
rect 124760 691920 124870 692160
rect 125110 691920 125200 692160
rect 125440 691920 125530 692160
rect 125770 691920 125860 692160
rect 126100 691920 126210 692160
rect 126450 691920 126540 692160
rect 126780 691920 126870 692160
rect 127110 691920 127200 692160
rect 127440 691920 127550 692160
rect 127790 691920 127880 692160
rect 128120 691920 128210 692160
rect 128450 691920 128540 692160
rect 128780 691920 128890 692160
rect 129130 691920 129220 692160
rect 129460 691920 129550 692160
rect 129790 691920 129880 692160
rect 130120 691920 130230 692160
rect 130470 691920 130560 692160
rect 130800 691920 130890 692160
rect 131130 691920 131220 692160
rect 131460 691920 131570 692160
rect 131810 691920 131900 692160
rect 132140 691920 132230 692160
rect 132470 691920 132560 692160
rect 132800 691920 132910 692160
rect 133150 691920 133570 692160
rect 133810 691920 133900 692160
rect 134140 691920 134230 692160
rect 134470 691920 134560 692160
rect 134800 691920 134910 692160
rect 135150 691920 135240 692160
rect 135480 691920 135570 692160
rect 135810 691920 135900 692160
rect 136140 691920 136250 692160
rect 136490 691920 136580 692160
rect 136820 691920 136910 692160
rect 137150 691920 137240 692160
rect 137480 691920 137590 692160
rect 137830 691920 137920 692160
rect 138160 691920 138250 692160
rect 138490 691920 138580 692160
rect 138820 691920 138930 692160
rect 139170 691920 139260 692160
rect 139500 691920 139590 692160
rect 139830 691920 139920 692160
rect 140160 691920 140270 692160
rect 140510 691920 140600 692160
rect 140840 691920 140930 692160
rect 141170 691920 141260 692160
rect 141500 691920 141610 692160
rect 141850 691920 141940 692160
rect 142180 691920 142270 692160
rect 142510 691920 142600 692160
rect 142840 691920 142950 692160
rect 143190 691920 143280 692160
rect 143520 691920 143610 692160
rect 143850 691920 143940 692160
rect 144180 691920 144290 692160
rect 144530 691920 144950 692160
rect 145190 691920 145280 692160
rect 145520 691920 145610 692160
rect 145850 691920 145940 692160
rect 146180 691920 146290 692160
rect 146530 691920 146620 692160
rect 146860 691920 146950 692160
rect 147190 691920 147280 692160
rect 147520 691920 147630 692160
rect 147870 691920 147960 692160
rect 148200 691920 148290 692160
rect 148530 691920 148620 692160
rect 148860 691920 148970 692160
rect 149210 691920 149300 692160
rect 149540 691920 149630 692160
rect 149870 691920 149960 692160
rect 150200 691920 150310 692160
rect 150550 691920 150640 692160
rect 150880 691920 150970 692160
rect 151210 691920 151300 692160
rect 151540 691920 151650 692160
rect 151890 691920 151980 692160
rect 152220 691920 152310 692160
rect 152550 691920 152640 692160
rect 152880 691920 152990 692160
rect 153230 691920 153320 692160
rect 153560 691920 153650 692160
rect 153890 691920 153980 692160
rect 154220 691920 154330 692160
rect 154570 691920 154660 692160
rect 154900 691920 154990 692160
rect 155230 691920 155320 692160
rect 155560 691920 155670 692160
rect 155910 691920 155960 692160
rect 110760 691810 155960 691920
rect 110760 691570 110810 691810
rect 111050 691570 111140 691810
rect 111380 691570 111470 691810
rect 111710 691570 111800 691810
rect 112040 691570 112150 691810
rect 112390 691570 112480 691810
rect 112720 691570 112810 691810
rect 113050 691570 113140 691810
rect 113380 691570 113490 691810
rect 113730 691570 113820 691810
rect 114060 691570 114150 691810
rect 114390 691570 114480 691810
rect 114720 691570 114830 691810
rect 115070 691570 115160 691810
rect 115400 691570 115490 691810
rect 115730 691570 115820 691810
rect 116060 691570 116170 691810
rect 116410 691570 116500 691810
rect 116740 691570 116830 691810
rect 117070 691570 117160 691810
rect 117400 691570 117510 691810
rect 117750 691570 117840 691810
rect 118080 691570 118170 691810
rect 118410 691570 118500 691810
rect 118740 691570 118850 691810
rect 119090 691570 119180 691810
rect 119420 691570 119510 691810
rect 119750 691570 119840 691810
rect 120080 691570 120190 691810
rect 120430 691570 120520 691810
rect 120760 691570 120850 691810
rect 121090 691570 121180 691810
rect 121420 691570 121530 691810
rect 121770 691570 122190 691810
rect 122430 691570 122520 691810
rect 122760 691570 122850 691810
rect 123090 691570 123180 691810
rect 123420 691570 123530 691810
rect 123770 691570 123860 691810
rect 124100 691570 124190 691810
rect 124430 691570 124520 691810
rect 124760 691570 124870 691810
rect 125110 691570 125200 691810
rect 125440 691570 125530 691810
rect 125770 691570 125860 691810
rect 126100 691570 126210 691810
rect 126450 691570 126540 691810
rect 126780 691570 126870 691810
rect 127110 691570 127200 691810
rect 127440 691570 127550 691810
rect 127790 691570 127880 691810
rect 128120 691570 128210 691810
rect 128450 691570 128540 691810
rect 128780 691570 128890 691810
rect 129130 691570 129220 691810
rect 129460 691570 129550 691810
rect 129790 691570 129880 691810
rect 130120 691570 130230 691810
rect 130470 691570 130560 691810
rect 130800 691570 130890 691810
rect 131130 691570 131220 691810
rect 131460 691570 131570 691810
rect 131810 691570 131900 691810
rect 132140 691570 132230 691810
rect 132470 691570 132560 691810
rect 132800 691570 132910 691810
rect 133150 691570 133570 691810
rect 133810 691570 133900 691810
rect 134140 691570 134230 691810
rect 134470 691570 134560 691810
rect 134800 691570 134910 691810
rect 135150 691570 135240 691810
rect 135480 691570 135570 691810
rect 135810 691570 135900 691810
rect 136140 691570 136250 691810
rect 136490 691570 136580 691810
rect 136820 691570 136910 691810
rect 137150 691570 137240 691810
rect 137480 691570 137590 691810
rect 137830 691570 137920 691810
rect 138160 691570 138250 691810
rect 138490 691570 138580 691810
rect 138820 691570 138930 691810
rect 139170 691570 139260 691810
rect 139500 691570 139590 691810
rect 139830 691570 139920 691810
rect 140160 691570 140270 691810
rect 140510 691570 140600 691810
rect 140840 691570 140930 691810
rect 141170 691570 141260 691810
rect 141500 691570 141610 691810
rect 141850 691570 141940 691810
rect 142180 691570 142270 691810
rect 142510 691570 142600 691810
rect 142840 691570 142950 691810
rect 143190 691570 143280 691810
rect 143520 691570 143610 691810
rect 143850 691570 143940 691810
rect 144180 691570 144290 691810
rect 144530 691570 144950 691810
rect 145190 691570 145280 691810
rect 145520 691570 145610 691810
rect 145850 691570 145940 691810
rect 146180 691570 146290 691810
rect 146530 691570 146620 691810
rect 146860 691570 146950 691810
rect 147190 691570 147280 691810
rect 147520 691570 147630 691810
rect 147870 691570 147960 691810
rect 148200 691570 148290 691810
rect 148530 691570 148620 691810
rect 148860 691570 148970 691810
rect 149210 691570 149300 691810
rect 149540 691570 149630 691810
rect 149870 691570 149960 691810
rect 150200 691570 150310 691810
rect 150550 691570 150640 691810
rect 150880 691570 150970 691810
rect 151210 691570 151300 691810
rect 151540 691570 151650 691810
rect 151890 691570 151980 691810
rect 152220 691570 152310 691810
rect 152550 691570 152640 691810
rect 152880 691570 152990 691810
rect 153230 691570 153320 691810
rect 153560 691570 153650 691810
rect 153890 691570 153980 691810
rect 154220 691570 154330 691810
rect 154570 691570 154660 691810
rect 154900 691570 154990 691810
rect 155230 691570 155320 691810
rect 155560 691570 155670 691810
rect 155910 691570 155960 691810
rect 110760 691480 155960 691570
rect 110760 691240 110810 691480
rect 111050 691240 111140 691480
rect 111380 691240 111470 691480
rect 111710 691240 111800 691480
rect 112040 691240 112150 691480
rect 112390 691240 112480 691480
rect 112720 691240 112810 691480
rect 113050 691240 113140 691480
rect 113380 691240 113490 691480
rect 113730 691240 113820 691480
rect 114060 691240 114150 691480
rect 114390 691240 114480 691480
rect 114720 691240 114830 691480
rect 115070 691240 115160 691480
rect 115400 691240 115490 691480
rect 115730 691240 115820 691480
rect 116060 691240 116170 691480
rect 116410 691240 116500 691480
rect 116740 691240 116830 691480
rect 117070 691240 117160 691480
rect 117400 691240 117510 691480
rect 117750 691240 117840 691480
rect 118080 691240 118170 691480
rect 118410 691240 118500 691480
rect 118740 691240 118850 691480
rect 119090 691240 119180 691480
rect 119420 691240 119510 691480
rect 119750 691240 119840 691480
rect 120080 691240 120190 691480
rect 120430 691240 120520 691480
rect 120760 691240 120850 691480
rect 121090 691240 121180 691480
rect 121420 691240 121530 691480
rect 121770 691240 122190 691480
rect 122430 691240 122520 691480
rect 122760 691240 122850 691480
rect 123090 691240 123180 691480
rect 123420 691240 123530 691480
rect 123770 691240 123860 691480
rect 124100 691240 124190 691480
rect 124430 691240 124520 691480
rect 124760 691240 124870 691480
rect 125110 691240 125200 691480
rect 125440 691240 125530 691480
rect 125770 691240 125860 691480
rect 126100 691240 126210 691480
rect 126450 691240 126540 691480
rect 126780 691240 126870 691480
rect 127110 691240 127200 691480
rect 127440 691240 127550 691480
rect 127790 691240 127880 691480
rect 128120 691240 128210 691480
rect 128450 691240 128540 691480
rect 128780 691240 128890 691480
rect 129130 691240 129220 691480
rect 129460 691240 129550 691480
rect 129790 691240 129880 691480
rect 130120 691240 130230 691480
rect 130470 691240 130560 691480
rect 130800 691240 130890 691480
rect 131130 691240 131220 691480
rect 131460 691240 131570 691480
rect 131810 691240 131900 691480
rect 132140 691240 132230 691480
rect 132470 691240 132560 691480
rect 132800 691240 132910 691480
rect 133150 691240 133570 691480
rect 133810 691240 133900 691480
rect 134140 691240 134230 691480
rect 134470 691240 134560 691480
rect 134800 691240 134910 691480
rect 135150 691240 135240 691480
rect 135480 691240 135570 691480
rect 135810 691240 135900 691480
rect 136140 691240 136250 691480
rect 136490 691240 136580 691480
rect 136820 691240 136910 691480
rect 137150 691240 137240 691480
rect 137480 691240 137590 691480
rect 137830 691240 137920 691480
rect 138160 691240 138250 691480
rect 138490 691240 138580 691480
rect 138820 691240 138930 691480
rect 139170 691240 139260 691480
rect 139500 691240 139590 691480
rect 139830 691240 139920 691480
rect 140160 691240 140270 691480
rect 140510 691240 140600 691480
rect 140840 691240 140930 691480
rect 141170 691240 141260 691480
rect 141500 691240 141610 691480
rect 141850 691240 141940 691480
rect 142180 691240 142270 691480
rect 142510 691240 142600 691480
rect 142840 691240 142950 691480
rect 143190 691240 143280 691480
rect 143520 691240 143610 691480
rect 143850 691240 143940 691480
rect 144180 691240 144290 691480
rect 144530 691240 144950 691480
rect 145190 691240 145280 691480
rect 145520 691240 145610 691480
rect 145850 691240 145940 691480
rect 146180 691240 146290 691480
rect 146530 691240 146620 691480
rect 146860 691240 146950 691480
rect 147190 691240 147280 691480
rect 147520 691240 147630 691480
rect 147870 691240 147960 691480
rect 148200 691240 148290 691480
rect 148530 691240 148620 691480
rect 148860 691240 148970 691480
rect 149210 691240 149300 691480
rect 149540 691240 149630 691480
rect 149870 691240 149960 691480
rect 150200 691240 150310 691480
rect 150550 691240 150640 691480
rect 150880 691240 150970 691480
rect 151210 691240 151300 691480
rect 151540 691240 151650 691480
rect 151890 691240 151980 691480
rect 152220 691240 152310 691480
rect 152550 691240 152640 691480
rect 152880 691240 152990 691480
rect 153230 691240 153320 691480
rect 153560 691240 153650 691480
rect 153890 691240 153980 691480
rect 154220 691240 154330 691480
rect 154570 691240 154660 691480
rect 154900 691240 154990 691480
rect 155230 691240 155320 691480
rect 155560 691240 155670 691480
rect 155910 691240 155960 691480
rect 110760 691150 155960 691240
rect 110760 691028 110810 691150
rect 103643 690910 110810 691028
rect 111050 690910 111140 691150
rect 111380 690910 111470 691150
rect 111710 690910 111800 691150
rect 112040 690910 112150 691150
rect 112390 690910 112480 691150
rect 112720 690910 112810 691150
rect 113050 690910 113140 691150
rect 113380 690910 113490 691150
rect 113730 690910 113820 691150
rect 114060 690910 114150 691150
rect 114390 690910 114480 691150
rect 114720 690910 114830 691150
rect 115070 690910 115160 691150
rect 115400 690910 115490 691150
rect 115730 690910 115820 691150
rect 116060 690910 116170 691150
rect 116410 690910 116500 691150
rect 116740 690910 116830 691150
rect 117070 690910 117160 691150
rect 117400 690910 117510 691150
rect 117750 690910 117840 691150
rect 118080 690910 118170 691150
rect 118410 690910 118500 691150
rect 118740 690910 118850 691150
rect 119090 690910 119180 691150
rect 119420 690910 119510 691150
rect 119750 690910 119840 691150
rect 120080 690910 120190 691150
rect 120430 690910 120520 691150
rect 120760 690910 120850 691150
rect 121090 690910 121180 691150
rect 121420 690910 121530 691150
rect 121770 690910 122190 691150
rect 122430 690910 122520 691150
rect 122760 690910 122850 691150
rect 123090 690910 123180 691150
rect 123420 690910 123530 691150
rect 123770 690910 123860 691150
rect 124100 690910 124190 691150
rect 124430 690910 124520 691150
rect 124760 690910 124870 691150
rect 125110 690910 125200 691150
rect 125440 690910 125530 691150
rect 125770 690910 125860 691150
rect 126100 690910 126210 691150
rect 126450 690910 126540 691150
rect 126780 690910 126870 691150
rect 127110 690910 127200 691150
rect 127440 690910 127550 691150
rect 127790 690910 127880 691150
rect 128120 690910 128210 691150
rect 128450 690910 128540 691150
rect 128780 690910 128890 691150
rect 129130 690910 129220 691150
rect 129460 690910 129550 691150
rect 129790 690910 129880 691150
rect 130120 690910 130230 691150
rect 130470 690910 130560 691150
rect 130800 690910 130890 691150
rect 131130 690910 131220 691150
rect 131460 690910 131570 691150
rect 131810 690910 131900 691150
rect 132140 690910 132230 691150
rect 132470 690910 132560 691150
rect 132800 690910 132910 691150
rect 133150 690910 133570 691150
rect 133810 690910 133900 691150
rect 134140 690910 134230 691150
rect 134470 690910 134560 691150
rect 134800 690910 134910 691150
rect 135150 690910 135240 691150
rect 135480 690910 135570 691150
rect 135810 690910 135900 691150
rect 136140 690910 136250 691150
rect 136490 690910 136580 691150
rect 136820 690910 136910 691150
rect 137150 690910 137240 691150
rect 137480 690910 137590 691150
rect 137830 690910 137920 691150
rect 138160 690910 138250 691150
rect 138490 690910 138580 691150
rect 138820 690910 138930 691150
rect 139170 690910 139260 691150
rect 139500 690910 139590 691150
rect 139830 690910 139920 691150
rect 140160 690910 140270 691150
rect 140510 690910 140600 691150
rect 140840 690910 140930 691150
rect 141170 690910 141260 691150
rect 141500 690910 141610 691150
rect 141850 690910 141940 691150
rect 142180 690910 142270 691150
rect 142510 690910 142600 691150
rect 142840 690910 142950 691150
rect 143190 690910 143280 691150
rect 143520 690910 143610 691150
rect 143850 690910 143940 691150
rect 144180 690910 144290 691150
rect 144530 690910 144950 691150
rect 145190 690910 145280 691150
rect 145520 690910 145610 691150
rect 145850 690910 145940 691150
rect 146180 690910 146290 691150
rect 146530 690910 146620 691150
rect 146860 690910 146950 691150
rect 147190 690910 147280 691150
rect 147520 690910 147630 691150
rect 147870 690910 147960 691150
rect 148200 690910 148290 691150
rect 148530 690910 148620 691150
rect 148860 690910 148970 691150
rect 149210 690910 149300 691150
rect 149540 690910 149630 691150
rect 149870 690910 149960 691150
rect 150200 690910 150310 691150
rect 150550 690910 150640 691150
rect 150880 690910 150970 691150
rect 151210 690910 151300 691150
rect 151540 690910 151650 691150
rect 151890 690910 151980 691150
rect 152220 690910 152310 691150
rect 152550 690910 152640 691150
rect 152880 690910 152990 691150
rect 153230 690910 153320 691150
rect 153560 690910 153650 691150
rect 153890 690910 153980 691150
rect 154220 690910 154330 691150
rect 154570 690910 154660 691150
rect 154900 690910 154990 691150
rect 155230 690910 155320 691150
rect 155560 690910 155670 691150
rect 155910 691028 155960 691150
rect 155910 690910 162436 691028
rect 103643 690820 162436 690910
rect 103643 690580 110810 690820
rect 111050 690580 111140 690820
rect 111380 690580 111470 690820
rect 111710 690580 111800 690820
rect 112040 690580 112150 690820
rect 112390 690580 112480 690820
rect 112720 690580 112810 690820
rect 113050 690580 113140 690820
rect 113380 690580 113490 690820
rect 113730 690580 113820 690820
rect 114060 690580 114150 690820
rect 114390 690580 114480 690820
rect 114720 690580 114830 690820
rect 115070 690580 115160 690820
rect 115400 690580 115490 690820
rect 115730 690580 115820 690820
rect 116060 690580 116170 690820
rect 116410 690580 116500 690820
rect 116740 690580 116830 690820
rect 117070 690580 117160 690820
rect 117400 690580 117510 690820
rect 117750 690580 117840 690820
rect 118080 690580 118170 690820
rect 118410 690580 118500 690820
rect 118740 690580 118850 690820
rect 119090 690580 119180 690820
rect 119420 690580 119510 690820
rect 119750 690580 119840 690820
rect 120080 690580 120190 690820
rect 120430 690580 120520 690820
rect 120760 690580 120850 690820
rect 121090 690580 121180 690820
rect 121420 690580 121530 690820
rect 121770 690580 122190 690820
rect 122430 690580 122520 690820
rect 122760 690580 122850 690820
rect 123090 690580 123180 690820
rect 123420 690580 123530 690820
rect 123770 690580 123860 690820
rect 124100 690580 124190 690820
rect 124430 690580 124520 690820
rect 124760 690580 124870 690820
rect 125110 690580 125200 690820
rect 125440 690580 125530 690820
rect 125770 690580 125860 690820
rect 126100 690580 126210 690820
rect 126450 690580 126540 690820
rect 126780 690580 126870 690820
rect 127110 690580 127200 690820
rect 127440 690580 127550 690820
rect 127790 690580 127880 690820
rect 128120 690580 128210 690820
rect 128450 690580 128540 690820
rect 128780 690580 128890 690820
rect 129130 690580 129220 690820
rect 129460 690580 129550 690820
rect 129790 690580 129880 690820
rect 130120 690580 130230 690820
rect 130470 690580 130560 690820
rect 130800 690580 130890 690820
rect 131130 690580 131220 690820
rect 131460 690580 131570 690820
rect 131810 690580 131900 690820
rect 132140 690580 132230 690820
rect 132470 690580 132560 690820
rect 132800 690580 132910 690820
rect 133150 690580 133570 690820
rect 133810 690580 133900 690820
rect 134140 690580 134230 690820
rect 134470 690580 134560 690820
rect 134800 690580 134910 690820
rect 135150 690580 135240 690820
rect 135480 690580 135570 690820
rect 135810 690580 135900 690820
rect 136140 690580 136250 690820
rect 136490 690580 136580 690820
rect 136820 690580 136910 690820
rect 137150 690580 137240 690820
rect 137480 690580 137590 690820
rect 137830 690580 137920 690820
rect 138160 690580 138250 690820
rect 138490 690580 138580 690820
rect 138820 690580 138930 690820
rect 139170 690580 139260 690820
rect 139500 690580 139590 690820
rect 139830 690580 139920 690820
rect 140160 690580 140270 690820
rect 140510 690580 140600 690820
rect 140840 690580 140930 690820
rect 141170 690580 141260 690820
rect 141500 690580 141610 690820
rect 141850 690580 141940 690820
rect 142180 690580 142270 690820
rect 142510 690580 142600 690820
rect 142840 690580 142950 690820
rect 143190 690580 143280 690820
rect 143520 690580 143610 690820
rect 143850 690580 143940 690820
rect 144180 690580 144290 690820
rect 144530 690580 144950 690820
rect 145190 690580 145280 690820
rect 145520 690580 145610 690820
rect 145850 690580 145940 690820
rect 146180 690580 146290 690820
rect 146530 690580 146620 690820
rect 146860 690580 146950 690820
rect 147190 690580 147280 690820
rect 147520 690580 147630 690820
rect 147870 690580 147960 690820
rect 148200 690580 148290 690820
rect 148530 690580 148620 690820
rect 148860 690580 148970 690820
rect 149210 690580 149300 690820
rect 149540 690580 149630 690820
rect 149870 690580 149960 690820
rect 150200 690580 150310 690820
rect 150550 690580 150640 690820
rect 150880 690580 150970 690820
rect 151210 690580 151300 690820
rect 151540 690580 151650 690820
rect 151890 690580 151980 690820
rect 152220 690580 152310 690820
rect 152550 690580 152640 690820
rect 152880 690580 152990 690820
rect 153230 690580 153320 690820
rect 153560 690580 153650 690820
rect 153890 690580 153980 690820
rect 154220 690580 154330 690820
rect 154570 690580 154660 690820
rect 154900 690580 154990 690820
rect 155230 690580 155320 690820
rect 155560 690580 155670 690820
rect 155910 690580 162436 690820
rect 103643 690470 162436 690580
rect 103643 690230 110810 690470
rect 111050 690230 111140 690470
rect 111380 690230 111470 690470
rect 111710 690230 111800 690470
rect 112040 690230 112150 690470
rect 112390 690230 112480 690470
rect 112720 690230 112810 690470
rect 113050 690230 113140 690470
rect 113380 690230 113490 690470
rect 113730 690230 113820 690470
rect 114060 690230 114150 690470
rect 114390 690230 114480 690470
rect 114720 690230 114830 690470
rect 115070 690230 115160 690470
rect 115400 690230 115490 690470
rect 115730 690230 115820 690470
rect 116060 690230 116170 690470
rect 116410 690230 116500 690470
rect 116740 690230 116830 690470
rect 117070 690230 117160 690470
rect 117400 690230 117510 690470
rect 117750 690230 117840 690470
rect 118080 690230 118170 690470
rect 118410 690230 118500 690470
rect 118740 690230 118850 690470
rect 119090 690230 119180 690470
rect 119420 690230 119510 690470
rect 119750 690230 119840 690470
rect 120080 690230 120190 690470
rect 120430 690230 120520 690470
rect 120760 690230 120850 690470
rect 121090 690230 121180 690470
rect 121420 690230 121530 690470
rect 121770 690230 122190 690470
rect 122430 690230 122520 690470
rect 122760 690230 122850 690470
rect 123090 690230 123180 690470
rect 123420 690230 123530 690470
rect 123770 690230 123860 690470
rect 124100 690230 124190 690470
rect 124430 690230 124520 690470
rect 124760 690230 124870 690470
rect 125110 690230 125200 690470
rect 125440 690230 125530 690470
rect 125770 690230 125860 690470
rect 126100 690230 126210 690470
rect 126450 690230 126540 690470
rect 126780 690230 126870 690470
rect 127110 690230 127200 690470
rect 127440 690230 127550 690470
rect 127790 690230 127880 690470
rect 128120 690230 128210 690470
rect 128450 690230 128540 690470
rect 128780 690230 128890 690470
rect 129130 690230 129220 690470
rect 129460 690230 129550 690470
rect 129790 690230 129880 690470
rect 130120 690230 130230 690470
rect 130470 690230 130560 690470
rect 130800 690230 130890 690470
rect 131130 690230 131220 690470
rect 131460 690230 131570 690470
rect 131810 690230 131900 690470
rect 132140 690230 132230 690470
rect 132470 690230 132560 690470
rect 132800 690230 132910 690470
rect 133150 690230 133570 690470
rect 133810 690230 133900 690470
rect 134140 690230 134230 690470
rect 134470 690230 134560 690470
rect 134800 690230 134910 690470
rect 135150 690230 135240 690470
rect 135480 690230 135570 690470
rect 135810 690230 135900 690470
rect 136140 690230 136250 690470
rect 136490 690230 136580 690470
rect 136820 690230 136910 690470
rect 137150 690230 137240 690470
rect 137480 690230 137590 690470
rect 137830 690230 137920 690470
rect 138160 690230 138250 690470
rect 138490 690230 138580 690470
rect 138820 690230 138930 690470
rect 139170 690230 139260 690470
rect 139500 690230 139590 690470
rect 139830 690230 139920 690470
rect 140160 690230 140270 690470
rect 140510 690230 140600 690470
rect 140840 690230 140930 690470
rect 141170 690230 141260 690470
rect 141500 690230 141610 690470
rect 141850 690230 141940 690470
rect 142180 690230 142270 690470
rect 142510 690230 142600 690470
rect 142840 690230 142950 690470
rect 143190 690230 143280 690470
rect 143520 690230 143610 690470
rect 143850 690230 143940 690470
rect 144180 690230 144290 690470
rect 144530 690230 144950 690470
rect 145190 690230 145280 690470
rect 145520 690230 145610 690470
rect 145850 690230 145940 690470
rect 146180 690230 146290 690470
rect 146530 690230 146620 690470
rect 146860 690230 146950 690470
rect 147190 690230 147280 690470
rect 147520 690230 147630 690470
rect 147870 690230 147960 690470
rect 148200 690230 148290 690470
rect 148530 690230 148620 690470
rect 148860 690230 148970 690470
rect 149210 690230 149300 690470
rect 149540 690230 149630 690470
rect 149870 690230 149960 690470
rect 150200 690230 150310 690470
rect 150550 690230 150640 690470
rect 150880 690230 150970 690470
rect 151210 690230 151300 690470
rect 151540 690230 151650 690470
rect 151890 690230 151980 690470
rect 152220 690230 152310 690470
rect 152550 690230 152640 690470
rect 152880 690230 152990 690470
rect 153230 690230 153320 690470
rect 153560 690230 153650 690470
rect 153890 690230 153980 690470
rect 154220 690230 154330 690470
rect 154570 690230 154660 690470
rect 154900 690230 154990 690470
rect 155230 690230 155320 690470
rect 155560 690230 155670 690470
rect 155910 690230 162436 690470
rect 103643 690140 162436 690230
rect 103643 689900 110810 690140
rect 111050 689900 111140 690140
rect 111380 689900 111470 690140
rect 111710 689900 111800 690140
rect 112040 689900 112150 690140
rect 112390 689900 112480 690140
rect 112720 689900 112810 690140
rect 113050 689900 113140 690140
rect 113380 689900 113490 690140
rect 113730 689900 113820 690140
rect 114060 689900 114150 690140
rect 114390 689900 114480 690140
rect 114720 689900 114830 690140
rect 115070 689900 115160 690140
rect 115400 689900 115490 690140
rect 115730 689900 115820 690140
rect 116060 689900 116170 690140
rect 116410 689900 116500 690140
rect 116740 689900 116830 690140
rect 117070 689900 117160 690140
rect 117400 689900 117510 690140
rect 117750 689900 117840 690140
rect 118080 689900 118170 690140
rect 118410 689900 118500 690140
rect 118740 689900 118850 690140
rect 119090 689900 119180 690140
rect 119420 689900 119510 690140
rect 119750 689900 119840 690140
rect 120080 689900 120190 690140
rect 120430 689900 120520 690140
rect 120760 689900 120850 690140
rect 121090 689900 121180 690140
rect 121420 689900 121530 690140
rect 121770 689900 122190 690140
rect 122430 689900 122520 690140
rect 122760 689900 122850 690140
rect 123090 689900 123180 690140
rect 123420 689900 123530 690140
rect 123770 689900 123860 690140
rect 124100 689900 124190 690140
rect 124430 689900 124520 690140
rect 124760 689900 124870 690140
rect 125110 689900 125200 690140
rect 125440 689900 125530 690140
rect 125770 689900 125860 690140
rect 126100 689900 126210 690140
rect 126450 689900 126540 690140
rect 126780 689900 126870 690140
rect 127110 689900 127200 690140
rect 127440 689900 127550 690140
rect 127790 689900 127880 690140
rect 128120 689900 128210 690140
rect 128450 689900 128540 690140
rect 128780 689900 128890 690140
rect 129130 689900 129220 690140
rect 129460 689900 129550 690140
rect 129790 689900 129880 690140
rect 130120 689900 130230 690140
rect 130470 689900 130560 690140
rect 130800 689900 130890 690140
rect 131130 689900 131220 690140
rect 131460 689900 131570 690140
rect 131810 689900 131900 690140
rect 132140 689900 132230 690140
rect 132470 689900 132560 690140
rect 132800 689900 132910 690140
rect 133150 689900 133570 690140
rect 133810 689900 133900 690140
rect 134140 689900 134230 690140
rect 134470 689900 134560 690140
rect 134800 689900 134910 690140
rect 135150 689900 135240 690140
rect 135480 689900 135570 690140
rect 135810 689900 135900 690140
rect 136140 689900 136250 690140
rect 136490 689900 136580 690140
rect 136820 689900 136910 690140
rect 137150 689900 137240 690140
rect 137480 689900 137590 690140
rect 137830 689900 137920 690140
rect 138160 689900 138250 690140
rect 138490 689900 138580 690140
rect 138820 689900 138930 690140
rect 139170 689900 139260 690140
rect 139500 689900 139590 690140
rect 139830 689900 139920 690140
rect 140160 689900 140270 690140
rect 140510 689900 140600 690140
rect 140840 689900 140930 690140
rect 141170 689900 141260 690140
rect 141500 689900 141610 690140
rect 141850 689900 141940 690140
rect 142180 689900 142270 690140
rect 142510 689900 142600 690140
rect 142840 689900 142950 690140
rect 143190 689900 143280 690140
rect 143520 689900 143610 690140
rect 143850 689900 143940 690140
rect 144180 689900 144290 690140
rect 144530 689900 144950 690140
rect 145190 689900 145280 690140
rect 145520 689900 145610 690140
rect 145850 689900 145940 690140
rect 146180 689900 146290 690140
rect 146530 689900 146620 690140
rect 146860 689900 146950 690140
rect 147190 689900 147280 690140
rect 147520 689900 147630 690140
rect 147870 689900 147960 690140
rect 148200 689900 148290 690140
rect 148530 689900 148620 690140
rect 148860 689900 148970 690140
rect 149210 689900 149300 690140
rect 149540 689900 149630 690140
rect 149870 689900 149960 690140
rect 150200 689900 150310 690140
rect 150550 689900 150640 690140
rect 150880 689900 150970 690140
rect 151210 689900 151300 690140
rect 151540 689900 151650 690140
rect 151890 689900 151980 690140
rect 152220 689900 152310 690140
rect 152550 689900 152640 690140
rect 152880 689900 152990 690140
rect 153230 689900 153320 690140
rect 153560 689900 153650 690140
rect 153890 689900 153980 690140
rect 154220 689900 154330 690140
rect 154570 689900 154660 690140
rect 154900 689900 154990 690140
rect 155230 689900 155320 690140
rect 155560 689900 155670 690140
rect 155910 689900 162436 690140
rect 103643 689810 162436 689900
rect 103643 689570 110810 689810
rect 111050 689570 111140 689810
rect 111380 689570 111470 689810
rect 111710 689570 111800 689810
rect 112040 689570 112150 689810
rect 112390 689570 112480 689810
rect 112720 689570 112810 689810
rect 113050 689570 113140 689810
rect 113380 689570 113490 689810
rect 113730 689570 113820 689810
rect 114060 689570 114150 689810
rect 114390 689570 114480 689810
rect 114720 689570 114830 689810
rect 115070 689570 115160 689810
rect 115400 689570 115490 689810
rect 115730 689570 115820 689810
rect 116060 689570 116170 689810
rect 116410 689570 116500 689810
rect 116740 689570 116830 689810
rect 117070 689570 117160 689810
rect 117400 689570 117510 689810
rect 117750 689570 117840 689810
rect 118080 689570 118170 689810
rect 118410 689570 118500 689810
rect 118740 689570 118850 689810
rect 119090 689570 119180 689810
rect 119420 689570 119510 689810
rect 119750 689570 119840 689810
rect 120080 689570 120190 689810
rect 120430 689570 120520 689810
rect 120760 689570 120850 689810
rect 121090 689570 121180 689810
rect 121420 689570 121530 689810
rect 121770 689570 122190 689810
rect 122430 689570 122520 689810
rect 122760 689570 122850 689810
rect 123090 689570 123180 689810
rect 123420 689570 123530 689810
rect 123770 689570 123860 689810
rect 124100 689570 124190 689810
rect 124430 689570 124520 689810
rect 124760 689570 124870 689810
rect 125110 689570 125200 689810
rect 125440 689570 125530 689810
rect 125770 689570 125860 689810
rect 126100 689570 126210 689810
rect 126450 689570 126540 689810
rect 126780 689570 126870 689810
rect 127110 689570 127200 689810
rect 127440 689570 127550 689810
rect 127790 689570 127880 689810
rect 128120 689570 128210 689810
rect 128450 689570 128540 689810
rect 128780 689570 128890 689810
rect 129130 689570 129220 689810
rect 129460 689570 129550 689810
rect 129790 689570 129880 689810
rect 130120 689570 130230 689810
rect 130470 689570 130560 689810
rect 130800 689570 130890 689810
rect 131130 689570 131220 689810
rect 131460 689570 131570 689810
rect 131810 689570 131900 689810
rect 132140 689570 132230 689810
rect 132470 689570 132560 689810
rect 132800 689570 132910 689810
rect 133150 689570 133570 689810
rect 133810 689570 133900 689810
rect 134140 689570 134230 689810
rect 134470 689570 134560 689810
rect 134800 689570 134910 689810
rect 135150 689570 135240 689810
rect 135480 689570 135570 689810
rect 135810 689570 135900 689810
rect 136140 689570 136250 689810
rect 136490 689570 136580 689810
rect 136820 689570 136910 689810
rect 137150 689570 137240 689810
rect 137480 689570 137590 689810
rect 137830 689570 137920 689810
rect 138160 689570 138250 689810
rect 138490 689570 138580 689810
rect 138820 689570 138930 689810
rect 139170 689570 139260 689810
rect 139500 689570 139590 689810
rect 139830 689570 139920 689810
rect 140160 689570 140270 689810
rect 140510 689570 140600 689810
rect 140840 689570 140930 689810
rect 141170 689570 141260 689810
rect 141500 689570 141610 689810
rect 141850 689570 141940 689810
rect 142180 689570 142270 689810
rect 142510 689570 142600 689810
rect 142840 689570 142950 689810
rect 143190 689570 143280 689810
rect 143520 689570 143610 689810
rect 143850 689570 143940 689810
rect 144180 689570 144290 689810
rect 144530 689570 144950 689810
rect 145190 689570 145280 689810
rect 145520 689570 145610 689810
rect 145850 689570 145940 689810
rect 146180 689570 146290 689810
rect 146530 689570 146620 689810
rect 146860 689570 146950 689810
rect 147190 689570 147280 689810
rect 147520 689570 147630 689810
rect 147870 689570 147960 689810
rect 148200 689570 148290 689810
rect 148530 689570 148620 689810
rect 148860 689570 148970 689810
rect 149210 689570 149300 689810
rect 149540 689570 149630 689810
rect 149870 689570 149960 689810
rect 150200 689570 150310 689810
rect 150550 689570 150640 689810
rect 150880 689570 150970 689810
rect 151210 689570 151300 689810
rect 151540 689570 151650 689810
rect 151890 689570 151980 689810
rect 152220 689570 152310 689810
rect 152550 689570 152640 689810
rect 152880 689570 152990 689810
rect 153230 689570 153320 689810
rect 153560 689570 153650 689810
rect 153890 689570 153980 689810
rect 154220 689570 154330 689810
rect 154570 689570 154660 689810
rect 154900 689570 154990 689810
rect 155230 689570 155320 689810
rect 155560 689570 155670 689810
rect 155910 689570 162436 689810
rect 103643 689480 162436 689570
rect 103643 689240 110810 689480
rect 111050 689240 111140 689480
rect 111380 689240 111470 689480
rect 111710 689240 111800 689480
rect 112040 689240 112150 689480
rect 112390 689240 112480 689480
rect 112720 689240 112810 689480
rect 113050 689240 113140 689480
rect 113380 689240 113490 689480
rect 113730 689240 113820 689480
rect 114060 689240 114150 689480
rect 114390 689240 114480 689480
rect 114720 689240 114830 689480
rect 115070 689240 115160 689480
rect 115400 689240 115490 689480
rect 115730 689240 115820 689480
rect 116060 689240 116170 689480
rect 116410 689240 116500 689480
rect 116740 689240 116830 689480
rect 117070 689240 117160 689480
rect 117400 689240 117510 689480
rect 117750 689240 117840 689480
rect 118080 689240 118170 689480
rect 118410 689240 118500 689480
rect 118740 689240 118850 689480
rect 119090 689240 119180 689480
rect 119420 689240 119510 689480
rect 119750 689240 119840 689480
rect 120080 689240 120190 689480
rect 120430 689240 120520 689480
rect 120760 689240 120850 689480
rect 121090 689240 121180 689480
rect 121420 689240 121530 689480
rect 121770 689240 122190 689480
rect 122430 689240 122520 689480
rect 122760 689240 122850 689480
rect 123090 689240 123180 689480
rect 123420 689240 123530 689480
rect 123770 689240 123860 689480
rect 124100 689240 124190 689480
rect 124430 689240 124520 689480
rect 124760 689240 124870 689480
rect 125110 689240 125200 689480
rect 125440 689240 125530 689480
rect 125770 689240 125860 689480
rect 126100 689240 126210 689480
rect 126450 689240 126540 689480
rect 126780 689240 126870 689480
rect 127110 689240 127200 689480
rect 127440 689240 127550 689480
rect 127790 689240 127880 689480
rect 128120 689240 128210 689480
rect 128450 689240 128540 689480
rect 128780 689240 128890 689480
rect 129130 689240 129220 689480
rect 129460 689240 129550 689480
rect 129790 689240 129880 689480
rect 130120 689240 130230 689480
rect 130470 689240 130560 689480
rect 130800 689240 130890 689480
rect 131130 689240 131220 689480
rect 131460 689240 131570 689480
rect 131810 689240 131900 689480
rect 132140 689240 132230 689480
rect 132470 689240 132560 689480
rect 132800 689240 132910 689480
rect 133150 689240 133570 689480
rect 133810 689240 133900 689480
rect 134140 689240 134230 689480
rect 134470 689240 134560 689480
rect 134800 689240 134910 689480
rect 135150 689240 135240 689480
rect 135480 689240 135570 689480
rect 135810 689240 135900 689480
rect 136140 689240 136250 689480
rect 136490 689240 136580 689480
rect 136820 689240 136910 689480
rect 137150 689240 137240 689480
rect 137480 689240 137590 689480
rect 137830 689240 137920 689480
rect 138160 689240 138250 689480
rect 138490 689240 138580 689480
rect 138820 689240 138930 689480
rect 139170 689240 139260 689480
rect 139500 689240 139590 689480
rect 139830 689240 139920 689480
rect 140160 689240 140270 689480
rect 140510 689240 140600 689480
rect 140840 689240 140930 689480
rect 141170 689240 141260 689480
rect 141500 689240 141610 689480
rect 141850 689240 141940 689480
rect 142180 689240 142270 689480
rect 142510 689240 142600 689480
rect 142840 689240 142950 689480
rect 143190 689240 143280 689480
rect 143520 689240 143610 689480
rect 143850 689240 143940 689480
rect 144180 689240 144290 689480
rect 144530 689240 144950 689480
rect 145190 689240 145280 689480
rect 145520 689240 145610 689480
rect 145850 689240 145940 689480
rect 146180 689240 146290 689480
rect 146530 689240 146620 689480
rect 146860 689240 146950 689480
rect 147190 689240 147280 689480
rect 147520 689240 147630 689480
rect 147870 689240 147960 689480
rect 148200 689240 148290 689480
rect 148530 689240 148620 689480
rect 148860 689240 148970 689480
rect 149210 689240 149300 689480
rect 149540 689240 149630 689480
rect 149870 689240 149960 689480
rect 150200 689240 150310 689480
rect 150550 689240 150640 689480
rect 150880 689240 150970 689480
rect 151210 689240 151300 689480
rect 151540 689240 151650 689480
rect 151890 689240 151980 689480
rect 152220 689240 152310 689480
rect 152550 689240 152640 689480
rect 152880 689240 152990 689480
rect 153230 689240 153320 689480
rect 153560 689240 153650 689480
rect 153890 689240 153980 689480
rect 154220 689240 154330 689480
rect 154570 689240 154660 689480
rect 154900 689240 154990 689480
rect 155230 689240 155320 689480
rect 155560 689240 155670 689480
rect 155910 689240 162436 689480
rect 103643 689130 162436 689240
rect 103643 688890 110810 689130
rect 111050 688890 111140 689130
rect 111380 688890 111470 689130
rect 111710 688890 111800 689130
rect 112040 688890 112150 689130
rect 112390 688890 112480 689130
rect 112720 688890 112810 689130
rect 113050 688890 113140 689130
rect 113380 688890 113490 689130
rect 113730 688890 113820 689130
rect 114060 688890 114150 689130
rect 114390 688890 114480 689130
rect 114720 688890 114830 689130
rect 115070 688890 115160 689130
rect 115400 688890 115490 689130
rect 115730 688890 115820 689130
rect 116060 688890 116170 689130
rect 116410 688890 116500 689130
rect 116740 688890 116830 689130
rect 117070 688890 117160 689130
rect 117400 688890 117510 689130
rect 117750 688890 117840 689130
rect 118080 688890 118170 689130
rect 118410 688890 118500 689130
rect 118740 688890 118850 689130
rect 119090 688890 119180 689130
rect 119420 688890 119510 689130
rect 119750 688890 119840 689130
rect 120080 688890 120190 689130
rect 120430 688890 120520 689130
rect 120760 688890 120850 689130
rect 121090 688890 121180 689130
rect 121420 688890 121530 689130
rect 121770 688890 122190 689130
rect 122430 688890 122520 689130
rect 122760 688890 122850 689130
rect 123090 688890 123180 689130
rect 123420 688890 123530 689130
rect 123770 688890 123860 689130
rect 124100 688890 124190 689130
rect 124430 688890 124520 689130
rect 124760 688890 124870 689130
rect 125110 688890 125200 689130
rect 125440 688890 125530 689130
rect 125770 688890 125860 689130
rect 126100 688890 126210 689130
rect 126450 688890 126540 689130
rect 126780 688890 126870 689130
rect 127110 688890 127200 689130
rect 127440 688890 127550 689130
rect 127790 688890 127880 689130
rect 128120 688890 128210 689130
rect 128450 688890 128540 689130
rect 128780 688890 128890 689130
rect 129130 688890 129220 689130
rect 129460 688890 129550 689130
rect 129790 688890 129880 689130
rect 130120 688890 130230 689130
rect 130470 688890 130560 689130
rect 130800 688890 130890 689130
rect 131130 688890 131220 689130
rect 131460 688890 131570 689130
rect 131810 688890 131900 689130
rect 132140 688890 132230 689130
rect 132470 688890 132560 689130
rect 132800 688890 132910 689130
rect 133150 688890 133570 689130
rect 133810 688890 133900 689130
rect 134140 688890 134230 689130
rect 134470 688890 134560 689130
rect 134800 688890 134910 689130
rect 135150 688890 135240 689130
rect 135480 688890 135570 689130
rect 135810 688890 135900 689130
rect 136140 688890 136250 689130
rect 136490 688890 136580 689130
rect 136820 688890 136910 689130
rect 137150 688890 137240 689130
rect 137480 688890 137590 689130
rect 137830 688890 137920 689130
rect 138160 688890 138250 689130
rect 138490 688890 138580 689130
rect 138820 688890 138930 689130
rect 139170 688890 139260 689130
rect 139500 688890 139590 689130
rect 139830 688890 139920 689130
rect 140160 688890 140270 689130
rect 140510 688890 140600 689130
rect 140840 688890 140930 689130
rect 141170 688890 141260 689130
rect 141500 688890 141610 689130
rect 141850 688890 141940 689130
rect 142180 688890 142270 689130
rect 142510 688890 142600 689130
rect 142840 688890 142950 689130
rect 143190 688890 143280 689130
rect 143520 688890 143610 689130
rect 143850 688890 143940 689130
rect 144180 688890 144290 689130
rect 144530 688890 144950 689130
rect 145190 688890 145280 689130
rect 145520 688890 145610 689130
rect 145850 688890 145940 689130
rect 146180 688890 146290 689130
rect 146530 688890 146620 689130
rect 146860 688890 146950 689130
rect 147190 688890 147280 689130
rect 147520 688890 147630 689130
rect 147870 688890 147960 689130
rect 148200 688890 148290 689130
rect 148530 688890 148620 689130
rect 148860 688890 148970 689130
rect 149210 688890 149300 689130
rect 149540 688890 149630 689130
rect 149870 688890 149960 689130
rect 150200 688890 150310 689130
rect 150550 688890 150640 689130
rect 150880 688890 150970 689130
rect 151210 688890 151300 689130
rect 151540 688890 151650 689130
rect 151890 688890 151980 689130
rect 152220 688890 152310 689130
rect 152550 688890 152640 689130
rect 152880 688890 152990 689130
rect 153230 688890 153320 689130
rect 153560 688890 153650 689130
rect 153890 688890 153980 689130
rect 154220 688890 154330 689130
rect 154570 688890 154660 689130
rect 154900 688890 154990 689130
rect 155230 688890 155320 689130
rect 155560 688890 155670 689130
rect 155910 688890 162436 689130
rect 103643 688800 162436 688890
rect 103643 688560 110810 688800
rect 111050 688560 111140 688800
rect 111380 688560 111470 688800
rect 111710 688560 111800 688800
rect 112040 688560 112150 688800
rect 112390 688560 112480 688800
rect 112720 688560 112810 688800
rect 113050 688560 113140 688800
rect 113380 688560 113490 688800
rect 113730 688560 113820 688800
rect 114060 688560 114150 688800
rect 114390 688560 114480 688800
rect 114720 688560 114830 688800
rect 115070 688560 115160 688800
rect 115400 688560 115490 688800
rect 115730 688560 115820 688800
rect 116060 688560 116170 688800
rect 116410 688560 116500 688800
rect 116740 688560 116830 688800
rect 117070 688560 117160 688800
rect 117400 688560 117510 688800
rect 117750 688560 117840 688800
rect 118080 688560 118170 688800
rect 118410 688560 118500 688800
rect 118740 688560 118850 688800
rect 119090 688560 119180 688800
rect 119420 688560 119510 688800
rect 119750 688560 119840 688800
rect 120080 688560 120190 688800
rect 120430 688560 120520 688800
rect 120760 688560 120850 688800
rect 121090 688560 121180 688800
rect 121420 688560 121530 688800
rect 121770 688560 122190 688800
rect 122430 688560 122520 688800
rect 122760 688560 122850 688800
rect 123090 688560 123180 688800
rect 123420 688560 123530 688800
rect 123770 688560 123860 688800
rect 124100 688560 124190 688800
rect 124430 688560 124520 688800
rect 124760 688560 124870 688800
rect 125110 688560 125200 688800
rect 125440 688560 125530 688800
rect 125770 688560 125860 688800
rect 126100 688560 126210 688800
rect 126450 688560 126540 688800
rect 126780 688560 126870 688800
rect 127110 688560 127200 688800
rect 127440 688560 127550 688800
rect 127790 688560 127880 688800
rect 128120 688560 128210 688800
rect 128450 688560 128540 688800
rect 128780 688560 128890 688800
rect 129130 688560 129220 688800
rect 129460 688560 129550 688800
rect 129790 688560 129880 688800
rect 130120 688560 130230 688800
rect 130470 688560 130560 688800
rect 130800 688560 130890 688800
rect 131130 688560 131220 688800
rect 131460 688560 131570 688800
rect 131810 688560 131900 688800
rect 132140 688560 132230 688800
rect 132470 688560 132560 688800
rect 132800 688560 132910 688800
rect 133150 688560 133570 688800
rect 133810 688560 133900 688800
rect 134140 688560 134230 688800
rect 134470 688560 134560 688800
rect 134800 688560 134910 688800
rect 135150 688560 135240 688800
rect 135480 688560 135570 688800
rect 135810 688560 135900 688800
rect 136140 688560 136250 688800
rect 136490 688560 136580 688800
rect 136820 688560 136910 688800
rect 137150 688560 137240 688800
rect 137480 688560 137590 688800
rect 137830 688560 137920 688800
rect 138160 688560 138250 688800
rect 138490 688560 138580 688800
rect 138820 688560 138930 688800
rect 139170 688560 139260 688800
rect 139500 688560 139590 688800
rect 139830 688560 139920 688800
rect 140160 688560 140270 688800
rect 140510 688560 140600 688800
rect 140840 688560 140930 688800
rect 141170 688560 141260 688800
rect 141500 688560 141610 688800
rect 141850 688560 141940 688800
rect 142180 688560 142270 688800
rect 142510 688560 142600 688800
rect 142840 688560 142950 688800
rect 143190 688560 143280 688800
rect 143520 688560 143610 688800
rect 143850 688560 143940 688800
rect 144180 688560 144290 688800
rect 144530 688560 144950 688800
rect 145190 688560 145280 688800
rect 145520 688560 145610 688800
rect 145850 688560 145940 688800
rect 146180 688560 146290 688800
rect 146530 688560 146620 688800
rect 146860 688560 146950 688800
rect 147190 688560 147280 688800
rect 147520 688560 147630 688800
rect 147870 688560 147960 688800
rect 148200 688560 148290 688800
rect 148530 688560 148620 688800
rect 148860 688560 148970 688800
rect 149210 688560 149300 688800
rect 149540 688560 149630 688800
rect 149870 688560 149960 688800
rect 150200 688560 150310 688800
rect 150550 688560 150640 688800
rect 150880 688560 150970 688800
rect 151210 688560 151300 688800
rect 151540 688560 151650 688800
rect 151890 688560 151980 688800
rect 152220 688560 152310 688800
rect 152550 688560 152640 688800
rect 152880 688560 152990 688800
rect 153230 688560 153320 688800
rect 153560 688560 153650 688800
rect 153890 688560 153980 688800
rect 154220 688560 154330 688800
rect 154570 688560 154660 688800
rect 154900 688560 154990 688800
rect 155230 688560 155320 688800
rect 155560 688560 155670 688800
rect 155910 688560 162436 688800
rect 103643 688470 162436 688560
rect 103643 688230 110810 688470
rect 111050 688230 111140 688470
rect 111380 688230 111470 688470
rect 111710 688230 111800 688470
rect 112040 688230 112150 688470
rect 112390 688230 112480 688470
rect 112720 688230 112810 688470
rect 113050 688230 113140 688470
rect 113380 688230 113490 688470
rect 113730 688230 113820 688470
rect 114060 688230 114150 688470
rect 114390 688230 114480 688470
rect 114720 688230 114830 688470
rect 115070 688230 115160 688470
rect 115400 688230 115490 688470
rect 115730 688230 115820 688470
rect 116060 688230 116170 688470
rect 116410 688230 116500 688470
rect 116740 688230 116830 688470
rect 117070 688230 117160 688470
rect 117400 688230 117510 688470
rect 117750 688230 117840 688470
rect 118080 688230 118170 688470
rect 118410 688230 118500 688470
rect 118740 688230 118850 688470
rect 119090 688230 119180 688470
rect 119420 688230 119510 688470
rect 119750 688230 119840 688470
rect 120080 688230 120190 688470
rect 120430 688230 120520 688470
rect 120760 688230 120850 688470
rect 121090 688230 121180 688470
rect 121420 688230 121530 688470
rect 121770 688230 122190 688470
rect 122430 688230 122520 688470
rect 122760 688230 122850 688470
rect 123090 688230 123180 688470
rect 123420 688230 123530 688470
rect 123770 688230 123860 688470
rect 124100 688230 124190 688470
rect 124430 688230 124520 688470
rect 124760 688230 124870 688470
rect 125110 688230 125200 688470
rect 125440 688230 125530 688470
rect 125770 688230 125860 688470
rect 126100 688230 126210 688470
rect 126450 688230 126540 688470
rect 126780 688230 126870 688470
rect 127110 688230 127200 688470
rect 127440 688230 127550 688470
rect 127790 688230 127880 688470
rect 128120 688230 128210 688470
rect 128450 688230 128540 688470
rect 128780 688230 128890 688470
rect 129130 688230 129220 688470
rect 129460 688230 129550 688470
rect 129790 688230 129880 688470
rect 130120 688230 130230 688470
rect 130470 688230 130560 688470
rect 130800 688230 130890 688470
rect 131130 688230 131220 688470
rect 131460 688230 131570 688470
rect 131810 688230 131900 688470
rect 132140 688230 132230 688470
rect 132470 688230 132560 688470
rect 132800 688230 132910 688470
rect 133150 688230 133570 688470
rect 133810 688230 133900 688470
rect 134140 688230 134230 688470
rect 134470 688230 134560 688470
rect 134800 688230 134910 688470
rect 135150 688230 135240 688470
rect 135480 688230 135570 688470
rect 135810 688230 135900 688470
rect 136140 688230 136250 688470
rect 136490 688230 136580 688470
rect 136820 688230 136910 688470
rect 137150 688230 137240 688470
rect 137480 688230 137590 688470
rect 137830 688230 137920 688470
rect 138160 688230 138250 688470
rect 138490 688230 138580 688470
rect 138820 688230 138930 688470
rect 139170 688230 139260 688470
rect 139500 688230 139590 688470
rect 139830 688230 139920 688470
rect 140160 688230 140270 688470
rect 140510 688230 140600 688470
rect 140840 688230 140930 688470
rect 141170 688230 141260 688470
rect 141500 688230 141610 688470
rect 141850 688230 141940 688470
rect 142180 688230 142270 688470
rect 142510 688230 142600 688470
rect 142840 688230 142950 688470
rect 143190 688230 143280 688470
rect 143520 688230 143610 688470
rect 143850 688230 143940 688470
rect 144180 688230 144290 688470
rect 144530 688230 144950 688470
rect 145190 688230 145280 688470
rect 145520 688230 145610 688470
rect 145850 688230 145940 688470
rect 146180 688230 146290 688470
rect 146530 688230 146620 688470
rect 146860 688230 146950 688470
rect 147190 688230 147280 688470
rect 147520 688230 147630 688470
rect 147870 688230 147960 688470
rect 148200 688230 148290 688470
rect 148530 688230 148620 688470
rect 148860 688230 148970 688470
rect 149210 688230 149300 688470
rect 149540 688230 149630 688470
rect 149870 688230 149960 688470
rect 150200 688230 150310 688470
rect 150550 688230 150640 688470
rect 150880 688230 150970 688470
rect 151210 688230 151300 688470
rect 151540 688230 151650 688470
rect 151890 688230 151980 688470
rect 152220 688230 152310 688470
rect 152550 688230 152640 688470
rect 152880 688230 152990 688470
rect 153230 688230 153320 688470
rect 153560 688230 153650 688470
rect 153890 688230 153980 688470
rect 154220 688230 154330 688470
rect 154570 688230 154660 688470
rect 154900 688230 154990 688470
rect 155230 688230 155320 688470
rect 155560 688230 155670 688470
rect 155910 688230 162436 688470
rect 103643 688140 162436 688230
rect 103643 687900 110810 688140
rect 111050 687900 111140 688140
rect 111380 687900 111470 688140
rect 111710 687900 111800 688140
rect 112040 687900 112150 688140
rect 112390 687900 112480 688140
rect 112720 687900 112810 688140
rect 113050 687900 113140 688140
rect 113380 687900 113490 688140
rect 113730 687900 113820 688140
rect 114060 687900 114150 688140
rect 114390 687900 114480 688140
rect 114720 687900 114830 688140
rect 115070 687900 115160 688140
rect 115400 687900 115490 688140
rect 115730 687900 115820 688140
rect 116060 687900 116170 688140
rect 116410 687900 116500 688140
rect 116740 687900 116830 688140
rect 117070 687900 117160 688140
rect 117400 687900 117510 688140
rect 117750 687900 117840 688140
rect 118080 687900 118170 688140
rect 118410 687900 118500 688140
rect 118740 687900 118850 688140
rect 119090 687900 119180 688140
rect 119420 687900 119510 688140
rect 119750 687900 119840 688140
rect 120080 687900 120190 688140
rect 120430 687900 120520 688140
rect 120760 687900 120850 688140
rect 121090 687900 121180 688140
rect 121420 687900 121530 688140
rect 121770 687900 122190 688140
rect 122430 687900 122520 688140
rect 122760 687900 122850 688140
rect 123090 687900 123180 688140
rect 123420 687900 123530 688140
rect 123770 687900 123860 688140
rect 124100 687900 124190 688140
rect 124430 687900 124520 688140
rect 124760 687900 124870 688140
rect 125110 687900 125200 688140
rect 125440 687900 125530 688140
rect 125770 687900 125860 688140
rect 126100 687900 126210 688140
rect 126450 687900 126540 688140
rect 126780 687900 126870 688140
rect 127110 687900 127200 688140
rect 127440 687900 127550 688140
rect 127790 687900 127880 688140
rect 128120 687900 128210 688140
rect 128450 687900 128540 688140
rect 128780 687900 128890 688140
rect 129130 687900 129220 688140
rect 129460 687900 129550 688140
rect 129790 687900 129880 688140
rect 130120 687900 130230 688140
rect 130470 687900 130560 688140
rect 130800 687900 130890 688140
rect 131130 687900 131220 688140
rect 131460 687900 131570 688140
rect 131810 687900 131900 688140
rect 132140 687900 132230 688140
rect 132470 687900 132560 688140
rect 132800 687900 132910 688140
rect 133150 687900 133570 688140
rect 133810 687900 133900 688140
rect 134140 687900 134230 688140
rect 134470 687900 134560 688140
rect 134800 687900 134910 688140
rect 135150 687900 135240 688140
rect 135480 687900 135570 688140
rect 135810 687900 135900 688140
rect 136140 687900 136250 688140
rect 136490 687900 136580 688140
rect 136820 687900 136910 688140
rect 137150 687900 137240 688140
rect 137480 687900 137590 688140
rect 137830 687900 137920 688140
rect 138160 687900 138250 688140
rect 138490 687900 138580 688140
rect 138820 687900 138930 688140
rect 139170 687900 139260 688140
rect 139500 687900 139590 688140
rect 139830 687900 139920 688140
rect 140160 687900 140270 688140
rect 140510 687900 140600 688140
rect 140840 687900 140930 688140
rect 141170 687900 141260 688140
rect 141500 687900 141610 688140
rect 141850 687900 141940 688140
rect 142180 687900 142270 688140
rect 142510 687900 142600 688140
rect 142840 687900 142950 688140
rect 143190 687900 143280 688140
rect 143520 687900 143610 688140
rect 143850 687900 143940 688140
rect 144180 687900 144290 688140
rect 144530 687900 144950 688140
rect 145190 687900 145280 688140
rect 145520 687900 145610 688140
rect 145850 687900 145940 688140
rect 146180 687900 146290 688140
rect 146530 687900 146620 688140
rect 146860 687900 146950 688140
rect 147190 687900 147280 688140
rect 147520 687900 147630 688140
rect 147870 687900 147960 688140
rect 148200 687900 148290 688140
rect 148530 687900 148620 688140
rect 148860 687900 148970 688140
rect 149210 687900 149300 688140
rect 149540 687900 149630 688140
rect 149870 687900 149960 688140
rect 150200 687900 150310 688140
rect 150550 687900 150640 688140
rect 150880 687900 150970 688140
rect 151210 687900 151300 688140
rect 151540 687900 151650 688140
rect 151890 687900 151980 688140
rect 152220 687900 152310 688140
rect 152550 687900 152640 688140
rect 152880 687900 152990 688140
rect 153230 687900 153320 688140
rect 153560 687900 153650 688140
rect 153890 687900 153980 688140
rect 154220 687900 154330 688140
rect 154570 687900 154660 688140
rect 154900 687900 154990 688140
rect 155230 687900 155320 688140
rect 155560 687900 155670 688140
rect 155910 687900 162436 688140
rect 103643 687790 162436 687900
rect 103643 687550 110810 687790
rect 111050 687550 111140 687790
rect 111380 687550 111470 687790
rect 111710 687550 111800 687790
rect 112040 687550 112150 687790
rect 112390 687550 112480 687790
rect 112720 687550 112810 687790
rect 113050 687550 113140 687790
rect 113380 687550 113490 687790
rect 113730 687550 113820 687790
rect 114060 687550 114150 687790
rect 114390 687550 114480 687790
rect 114720 687550 114830 687790
rect 115070 687550 115160 687790
rect 115400 687550 115490 687790
rect 115730 687550 115820 687790
rect 116060 687550 116170 687790
rect 116410 687550 116500 687790
rect 116740 687550 116830 687790
rect 117070 687550 117160 687790
rect 117400 687550 117510 687790
rect 117750 687550 117840 687790
rect 118080 687550 118170 687790
rect 118410 687550 118500 687790
rect 118740 687550 118850 687790
rect 119090 687550 119180 687790
rect 119420 687550 119510 687790
rect 119750 687550 119840 687790
rect 120080 687550 120190 687790
rect 120430 687550 120520 687790
rect 120760 687550 120850 687790
rect 121090 687550 121180 687790
rect 121420 687550 121530 687790
rect 121770 687550 122190 687790
rect 122430 687550 122520 687790
rect 122760 687550 122850 687790
rect 123090 687550 123180 687790
rect 123420 687550 123530 687790
rect 123770 687550 123860 687790
rect 124100 687550 124190 687790
rect 124430 687550 124520 687790
rect 124760 687550 124870 687790
rect 125110 687550 125200 687790
rect 125440 687550 125530 687790
rect 125770 687550 125860 687790
rect 126100 687550 126210 687790
rect 126450 687550 126540 687790
rect 126780 687550 126870 687790
rect 127110 687550 127200 687790
rect 127440 687550 127550 687790
rect 127790 687550 127880 687790
rect 128120 687550 128210 687790
rect 128450 687550 128540 687790
rect 128780 687550 128890 687790
rect 129130 687550 129220 687790
rect 129460 687550 129550 687790
rect 129790 687550 129880 687790
rect 130120 687550 130230 687790
rect 130470 687550 130560 687790
rect 130800 687550 130890 687790
rect 131130 687550 131220 687790
rect 131460 687550 131570 687790
rect 131810 687550 131900 687790
rect 132140 687550 132230 687790
rect 132470 687550 132560 687790
rect 132800 687550 132910 687790
rect 133150 687550 133570 687790
rect 133810 687550 133900 687790
rect 134140 687550 134230 687790
rect 134470 687550 134560 687790
rect 134800 687550 134910 687790
rect 135150 687550 135240 687790
rect 135480 687550 135570 687790
rect 135810 687550 135900 687790
rect 136140 687550 136250 687790
rect 136490 687550 136580 687790
rect 136820 687550 136910 687790
rect 137150 687550 137240 687790
rect 137480 687550 137590 687790
rect 137830 687550 137920 687790
rect 138160 687550 138250 687790
rect 138490 687550 138580 687790
rect 138820 687550 138930 687790
rect 139170 687550 139260 687790
rect 139500 687550 139590 687790
rect 139830 687550 139920 687790
rect 140160 687550 140270 687790
rect 140510 687550 140600 687790
rect 140840 687550 140930 687790
rect 141170 687550 141260 687790
rect 141500 687550 141610 687790
rect 141850 687550 141940 687790
rect 142180 687550 142270 687790
rect 142510 687550 142600 687790
rect 142840 687550 142950 687790
rect 143190 687550 143280 687790
rect 143520 687550 143610 687790
rect 143850 687550 143940 687790
rect 144180 687550 144290 687790
rect 144530 687550 144950 687790
rect 145190 687550 145280 687790
rect 145520 687550 145610 687790
rect 145850 687550 145940 687790
rect 146180 687550 146290 687790
rect 146530 687550 146620 687790
rect 146860 687550 146950 687790
rect 147190 687550 147280 687790
rect 147520 687550 147630 687790
rect 147870 687550 147960 687790
rect 148200 687550 148290 687790
rect 148530 687550 148620 687790
rect 148860 687550 148970 687790
rect 149210 687550 149300 687790
rect 149540 687550 149630 687790
rect 149870 687550 149960 687790
rect 150200 687550 150310 687790
rect 150550 687550 150640 687790
rect 150880 687550 150970 687790
rect 151210 687550 151300 687790
rect 151540 687550 151650 687790
rect 151890 687550 151980 687790
rect 152220 687550 152310 687790
rect 152550 687550 152640 687790
rect 152880 687550 152990 687790
rect 153230 687550 153320 687790
rect 153560 687550 153650 687790
rect 153890 687550 153980 687790
rect 154220 687550 154330 687790
rect 154570 687550 154660 687790
rect 154900 687550 154990 687790
rect 155230 687550 155320 687790
rect 155560 687550 155670 687790
rect 155910 687550 162436 687790
rect 103643 687460 162436 687550
rect 103643 687220 110810 687460
rect 111050 687220 111140 687460
rect 111380 687220 111470 687460
rect 111710 687220 111800 687460
rect 112040 687220 112150 687460
rect 112390 687220 112480 687460
rect 112720 687220 112810 687460
rect 113050 687220 113140 687460
rect 113380 687220 113490 687460
rect 113730 687220 113820 687460
rect 114060 687220 114150 687460
rect 114390 687220 114480 687460
rect 114720 687220 114830 687460
rect 115070 687220 115160 687460
rect 115400 687220 115490 687460
rect 115730 687220 115820 687460
rect 116060 687220 116170 687460
rect 116410 687220 116500 687460
rect 116740 687220 116830 687460
rect 117070 687220 117160 687460
rect 117400 687220 117510 687460
rect 117750 687220 117840 687460
rect 118080 687220 118170 687460
rect 118410 687220 118500 687460
rect 118740 687220 118850 687460
rect 119090 687220 119180 687460
rect 119420 687220 119510 687460
rect 119750 687220 119840 687460
rect 120080 687220 120190 687460
rect 120430 687220 120520 687460
rect 120760 687220 120850 687460
rect 121090 687220 121180 687460
rect 121420 687220 121530 687460
rect 121770 687220 122190 687460
rect 122430 687220 122520 687460
rect 122760 687220 122850 687460
rect 123090 687220 123180 687460
rect 123420 687220 123530 687460
rect 123770 687220 123860 687460
rect 124100 687220 124190 687460
rect 124430 687220 124520 687460
rect 124760 687220 124870 687460
rect 125110 687220 125200 687460
rect 125440 687220 125530 687460
rect 125770 687220 125860 687460
rect 126100 687220 126210 687460
rect 126450 687220 126540 687460
rect 126780 687220 126870 687460
rect 127110 687220 127200 687460
rect 127440 687220 127550 687460
rect 127790 687220 127880 687460
rect 128120 687220 128210 687460
rect 128450 687220 128540 687460
rect 128780 687220 128890 687460
rect 129130 687220 129220 687460
rect 129460 687220 129550 687460
rect 129790 687220 129880 687460
rect 130120 687220 130230 687460
rect 130470 687220 130560 687460
rect 130800 687220 130890 687460
rect 131130 687220 131220 687460
rect 131460 687220 131570 687460
rect 131810 687220 131900 687460
rect 132140 687220 132230 687460
rect 132470 687220 132560 687460
rect 132800 687220 132910 687460
rect 133150 687220 133570 687460
rect 133810 687220 133900 687460
rect 134140 687220 134230 687460
rect 134470 687220 134560 687460
rect 134800 687220 134910 687460
rect 135150 687220 135240 687460
rect 135480 687220 135570 687460
rect 135810 687220 135900 687460
rect 136140 687220 136250 687460
rect 136490 687220 136580 687460
rect 136820 687220 136910 687460
rect 137150 687220 137240 687460
rect 137480 687220 137590 687460
rect 137830 687220 137920 687460
rect 138160 687220 138250 687460
rect 138490 687220 138580 687460
rect 138820 687220 138930 687460
rect 139170 687220 139260 687460
rect 139500 687220 139590 687460
rect 139830 687220 139920 687460
rect 140160 687220 140270 687460
rect 140510 687220 140600 687460
rect 140840 687220 140930 687460
rect 141170 687220 141260 687460
rect 141500 687220 141610 687460
rect 141850 687220 141940 687460
rect 142180 687220 142270 687460
rect 142510 687220 142600 687460
rect 142840 687220 142950 687460
rect 143190 687220 143280 687460
rect 143520 687220 143610 687460
rect 143850 687220 143940 687460
rect 144180 687220 144290 687460
rect 144530 687220 144950 687460
rect 145190 687220 145280 687460
rect 145520 687220 145610 687460
rect 145850 687220 145940 687460
rect 146180 687220 146290 687460
rect 146530 687220 146620 687460
rect 146860 687220 146950 687460
rect 147190 687220 147280 687460
rect 147520 687220 147630 687460
rect 147870 687220 147960 687460
rect 148200 687220 148290 687460
rect 148530 687220 148620 687460
rect 148860 687220 148970 687460
rect 149210 687220 149300 687460
rect 149540 687220 149630 687460
rect 149870 687220 149960 687460
rect 150200 687220 150310 687460
rect 150550 687220 150640 687460
rect 150880 687220 150970 687460
rect 151210 687220 151300 687460
rect 151540 687220 151650 687460
rect 151890 687220 151980 687460
rect 152220 687220 152310 687460
rect 152550 687220 152640 687460
rect 152880 687220 152990 687460
rect 153230 687220 153320 687460
rect 153560 687220 153650 687460
rect 153890 687220 153980 687460
rect 154220 687220 154330 687460
rect 154570 687220 154660 687460
rect 154900 687220 154990 687460
rect 155230 687220 155320 687460
rect 155560 687220 155670 687460
rect 155910 687220 162436 687460
rect 103643 687130 162436 687220
rect 103643 686890 110810 687130
rect 111050 686890 111140 687130
rect 111380 686890 111470 687130
rect 111710 686890 111800 687130
rect 112040 686890 112150 687130
rect 112390 686890 112480 687130
rect 112720 686890 112810 687130
rect 113050 686890 113140 687130
rect 113380 686890 113490 687130
rect 113730 686890 113820 687130
rect 114060 686890 114150 687130
rect 114390 686890 114480 687130
rect 114720 686890 114830 687130
rect 115070 686890 115160 687130
rect 115400 686890 115490 687130
rect 115730 686890 115820 687130
rect 116060 686890 116170 687130
rect 116410 686890 116500 687130
rect 116740 686890 116830 687130
rect 117070 686890 117160 687130
rect 117400 686890 117510 687130
rect 117750 686890 117840 687130
rect 118080 686890 118170 687130
rect 118410 686890 118500 687130
rect 118740 686890 118850 687130
rect 119090 686890 119180 687130
rect 119420 686890 119510 687130
rect 119750 686890 119840 687130
rect 120080 686890 120190 687130
rect 120430 686890 120520 687130
rect 120760 686890 120850 687130
rect 121090 686890 121180 687130
rect 121420 686890 121530 687130
rect 121770 686890 122190 687130
rect 122430 686890 122520 687130
rect 122760 686890 122850 687130
rect 123090 686890 123180 687130
rect 123420 686890 123530 687130
rect 123770 686890 123860 687130
rect 124100 686890 124190 687130
rect 124430 686890 124520 687130
rect 124760 686890 124870 687130
rect 125110 686890 125200 687130
rect 125440 686890 125530 687130
rect 125770 686890 125860 687130
rect 126100 686890 126210 687130
rect 126450 686890 126540 687130
rect 126780 686890 126870 687130
rect 127110 686890 127200 687130
rect 127440 686890 127550 687130
rect 127790 686890 127880 687130
rect 128120 686890 128210 687130
rect 128450 686890 128540 687130
rect 128780 686890 128890 687130
rect 129130 686890 129220 687130
rect 129460 686890 129550 687130
rect 129790 686890 129880 687130
rect 130120 686890 130230 687130
rect 130470 686890 130560 687130
rect 130800 686890 130890 687130
rect 131130 686890 131220 687130
rect 131460 686890 131570 687130
rect 131810 686890 131900 687130
rect 132140 686890 132230 687130
rect 132470 686890 132560 687130
rect 132800 686890 132910 687130
rect 133150 686890 133570 687130
rect 133810 686890 133900 687130
rect 134140 686890 134230 687130
rect 134470 686890 134560 687130
rect 134800 686890 134910 687130
rect 135150 686890 135240 687130
rect 135480 686890 135570 687130
rect 135810 686890 135900 687130
rect 136140 686890 136250 687130
rect 136490 686890 136580 687130
rect 136820 686890 136910 687130
rect 137150 686890 137240 687130
rect 137480 686890 137590 687130
rect 137830 686890 137920 687130
rect 138160 686890 138250 687130
rect 138490 686890 138580 687130
rect 138820 686890 138930 687130
rect 139170 686890 139260 687130
rect 139500 686890 139590 687130
rect 139830 686890 139920 687130
rect 140160 686890 140270 687130
rect 140510 686890 140600 687130
rect 140840 686890 140930 687130
rect 141170 686890 141260 687130
rect 141500 686890 141610 687130
rect 141850 686890 141940 687130
rect 142180 686890 142270 687130
rect 142510 686890 142600 687130
rect 142840 686890 142950 687130
rect 143190 686890 143280 687130
rect 143520 686890 143610 687130
rect 143850 686890 143940 687130
rect 144180 686890 144290 687130
rect 144530 686890 144950 687130
rect 145190 686890 145280 687130
rect 145520 686890 145610 687130
rect 145850 686890 145940 687130
rect 146180 686890 146290 687130
rect 146530 686890 146620 687130
rect 146860 686890 146950 687130
rect 147190 686890 147280 687130
rect 147520 686890 147630 687130
rect 147870 686890 147960 687130
rect 148200 686890 148290 687130
rect 148530 686890 148620 687130
rect 148860 686890 148970 687130
rect 149210 686890 149300 687130
rect 149540 686890 149630 687130
rect 149870 686890 149960 687130
rect 150200 686890 150310 687130
rect 150550 686890 150640 687130
rect 150880 686890 150970 687130
rect 151210 686890 151300 687130
rect 151540 686890 151650 687130
rect 151890 686890 151980 687130
rect 152220 686890 152310 687130
rect 152550 686890 152640 687130
rect 152880 686890 152990 687130
rect 153230 686890 153320 687130
rect 153560 686890 153650 687130
rect 153890 686890 153980 687130
rect 154220 686890 154330 687130
rect 154570 686890 154660 687130
rect 154900 686890 154990 687130
rect 155230 686890 155320 687130
rect 155560 686890 155670 687130
rect 155910 686890 162436 687130
rect 103643 686800 162436 686890
rect 103643 686560 110810 686800
rect 111050 686560 111140 686800
rect 111380 686560 111470 686800
rect 111710 686560 111800 686800
rect 112040 686560 112150 686800
rect 112390 686560 112480 686800
rect 112720 686560 112810 686800
rect 113050 686560 113140 686800
rect 113380 686560 113490 686800
rect 113730 686560 113820 686800
rect 114060 686560 114150 686800
rect 114390 686560 114480 686800
rect 114720 686560 114830 686800
rect 115070 686560 115160 686800
rect 115400 686560 115490 686800
rect 115730 686560 115820 686800
rect 116060 686560 116170 686800
rect 116410 686560 116500 686800
rect 116740 686560 116830 686800
rect 117070 686560 117160 686800
rect 117400 686560 117510 686800
rect 117750 686560 117840 686800
rect 118080 686560 118170 686800
rect 118410 686560 118500 686800
rect 118740 686560 118850 686800
rect 119090 686560 119180 686800
rect 119420 686560 119510 686800
rect 119750 686560 119840 686800
rect 120080 686560 120190 686800
rect 120430 686560 120520 686800
rect 120760 686560 120850 686800
rect 121090 686560 121180 686800
rect 121420 686560 121530 686800
rect 121770 686560 122190 686800
rect 122430 686560 122520 686800
rect 122760 686560 122850 686800
rect 123090 686560 123180 686800
rect 123420 686560 123530 686800
rect 123770 686560 123860 686800
rect 124100 686560 124190 686800
rect 124430 686560 124520 686800
rect 124760 686560 124870 686800
rect 125110 686560 125200 686800
rect 125440 686560 125530 686800
rect 125770 686560 125860 686800
rect 126100 686560 126210 686800
rect 126450 686560 126540 686800
rect 126780 686560 126870 686800
rect 127110 686560 127200 686800
rect 127440 686560 127550 686800
rect 127790 686560 127880 686800
rect 128120 686560 128210 686800
rect 128450 686560 128540 686800
rect 128780 686560 128890 686800
rect 129130 686560 129220 686800
rect 129460 686560 129550 686800
rect 129790 686560 129880 686800
rect 130120 686560 130230 686800
rect 130470 686560 130560 686800
rect 130800 686560 130890 686800
rect 131130 686560 131220 686800
rect 131460 686560 131570 686800
rect 131810 686560 131900 686800
rect 132140 686560 132230 686800
rect 132470 686560 132560 686800
rect 132800 686560 132910 686800
rect 133150 686560 133570 686800
rect 133810 686560 133900 686800
rect 134140 686560 134230 686800
rect 134470 686560 134560 686800
rect 134800 686560 134910 686800
rect 135150 686560 135240 686800
rect 135480 686560 135570 686800
rect 135810 686560 135900 686800
rect 136140 686560 136250 686800
rect 136490 686560 136580 686800
rect 136820 686560 136910 686800
rect 137150 686560 137240 686800
rect 137480 686560 137590 686800
rect 137830 686560 137920 686800
rect 138160 686560 138250 686800
rect 138490 686560 138580 686800
rect 138820 686560 138930 686800
rect 139170 686560 139260 686800
rect 139500 686560 139590 686800
rect 139830 686560 139920 686800
rect 140160 686560 140270 686800
rect 140510 686560 140600 686800
rect 140840 686560 140930 686800
rect 141170 686560 141260 686800
rect 141500 686560 141610 686800
rect 141850 686560 141940 686800
rect 142180 686560 142270 686800
rect 142510 686560 142600 686800
rect 142840 686560 142950 686800
rect 143190 686560 143280 686800
rect 143520 686560 143610 686800
rect 143850 686560 143940 686800
rect 144180 686560 144290 686800
rect 144530 686560 144950 686800
rect 145190 686560 145280 686800
rect 145520 686560 145610 686800
rect 145850 686560 145940 686800
rect 146180 686560 146290 686800
rect 146530 686560 146620 686800
rect 146860 686560 146950 686800
rect 147190 686560 147280 686800
rect 147520 686560 147630 686800
rect 147870 686560 147960 686800
rect 148200 686560 148290 686800
rect 148530 686560 148620 686800
rect 148860 686560 148970 686800
rect 149210 686560 149300 686800
rect 149540 686560 149630 686800
rect 149870 686560 149960 686800
rect 150200 686560 150310 686800
rect 150550 686560 150640 686800
rect 150880 686560 150970 686800
rect 151210 686560 151300 686800
rect 151540 686560 151650 686800
rect 151890 686560 151980 686800
rect 152220 686560 152310 686800
rect 152550 686560 152640 686800
rect 152880 686560 152990 686800
rect 153230 686560 153320 686800
rect 153560 686560 153650 686800
rect 153890 686560 153980 686800
rect 154220 686560 154330 686800
rect 154570 686560 154660 686800
rect 154900 686560 154990 686800
rect 155230 686560 155320 686800
rect 155560 686560 155670 686800
rect 155910 686560 162436 686800
rect 103643 686450 162436 686560
rect 103643 686210 110810 686450
rect 111050 686210 111140 686450
rect 111380 686210 111470 686450
rect 111710 686210 111800 686450
rect 112040 686210 112150 686450
rect 112390 686210 112480 686450
rect 112720 686210 112810 686450
rect 113050 686210 113140 686450
rect 113380 686210 113490 686450
rect 113730 686210 113820 686450
rect 114060 686210 114150 686450
rect 114390 686210 114480 686450
rect 114720 686210 114830 686450
rect 115070 686210 115160 686450
rect 115400 686210 115490 686450
rect 115730 686210 115820 686450
rect 116060 686210 116170 686450
rect 116410 686210 116500 686450
rect 116740 686210 116830 686450
rect 117070 686210 117160 686450
rect 117400 686210 117510 686450
rect 117750 686210 117840 686450
rect 118080 686210 118170 686450
rect 118410 686210 118500 686450
rect 118740 686210 118850 686450
rect 119090 686210 119180 686450
rect 119420 686210 119510 686450
rect 119750 686210 119840 686450
rect 120080 686210 120190 686450
rect 120430 686210 120520 686450
rect 120760 686210 120850 686450
rect 121090 686210 121180 686450
rect 121420 686210 121530 686450
rect 121770 686210 122190 686450
rect 122430 686210 122520 686450
rect 122760 686210 122850 686450
rect 123090 686210 123180 686450
rect 123420 686210 123530 686450
rect 123770 686210 123860 686450
rect 124100 686210 124190 686450
rect 124430 686210 124520 686450
rect 124760 686210 124870 686450
rect 125110 686210 125200 686450
rect 125440 686210 125530 686450
rect 125770 686210 125860 686450
rect 126100 686210 126210 686450
rect 126450 686210 126540 686450
rect 126780 686210 126870 686450
rect 127110 686210 127200 686450
rect 127440 686210 127550 686450
rect 127790 686210 127880 686450
rect 128120 686210 128210 686450
rect 128450 686210 128540 686450
rect 128780 686210 128890 686450
rect 129130 686210 129220 686450
rect 129460 686210 129550 686450
rect 129790 686210 129880 686450
rect 130120 686210 130230 686450
rect 130470 686210 130560 686450
rect 130800 686210 130890 686450
rect 131130 686210 131220 686450
rect 131460 686210 131570 686450
rect 131810 686210 131900 686450
rect 132140 686210 132230 686450
rect 132470 686210 132560 686450
rect 132800 686210 132910 686450
rect 133150 686210 133570 686450
rect 133810 686210 133900 686450
rect 134140 686210 134230 686450
rect 134470 686210 134560 686450
rect 134800 686210 134910 686450
rect 135150 686210 135240 686450
rect 135480 686210 135570 686450
rect 135810 686210 135900 686450
rect 136140 686210 136250 686450
rect 136490 686210 136580 686450
rect 136820 686210 136910 686450
rect 137150 686210 137240 686450
rect 137480 686210 137590 686450
rect 137830 686210 137920 686450
rect 138160 686210 138250 686450
rect 138490 686210 138580 686450
rect 138820 686210 138930 686450
rect 139170 686210 139260 686450
rect 139500 686210 139590 686450
rect 139830 686210 139920 686450
rect 140160 686210 140270 686450
rect 140510 686210 140600 686450
rect 140840 686210 140930 686450
rect 141170 686210 141260 686450
rect 141500 686210 141610 686450
rect 141850 686210 141940 686450
rect 142180 686210 142270 686450
rect 142510 686210 142600 686450
rect 142840 686210 142950 686450
rect 143190 686210 143280 686450
rect 143520 686210 143610 686450
rect 143850 686210 143940 686450
rect 144180 686210 144290 686450
rect 144530 686210 144950 686450
rect 145190 686210 145280 686450
rect 145520 686210 145610 686450
rect 145850 686210 145940 686450
rect 146180 686210 146290 686450
rect 146530 686210 146620 686450
rect 146860 686210 146950 686450
rect 147190 686210 147280 686450
rect 147520 686210 147630 686450
rect 147870 686210 147960 686450
rect 148200 686210 148290 686450
rect 148530 686210 148620 686450
rect 148860 686210 148970 686450
rect 149210 686210 149300 686450
rect 149540 686210 149630 686450
rect 149870 686210 149960 686450
rect 150200 686210 150310 686450
rect 150550 686210 150640 686450
rect 150880 686210 150970 686450
rect 151210 686210 151300 686450
rect 151540 686210 151650 686450
rect 151890 686210 151980 686450
rect 152220 686210 152310 686450
rect 152550 686210 152640 686450
rect 152880 686210 152990 686450
rect 153230 686210 153320 686450
rect 153560 686210 153650 686450
rect 153890 686210 153980 686450
rect 154220 686210 154330 686450
rect 154570 686210 154660 686450
rect 154900 686210 154990 686450
rect 155230 686210 155320 686450
rect 155560 686210 155670 686450
rect 155910 686210 162436 686450
rect 103643 686120 162436 686210
rect 103643 686032 110810 686120
rect 103643 679147 108640 686032
rect 110760 685880 110810 686032
rect 111050 685880 111140 686120
rect 111380 685880 111470 686120
rect 111710 685880 111800 686120
rect 112040 685880 112150 686120
rect 112390 685880 112480 686120
rect 112720 685880 112810 686120
rect 113050 685880 113140 686120
rect 113380 685880 113490 686120
rect 113730 685880 113820 686120
rect 114060 685880 114150 686120
rect 114390 685880 114480 686120
rect 114720 685880 114830 686120
rect 115070 685880 115160 686120
rect 115400 685880 115490 686120
rect 115730 685880 115820 686120
rect 116060 685880 116170 686120
rect 116410 685880 116500 686120
rect 116740 685880 116830 686120
rect 117070 685880 117160 686120
rect 117400 685880 117510 686120
rect 117750 685880 117840 686120
rect 118080 685880 118170 686120
rect 118410 685880 118500 686120
rect 118740 685880 118850 686120
rect 119090 685880 119180 686120
rect 119420 685880 119510 686120
rect 119750 685880 119840 686120
rect 120080 685880 120190 686120
rect 120430 685880 120520 686120
rect 120760 685880 120850 686120
rect 121090 685880 121180 686120
rect 121420 685880 121530 686120
rect 121770 685880 122190 686120
rect 122430 685880 122520 686120
rect 122760 685880 122850 686120
rect 123090 685880 123180 686120
rect 123420 685880 123530 686120
rect 123770 685880 123860 686120
rect 124100 685880 124190 686120
rect 124430 685880 124520 686120
rect 124760 685880 124870 686120
rect 125110 685880 125200 686120
rect 125440 685880 125530 686120
rect 125770 685880 125860 686120
rect 126100 685880 126210 686120
rect 126450 685880 126540 686120
rect 126780 685880 126870 686120
rect 127110 685880 127200 686120
rect 127440 685880 127550 686120
rect 127790 685880 127880 686120
rect 128120 685880 128210 686120
rect 128450 685880 128540 686120
rect 128780 685880 128890 686120
rect 129130 685880 129220 686120
rect 129460 685880 129550 686120
rect 129790 685880 129880 686120
rect 130120 685880 130230 686120
rect 130470 685880 130560 686120
rect 130800 685880 130890 686120
rect 131130 685880 131220 686120
rect 131460 685880 131570 686120
rect 131810 685880 131900 686120
rect 132140 685880 132230 686120
rect 132470 685880 132560 686120
rect 132800 685880 132910 686120
rect 133150 685880 133570 686120
rect 133810 685880 133900 686120
rect 134140 685880 134230 686120
rect 134470 685880 134560 686120
rect 134800 685880 134910 686120
rect 135150 685880 135240 686120
rect 135480 685880 135570 686120
rect 135810 685880 135900 686120
rect 136140 685880 136250 686120
rect 136490 685880 136580 686120
rect 136820 685880 136910 686120
rect 137150 685880 137240 686120
rect 137480 685880 137590 686120
rect 137830 685880 137920 686120
rect 138160 685880 138250 686120
rect 138490 685880 138580 686120
rect 138820 685880 138930 686120
rect 139170 685880 139260 686120
rect 139500 685880 139590 686120
rect 139830 685880 139920 686120
rect 140160 685880 140270 686120
rect 140510 685880 140600 686120
rect 140840 685880 140930 686120
rect 141170 685880 141260 686120
rect 141500 685880 141610 686120
rect 141850 685880 141940 686120
rect 142180 685880 142270 686120
rect 142510 685880 142600 686120
rect 142840 685880 142950 686120
rect 143190 685880 143280 686120
rect 143520 685880 143610 686120
rect 143850 685880 143940 686120
rect 144180 685880 144290 686120
rect 144530 685880 144950 686120
rect 145190 685880 145280 686120
rect 145520 685880 145610 686120
rect 145850 685880 145940 686120
rect 146180 685880 146290 686120
rect 146530 685880 146620 686120
rect 146860 685880 146950 686120
rect 147190 685880 147280 686120
rect 147520 685880 147630 686120
rect 147870 685880 147960 686120
rect 148200 685880 148290 686120
rect 148530 685880 148620 686120
rect 148860 685880 148970 686120
rect 149210 685880 149300 686120
rect 149540 685880 149630 686120
rect 149870 685880 149960 686120
rect 150200 685880 150310 686120
rect 150550 685880 150640 686120
rect 150880 685880 150970 686120
rect 151210 685880 151300 686120
rect 151540 685880 151650 686120
rect 151890 685880 151980 686120
rect 152220 685880 152310 686120
rect 152550 685880 152640 686120
rect 152880 685880 152990 686120
rect 153230 685880 153320 686120
rect 153560 685880 153650 686120
rect 153890 685880 153980 686120
rect 154220 685880 154330 686120
rect 154570 685880 154660 686120
rect 154900 685880 154990 686120
rect 155230 685880 155320 686120
rect 155560 685880 155670 686120
rect 155910 686032 162436 686120
rect 155910 685880 155960 686032
rect 110760 685790 155960 685880
rect 110760 685550 110810 685790
rect 111050 685550 111140 685790
rect 111380 685550 111470 685790
rect 111710 685550 111800 685790
rect 112040 685550 112150 685790
rect 112390 685550 112480 685790
rect 112720 685550 112810 685790
rect 113050 685550 113140 685790
rect 113380 685550 113490 685790
rect 113730 685550 113820 685790
rect 114060 685550 114150 685790
rect 114390 685550 114480 685790
rect 114720 685550 114830 685790
rect 115070 685550 115160 685790
rect 115400 685550 115490 685790
rect 115730 685550 115820 685790
rect 116060 685550 116170 685790
rect 116410 685550 116500 685790
rect 116740 685550 116830 685790
rect 117070 685550 117160 685790
rect 117400 685550 117510 685790
rect 117750 685550 117840 685790
rect 118080 685550 118170 685790
rect 118410 685550 118500 685790
rect 118740 685550 118850 685790
rect 119090 685550 119180 685790
rect 119420 685550 119510 685790
rect 119750 685550 119840 685790
rect 120080 685550 120190 685790
rect 120430 685550 120520 685790
rect 120760 685550 120850 685790
rect 121090 685550 121180 685790
rect 121420 685550 121530 685790
rect 121770 685550 122190 685790
rect 122430 685550 122520 685790
rect 122760 685550 122850 685790
rect 123090 685550 123180 685790
rect 123420 685550 123530 685790
rect 123770 685550 123860 685790
rect 124100 685550 124190 685790
rect 124430 685550 124520 685790
rect 124760 685550 124870 685790
rect 125110 685550 125200 685790
rect 125440 685550 125530 685790
rect 125770 685550 125860 685790
rect 126100 685550 126210 685790
rect 126450 685550 126540 685790
rect 126780 685550 126870 685790
rect 127110 685550 127200 685790
rect 127440 685550 127550 685790
rect 127790 685550 127880 685790
rect 128120 685550 128210 685790
rect 128450 685550 128540 685790
rect 128780 685550 128890 685790
rect 129130 685550 129220 685790
rect 129460 685550 129550 685790
rect 129790 685550 129880 685790
rect 130120 685550 130230 685790
rect 130470 685550 130560 685790
rect 130800 685550 130890 685790
rect 131130 685550 131220 685790
rect 131460 685550 131570 685790
rect 131810 685550 131900 685790
rect 132140 685550 132230 685790
rect 132470 685550 132560 685790
rect 132800 685550 132910 685790
rect 133150 685550 133570 685790
rect 133810 685550 133900 685790
rect 134140 685550 134230 685790
rect 134470 685550 134560 685790
rect 134800 685550 134910 685790
rect 135150 685550 135240 685790
rect 135480 685550 135570 685790
rect 135810 685550 135900 685790
rect 136140 685550 136250 685790
rect 136490 685550 136580 685790
rect 136820 685550 136910 685790
rect 137150 685550 137240 685790
rect 137480 685550 137590 685790
rect 137830 685550 137920 685790
rect 138160 685550 138250 685790
rect 138490 685550 138580 685790
rect 138820 685550 138930 685790
rect 139170 685550 139260 685790
rect 139500 685550 139590 685790
rect 139830 685550 139920 685790
rect 140160 685550 140270 685790
rect 140510 685550 140600 685790
rect 140840 685550 140930 685790
rect 141170 685550 141260 685790
rect 141500 685550 141610 685790
rect 141850 685550 141940 685790
rect 142180 685550 142270 685790
rect 142510 685550 142600 685790
rect 142840 685550 142950 685790
rect 143190 685550 143280 685790
rect 143520 685550 143610 685790
rect 143850 685550 143940 685790
rect 144180 685550 144290 685790
rect 144530 685550 144950 685790
rect 145190 685550 145280 685790
rect 145520 685550 145610 685790
rect 145850 685550 145940 685790
rect 146180 685550 146290 685790
rect 146530 685550 146620 685790
rect 146860 685550 146950 685790
rect 147190 685550 147280 685790
rect 147520 685550 147630 685790
rect 147870 685550 147960 685790
rect 148200 685550 148290 685790
rect 148530 685550 148620 685790
rect 148860 685550 148970 685790
rect 149210 685550 149300 685790
rect 149540 685550 149630 685790
rect 149870 685550 149960 685790
rect 150200 685550 150310 685790
rect 150550 685550 150640 685790
rect 150880 685550 150970 685790
rect 151210 685550 151300 685790
rect 151540 685550 151650 685790
rect 151890 685550 151980 685790
rect 152220 685550 152310 685790
rect 152550 685550 152640 685790
rect 152880 685550 152990 685790
rect 153230 685550 153320 685790
rect 153560 685550 153650 685790
rect 153890 685550 153980 685790
rect 154220 685550 154330 685790
rect 154570 685550 154660 685790
rect 154900 685550 154990 685790
rect 155230 685550 155320 685790
rect 155560 685550 155670 685790
rect 155910 685550 155960 685790
rect 110760 685460 155960 685550
rect 110760 685220 110810 685460
rect 111050 685220 111140 685460
rect 111380 685220 111470 685460
rect 111710 685220 111800 685460
rect 112040 685220 112150 685460
rect 112390 685220 112480 685460
rect 112720 685220 112810 685460
rect 113050 685220 113140 685460
rect 113380 685220 113490 685460
rect 113730 685220 113820 685460
rect 114060 685220 114150 685460
rect 114390 685220 114480 685460
rect 114720 685220 114830 685460
rect 115070 685220 115160 685460
rect 115400 685220 115490 685460
rect 115730 685220 115820 685460
rect 116060 685220 116170 685460
rect 116410 685220 116500 685460
rect 116740 685220 116830 685460
rect 117070 685220 117160 685460
rect 117400 685220 117510 685460
rect 117750 685220 117840 685460
rect 118080 685220 118170 685460
rect 118410 685220 118500 685460
rect 118740 685220 118850 685460
rect 119090 685220 119180 685460
rect 119420 685220 119510 685460
rect 119750 685220 119840 685460
rect 120080 685220 120190 685460
rect 120430 685220 120520 685460
rect 120760 685220 120850 685460
rect 121090 685220 121180 685460
rect 121420 685220 121530 685460
rect 121770 685220 122190 685460
rect 122430 685220 122520 685460
rect 122760 685220 122850 685460
rect 123090 685220 123180 685460
rect 123420 685220 123530 685460
rect 123770 685220 123860 685460
rect 124100 685220 124190 685460
rect 124430 685220 124520 685460
rect 124760 685220 124870 685460
rect 125110 685220 125200 685460
rect 125440 685220 125530 685460
rect 125770 685220 125860 685460
rect 126100 685220 126210 685460
rect 126450 685220 126540 685460
rect 126780 685220 126870 685460
rect 127110 685220 127200 685460
rect 127440 685220 127550 685460
rect 127790 685220 127880 685460
rect 128120 685220 128210 685460
rect 128450 685220 128540 685460
rect 128780 685220 128890 685460
rect 129130 685220 129220 685460
rect 129460 685220 129550 685460
rect 129790 685220 129880 685460
rect 130120 685220 130230 685460
rect 130470 685220 130560 685460
rect 130800 685220 130890 685460
rect 131130 685220 131220 685460
rect 131460 685220 131570 685460
rect 131810 685220 131900 685460
rect 132140 685220 132230 685460
rect 132470 685220 132560 685460
rect 132800 685220 132910 685460
rect 133150 685220 133570 685460
rect 133810 685220 133900 685460
rect 134140 685220 134230 685460
rect 134470 685220 134560 685460
rect 134800 685220 134910 685460
rect 135150 685220 135240 685460
rect 135480 685220 135570 685460
rect 135810 685220 135900 685460
rect 136140 685220 136250 685460
rect 136490 685220 136580 685460
rect 136820 685220 136910 685460
rect 137150 685220 137240 685460
rect 137480 685220 137590 685460
rect 137830 685220 137920 685460
rect 138160 685220 138250 685460
rect 138490 685220 138580 685460
rect 138820 685220 138930 685460
rect 139170 685220 139260 685460
rect 139500 685220 139590 685460
rect 139830 685220 139920 685460
rect 140160 685220 140270 685460
rect 140510 685220 140600 685460
rect 140840 685220 140930 685460
rect 141170 685220 141260 685460
rect 141500 685220 141610 685460
rect 141850 685220 141940 685460
rect 142180 685220 142270 685460
rect 142510 685220 142600 685460
rect 142840 685220 142950 685460
rect 143190 685220 143280 685460
rect 143520 685220 143610 685460
rect 143850 685220 143940 685460
rect 144180 685220 144290 685460
rect 144530 685220 144950 685460
rect 145190 685220 145280 685460
rect 145520 685220 145610 685460
rect 145850 685220 145940 685460
rect 146180 685220 146290 685460
rect 146530 685220 146620 685460
rect 146860 685220 146950 685460
rect 147190 685220 147280 685460
rect 147520 685220 147630 685460
rect 147870 685220 147960 685460
rect 148200 685220 148290 685460
rect 148530 685220 148620 685460
rect 148860 685220 148970 685460
rect 149210 685220 149300 685460
rect 149540 685220 149630 685460
rect 149870 685220 149960 685460
rect 150200 685220 150310 685460
rect 150550 685220 150640 685460
rect 150880 685220 150970 685460
rect 151210 685220 151300 685460
rect 151540 685220 151650 685460
rect 151890 685220 151980 685460
rect 152220 685220 152310 685460
rect 152550 685220 152640 685460
rect 152880 685220 152990 685460
rect 153230 685220 153320 685460
rect 153560 685220 153650 685460
rect 153890 685220 153980 685460
rect 154220 685220 154330 685460
rect 154570 685220 154660 685460
rect 154900 685220 154990 685460
rect 155230 685220 155320 685460
rect 155560 685220 155670 685460
rect 155910 685220 155960 685460
rect 110760 685110 155960 685220
rect 110760 684870 110810 685110
rect 111050 684870 111140 685110
rect 111380 684870 111470 685110
rect 111710 684870 111800 685110
rect 112040 684870 112150 685110
rect 112390 684870 112480 685110
rect 112720 684870 112810 685110
rect 113050 684870 113140 685110
rect 113380 684870 113490 685110
rect 113730 684870 113820 685110
rect 114060 684870 114150 685110
rect 114390 684870 114480 685110
rect 114720 684870 114830 685110
rect 115070 684870 115160 685110
rect 115400 684870 115490 685110
rect 115730 684870 115820 685110
rect 116060 684870 116170 685110
rect 116410 684870 116500 685110
rect 116740 684870 116830 685110
rect 117070 684870 117160 685110
rect 117400 684870 117510 685110
rect 117750 684870 117840 685110
rect 118080 684870 118170 685110
rect 118410 684870 118500 685110
rect 118740 684870 118850 685110
rect 119090 684870 119180 685110
rect 119420 684870 119510 685110
rect 119750 684870 119840 685110
rect 120080 684870 120190 685110
rect 120430 684870 120520 685110
rect 120760 684870 120850 685110
rect 121090 684870 121180 685110
rect 121420 684870 121530 685110
rect 121770 684870 122190 685110
rect 122430 684870 122520 685110
rect 122760 684870 122850 685110
rect 123090 684870 123180 685110
rect 123420 684870 123530 685110
rect 123770 684870 123860 685110
rect 124100 684870 124190 685110
rect 124430 684870 124520 685110
rect 124760 684870 124870 685110
rect 125110 684870 125200 685110
rect 125440 684870 125530 685110
rect 125770 684870 125860 685110
rect 126100 684870 126210 685110
rect 126450 684870 126540 685110
rect 126780 684870 126870 685110
rect 127110 684870 127200 685110
rect 127440 684870 127550 685110
rect 127790 684870 127880 685110
rect 128120 684870 128210 685110
rect 128450 684870 128540 685110
rect 128780 684870 128890 685110
rect 129130 684870 129220 685110
rect 129460 684870 129550 685110
rect 129790 684870 129880 685110
rect 130120 684870 130230 685110
rect 130470 684870 130560 685110
rect 130800 684870 130890 685110
rect 131130 684870 131220 685110
rect 131460 684870 131570 685110
rect 131810 684870 131900 685110
rect 132140 684870 132230 685110
rect 132470 684870 132560 685110
rect 132800 684870 132910 685110
rect 133150 684870 133570 685110
rect 133810 684870 133900 685110
rect 134140 684870 134230 685110
rect 134470 684870 134560 685110
rect 134800 684870 134910 685110
rect 135150 684870 135240 685110
rect 135480 684870 135570 685110
rect 135810 684870 135900 685110
rect 136140 684870 136250 685110
rect 136490 684870 136580 685110
rect 136820 684870 136910 685110
rect 137150 684870 137240 685110
rect 137480 684870 137590 685110
rect 137830 684870 137920 685110
rect 138160 684870 138250 685110
rect 138490 684870 138580 685110
rect 138820 684870 138930 685110
rect 139170 684870 139260 685110
rect 139500 684870 139590 685110
rect 139830 684870 139920 685110
rect 140160 684870 140270 685110
rect 140510 684870 140600 685110
rect 140840 684870 140930 685110
rect 141170 684870 141260 685110
rect 141500 684870 141610 685110
rect 141850 684870 141940 685110
rect 142180 684870 142270 685110
rect 142510 684870 142600 685110
rect 142840 684870 142950 685110
rect 143190 684870 143280 685110
rect 143520 684870 143610 685110
rect 143850 684870 143940 685110
rect 144180 684870 144290 685110
rect 144530 684870 144950 685110
rect 145190 684870 145280 685110
rect 145520 684870 145610 685110
rect 145850 684870 145940 685110
rect 146180 684870 146290 685110
rect 146530 684870 146620 685110
rect 146860 684870 146950 685110
rect 147190 684870 147280 685110
rect 147520 684870 147630 685110
rect 147870 684870 147960 685110
rect 148200 684870 148290 685110
rect 148530 684870 148620 685110
rect 148860 684870 148970 685110
rect 149210 684870 149300 685110
rect 149540 684870 149630 685110
rect 149870 684870 149960 685110
rect 150200 684870 150310 685110
rect 150550 684870 150640 685110
rect 150880 684870 150970 685110
rect 151210 684870 151300 685110
rect 151540 684870 151650 685110
rect 151890 684870 151980 685110
rect 152220 684870 152310 685110
rect 152550 684870 152640 685110
rect 152880 684870 152990 685110
rect 153230 684870 153320 685110
rect 153560 684870 153650 685110
rect 153890 684870 153980 685110
rect 154220 684870 154330 685110
rect 154570 684870 154660 685110
rect 154900 684870 154990 685110
rect 155230 684870 155320 685110
rect 155560 684870 155670 685110
rect 155910 684870 155960 685110
rect 110760 684780 155960 684870
rect 110760 684540 110810 684780
rect 111050 684540 111140 684780
rect 111380 684540 111470 684780
rect 111710 684540 111800 684780
rect 112040 684540 112150 684780
rect 112390 684540 112480 684780
rect 112720 684540 112810 684780
rect 113050 684540 113140 684780
rect 113380 684540 113490 684780
rect 113730 684540 113820 684780
rect 114060 684540 114150 684780
rect 114390 684540 114480 684780
rect 114720 684540 114830 684780
rect 115070 684540 115160 684780
rect 115400 684540 115490 684780
rect 115730 684540 115820 684780
rect 116060 684540 116170 684780
rect 116410 684540 116500 684780
rect 116740 684540 116830 684780
rect 117070 684540 117160 684780
rect 117400 684540 117510 684780
rect 117750 684540 117840 684780
rect 118080 684540 118170 684780
rect 118410 684540 118500 684780
rect 118740 684540 118850 684780
rect 119090 684540 119180 684780
rect 119420 684540 119510 684780
rect 119750 684540 119840 684780
rect 120080 684540 120190 684780
rect 120430 684540 120520 684780
rect 120760 684540 120850 684780
rect 121090 684540 121180 684780
rect 121420 684540 121530 684780
rect 121770 684540 122190 684780
rect 122430 684540 122520 684780
rect 122760 684540 122850 684780
rect 123090 684540 123180 684780
rect 123420 684540 123530 684780
rect 123770 684540 123860 684780
rect 124100 684540 124190 684780
rect 124430 684540 124520 684780
rect 124760 684540 124870 684780
rect 125110 684540 125200 684780
rect 125440 684540 125530 684780
rect 125770 684540 125860 684780
rect 126100 684540 126210 684780
rect 126450 684540 126540 684780
rect 126780 684540 126870 684780
rect 127110 684540 127200 684780
rect 127440 684540 127550 684780
rect 127790 684540 127880 684780
rect 128120 684540 128210 684780
rect 128450 684540 128540 684780
rect 128780 684540 128890 684780
rect 129130 684540 129220 684780
rect 129460 684540 129550 684780
rect 129790 684540 129880 684780
rect 130120 684540 130230 684780
rect 130470 684540 130560 684780
rect 130800 684540 130890 684780
rect 131130 684540 131220 684780
rect 131460 684540 131570 684780
rect 131810 684540 131900 684780
rect 132140 684540 132230 684780
rect 132470 684540 132560 684780
rect 132800 684540 132910 684780
rect 133150 684540 133570 684780
rect 133810 684540 133900 684780
rect 134140 684540 134230 684780
rect 134470 684540 134560 684780
rect 134800 684540 134910 684780
rect 135150 684540 135240 684780
rect 135480 684540 135570 684780
rect 135810 684540 135900 684780
rect 136140 684540 136250 684780
rect 136490 684540 136580 684780
rect 136820 684540 136910 684780
rect 137150 684540 137240 684780
rect 137480 684540 137590 684780
rect 137830 684540 137920 684780
rect 138160 684540 138250 684780
rect 138490 684540 138580 684780
rect 138820 684540 138930 684780
rect 139170 684540 139260 684780
rect 139500 684540 139590 684780
rect 139830 684540 139920 684780
rect 140160 684540 140270 684780
rect 140510 684540 140600 684780
rect 140840 684540 140930 684780
rect 141170 684540 141260 684780
rect 141500 684540 141610 684780
rect 141850 684540 141940 684780
rect 142180 684540 142270 684780
rect 142510 684540 142600 684780
rect 142840 684540 142950 684780
rect 143190 684540 143280 684780
rect 143520 684540 143610 684780
rect 143850 684540 143940 684780
rect 144180 684540 144290 684780
rect 144530 684540 144950 684780
rect 145190 684540 145280 684780
rect 145520 684540 145610 684780
rect 145850 684540 145940 684780
rect 146180 684540 146290 684780
rect 146530 684540 146620 684780
rect 146860 684540 146950 684780
rect 147190 684540 147280 684780
rect 147520 684540 147630 684780
rect 147870 684540 147960 684780
rect 148200 684540 148290 684780
rect 148530 684540 148620 684780
rect 148860 684540 148970 684780
rect 149210 684540 149300 684780
rect 149540 684540 149630 684780
rect 149870 684540 149960 684780
rect 150200 684540 150310 684780
rect 150550 684540 150640 684780
rect 150880 684540 150970 684780
rect 151210 684540 151300 684780
rect 151540 684540 151650 684780
rect 151890 684540 151980 684780
rect 152220 684540 152310 684780
rect 152550 684540 152640 684780
rect 152880 684540 152990 684780
rect 153230 684540 153320 684780
rect 153560 684540 153650 684780
rect 153890 684540 153980 684780
rect 154220 684540 154330 684780
rect 154570 684540 154660 684780
rect 154900 684540 154990 684780
rect 155230 684540 155320 684780
rect 155560 684540 155670 684780
rect 155910 684540 155960 684780
rect 110760 684450 155960 684540
rect 110760 684210 110810 684450
rect 111050 684210 111140 684450
rect 111380 684210 111470 684450
rect 111710 684210 111800 684450
rect 112040 684210 112150 684450
rect 112390 684210 112480 684450
rect 112720 684210 112810 684450
rect 113050 684210 113140 684450
rect 113380 684210 113490 684450
rect 113730 684210 113820 684450
rect 114060 684210 114150 684450
rect 114390 684210 114480 684450
rect 114720 684210 114830 684450
rect 115070 684210 115160 684450
rect 115400 684210 115490 684450
rect 115730 684210 115820 684450
rect 116060 684210 116170 684450
rect 116410 684210 116500 684450
rect 116740 684210 116830 684450
rect 117070 684210 117160 684450
rect 117400 684210 117510 684450
rect 117750 684210 117840 684450
rect 118080 684210 118170 684450
rect 118410 684210 118500 684450
rect 118740 684210 118850 684450
rect 119090 684210 119180 684450
rect 119420 684210 119510 684450
rect 119750 684210 119840 684450
rect 120080 684210 120190 684450
rect 120430 684210 120520 684450
rect 120760 684210 120850 684450
rect 121090 684210 121180 684450
rect 121420 684210 121530 684450
rect 121770 684210 122190 684450
rect 122430 684210 122520 684450
rect 122760 684210 122850 684450
rect 123090 684210 123180 684450
rect 123420 684210 123530 684450
rect 123770 684210 123860 684450
rect 124100 684210 124190 684450
rect 124430 684210 124520 684450
rect 124760 684210 124870 684450
rect 125110 684210 125200 684450
rect 125440 684210 125530 684450
rect 125770 684210 125860 684450
rect 126100 684210 126210 684450
rect 126450 684210 126540 684450
rect 126780 684210 126870 684450
rect 127110 684210 127200 684450
rect 127440 684210 127550 684450
rect 127790 684210 127880 684450
rect 128120 684210 128210 684450
rect 128450 684210 128540 684450
rect 128780 684210 128890 684450
rect 129130 684210 129220 684450
rect 129460 684210 129550 684450
rect 129790 684210 129880 684450
rect 130120 684210 130230 684450
rect 130470 684210 130560 684450
rect 130800 684210 130890 684450
rect 131130 684210 131220 684450
rect 131460 684210 131570 684450
rect 131810 684210 131900 684450
rect 132140 684210 132230 684450
rect 132470 684210 132560 684450
rect 132800 684210 132910 684450
rect 133150 684210 133570 684450
rect 133810 684210 133900 684450
rect 134140 684210 134230 684450
rect 134470 684210 134560 684450
rect 134800 684210 134910 684450
rect 135150 684210 135240 684450
rect 135480 684210 135570 684450
rect 135810 684210 135900 684450
rect 136140 684210 136250 684450
rect 136490 684210 136580 684450
rect 136820 684210 136910 684450
rect 137150 684210 137240 684450
rect 137480 684210 137590 684450
rect 137830 684210 137920 684450
rect 138160 684210 138250 684450
rect 138490 684210 138580 684450
rect 138820 684210 138930 684450
rect 139170 684210 139260 684450
rect 139500 684210 139590 684450
rect 139830 684210 139920 684450
rect 140160 684210 140270 684450
rect 140510 684210 140600 684450
rect 140840 684210 140930 684450
rect 141170 684210 141260 684450
rect 141500 684210 141610 684450
rect 141850 684210 141940 684450
rect 142180 684210 142270 684450
rect 142510 684210 142600 684450
rect 142840 684210 142950 684450
rect 143190 684210 143280 684450
rect 143520 684210 143610 684450
rect 143850 684210 143940 684450
rect 144180 684210 144290 684450
rect 144530 684210 144950 684450
rect 145190 684210 145280 684450
rect 145520 684210 145610 684450
rect 145850 684210 145940 684450
rect 146180 684210 146290 684450
rect 146530 684210 146620 684450
rect 146860 684210 146950 684450
rect 147190 684210 147280 684450
rect 147520 684210 147630 684450
rect 147870 684210 147960 684450
rect 148200 684210 148290 684450
rect 148530 684210 148620 684450
rect 148860 684210 148970 684450
rect 149210 684210 149300 684450
rect 149540 684210 149630 684450
rect 149870 684210 149960 684450
rect 150200 684210 150310 684450
rect 150550 684210 150640 684450
rect 150880 684210 150970 684450
rect 151210 684210 151300 684450
rect 151540 684210 151650 684450
rect 151890 684210 151980 684450
rect 152220 684210 152310 684450
rect 152550 684210 152640 684450
rect 152880 684210 152990 684450
rect 153230 684210 153320 684450
rect 153560 684210 153650 684450
rect 153890 684210 153980 684450
rect 154220 684210 154330 684450
rect 154570 684210 154660 684450
rect 154900 684210 154990 684450
rect 155230 684210 155320 684450
rect 155560 684210 155670 684450
rect 155910 684210 155960 684450
rect 110760 684120 155960 684210
rect 110760 683880 110810 684120
rect 111050 683880 111140 684120
rect 111380 683880 111470 684120
rect 111710 683880 111800 684120
rect 112040 683880 112150 684120
rect 112390 683880 112480 684120
rect 112720 683880 112810 684120
rect 113050 683880 113140 684120
rect 113380 683880 113490 684120
rect 113730 683880 113820 684120
rect 114060 683880 114150 684120
rect 114390 683880 114480 684120
rect 114720 683880 114830 684120
rect 115070 683880 115160 684120
rect 115400 683880 115490 684120
rect 115730 683880 115820 684120
rect 116060 683880 116170 684120
rect 116410 683880 116500 684120
rect 116740 683880 116830 684120
rect 117070 683880 117160 684120
rect 117400 683880 117510 684120
rect 117750 683880 117840 684120
rect 118080 683880 118170 684120
rect 118410 683880 118500 684120
rect 118740 683880 118850 684120
rect 119090 683880 119180 684120
rect 119420 683880 119510 684120
rect 119750 683880 119840 684120
rect 120080 683880 120190 684120
rect 120430 683880 120520 684120
rect 120760 683880 120850 684120
rect 121090 683880 121180 684120
rect 121420 683880 121530 684120
rect 121770 683880 122190 684120
rect 122430 683880 122520 684120
rect 122760 683880 122850 684120
rect 123090 683880 123180 684120
rect 123420 683880 123530 684120
rect 123770 683880 123860 684120
rect 124100 683880 124190 684120
rect 124430 683880 124520 684120
rect 124760 683880 124870 684120
rect 125110 683880 125200 684120
rect 125440 683880 125530 684120
rect 125770 683880 125860 684120
rect 126100 683880 126210 684120
rect 126450 683880 126540 684120
rect 126780 683880 126870 684120
rect 127110 683880 127200 684120
rect 127440 683880 127550 684120
rect 127790 683880 127880 684120
rect 128120 683880 128210 684120
rect 128450 683880 128540 684120
rect 128780 683880 128890 684120
rect 129130 683880 129220 684120
rect 129460 683880 129550 684120
rect 129790 683880 129880 684120
rect 130120 683880 130230 684120
rect 130470 683880 130560 684120
rect 130800 683880 130890 684120
rect 131130 683880 131220 684120
rect 131460 683880 131570 684120
rect 131810 683880 131900 684120
rect 132140 683880 132230 684120
rect 132470 683880 132560 684120
rect 132800 683880 132910 684120
rect 133150 683880 133570 684120
rect 133810 683880 133900 684120
rect 134140 683880 134230 684120
rect 134470 683880 134560 684120
rect 134800 683880 134910 684120
rect 135150 683880 135240 684120
rect 135480 683880 135570 684120
rect 135810 683880 135900 684120
rect 136140 683880 136250 684120
rect 136490 683880 136580 684120
rect 136820 683880 136910 684120
rect 137150 683880 137240 684120
rect 137480 683880 137590 684120
rect 137830 683880 137920 684120
rect 138160 683880 138250 684120
rect 138490 683880 138580 684120
rect 138820 683880 138930 684120
rect 139170 683880 139260 684120
rect 139500 683880 139590 684120
rect 139830 683880 139920 684120
rect 140160 683880 140270 684120
rect 140510 683880 140600 684120
rect 140840 683880 140930 684120
rect 141170 683880 141260 684120
rect 141500 683880 141610 684120
rect 141850 683880 141940 684120
rect 142180 683880 142270 684120
rect 142510 683880 142600 684120
rect 142840 683880 142950 684120
rect 143190 683880 143280 684120
rect 143520 683880 143610 684120
rect 143850 683880 143940 684120
rect 144180 683880 144290 684120
rect 144530 683880 144950 684120
rect 145190 683880 145280 684120
rect 145520 683880 145610 684120
rect 145850 683880 145940 684120
rect 146180 683880 146290 684120
rect 146530 683880 146620 684120
rect 146860 683880 146950 684120
rect 147190 683880 147280 684120
rect 147520 683880 147630 684120
rect 147870 683880 147960 684120
rect 148200 683880 148290 684120
rect 148530 683880 148620 684120
rect 148860 683880 148970 684120
rect 149210 683880 149300 684120
rect 149540 683880 149630 684120
rect 149870 683880 149960 684120
rect 150200 683880 150310 684120
rect 150550 683880 150640 684120
rect 150880 683880 150970 684120
rect 151210 683880 151300 684120
rect 151540 683880 151650 684120
rect 151890 683880 151980 684120
rect 152220 683880 152310 684120
rect 152550 683880 152640 684120
rect 152880 683880 152990 684120
rect 153230 683880 153320 684120
rect 153560 683880 153650 684120
rect 153890 683880 153980 684120
rect 154220 683880 154330 684120
rect 154570 683880 154660 684120
rect 154900 683880 154990 684120
rect 155230 683880 155320 684120
rect 155560 683880 155670 684120
rect 155910 683880 155960 684120
rect 110760 683830 155960 683880
rect 121820 683730 122140 683740
rect 133200 683730 133520 683740
rect 144580 683730 144900 683740
rect 110760 683700 155960 683730
rect 110760 683460 110890 683700
rect 111130 683460 111220 683700
rect 111460 683460 111550 683700
rect 111790 683460 111880 683700
rect 112120 683460 112210 683700
rect 112450 683460 112540 683700
rect 112780 683460 112870 683700
rect 113110 683460 113200 683700
rect 113440 683460 113530 683700
rect 113770 683460 113860 683700
rect 114100 683460 114190 683700
rect 114430 683460 114520 683700
rect 114760 683460 114850 683700
rect 115090 683460 115180 683700
rect 115420 683460 115510 683700
rect 115750 683460 115840 683700
rect 116080 683460 116170 683700
rect 116410 683460 116500 683700
rect 116740 683460 116830 683700
rect 117070 683460 117160 683700
rect 117400 683460 117490 683700
rect 117730 683460 117820 683700
rect 118060 683460 118150 683700
rect 118390 683460 118480 683700
rect 118720 683460 118810 683700
rect 119050 683460 119140 683700
rect 119380 683460 119470 683700
rect 119710 683460 119800 683700
rect 120040 683460 120130 683700
rect 120370 683460 120460 683700
rect 120700 683460 120790 683700
rect 121030 683460 121120 683700
rect 121360 683460 121450 683700
rect 121690 683460 122270 683700
rect 122510 683460 122600 683700
rect 122840 683460 122930 683700
rect 123170 683460 123260 683700
rect 123500 683460 123590 683700
rect 123830 683460 123920 683700
rect 124160 683460 124250 683700
rect 124490 683460 124580 683700
rect 124820 683460 124910 683700
rect 125150 683460 125240 683700
rect 125480 683460 125570 683700
rect 125810 683460 125900 683700
rect 126140 683460 126230 683700
rect 126470 683460 126560 683700
rect 126800 683460 126890 683700
rect 127130 683460 127220 683700
rect 127460 683460 127550 683700
rect 127790 683460 127880 683700
rect 128120 683460 128210 683700
rect 128450 683460 128540 683700
rect 128780 683460 128870 683700
rect 129110 683460 129200 683700
rect 129440 683460 129530 683700
rect 129770 683460 129860 683700
rect 130100 683460 130190 683700
rect 130430 683460 130520 683700
rect 130760 683460 130850 683700
rect 131090 683460 131180 683700
rect 131420 683460 131510 683700
rect 131750 683460 131840 683700
rect 132080 683460 132170 683700
rect 132410 683460 132500 683700
rect 132740 683460 132830 683700
rect 133070 683460 133650 683700
rect 133890 683460 133980 683700
rect 134220 683460 134310 683700
rect 134550 683460 134640 683700
rect 134880 683460 134970 683700
rect 135210 683460 135300 683700
rect 135540 683460 135630 683700
rect 135870 683460 135960 683700
rect 136200 683460 136290 683700
rect 136530 683460 136620 683700
rect 136860 683460 136950 683700
rect 137190 683460 137280 683700
rect 137520 683460 137610 683700
rect 137850 683460 137940 683700
rect 138180 683460 138270 683700
rect 138510 683460 138600 683700
rect 138840 683460 138930 683700
rect 139170 683460 139260 683700
rect 139500 683460 139590 683700
rect 139830 683460 139920 683700
rect 140160 683460 140250 683700
rect 140490 683460 140580 683700
rect 140820 683460 140910 683700
rect 141150 683460 141240 683700
rect 141480 683460 141570 683700
rect 141810 683460 141900 683700
rect 142140 683460 142230 683700
rect 142470 683460 142560 683700
rect 142800 683460 142890 683700
rect 143130 683460 143220 683700
rect 143460 683460 143550 683700
rect 143790 683460 143880 683700
rect 144120 683460 144210 683700
rect 144450 683460 145030 683700
rect 145270 683460 145360 683700
rect 145600 683460 145690 683700
rect 145930 683460 146020 683700
rect 146260 683460 146350 683700
rect 146590 683460 146680 683700
rect 146920 683460 147010 683700
rect 147250 683460 147340 683700
rect 147580 683460 147670 683700
rect 147910 683460 148000 683700
rect 148240 683460 148330 683700
rect 148570 683460 148660 683700
rect 148900 683460 148990 683700
rect 149230 683460 149320 683700
rect 149560 683460 149650 683700
rect 149890 683460 149980 683700
rect 150220 683460 150310 683700
rect 150550 683460 150640 683700
rect 150880 683460 150970 683700
rect 151210 683460 151300 683700
rect 151540 683460 151630 683700
rect 151870 683460 151960 683700
rect 152200 683460 152290 683700
rect 152530 683460 152620 683700
rect 152860 683460 152950 683700
rect 153190 683460 153280 683700
rect 153520 683460 153610 683700
rect 153850 683460 153940 683700
rect 154180 683460 154270 683700
rect 154510 683460 154600 683700
rect 154840 683460 154930 683700
rect 155170 683460 155260 683700
rect 155500 683460 155590 683700
rect 155830 683460 155960 683700
rect 110760 683430 155960 683460
rect 121820 683420 122140 683430
rect 133200 683420 133520 683430
rect 144580 683420 144900 683430
rect 110760 683280 155960 683330
rect 110760 683040 110810 683280
rect 111050 683040 111160 683280
rect 111400 683040 111490 683280
rect 111730 683040 111820 683280
rect 112060 683040 112150 683280
rect 112390 683040 112500 683280
rect 112740 683040 112830 683280
rect 113070 683040 113160 683280
rect 113400 683040 113490 683280
rect 113730 683040 113840 683280
rect 114080 683040 114170 683280
rect 114410 683040 114500 683280
rect 114740 683040 114830 683280
rect 115070 683040 115180 683280
rect 115420 683040 115510 683280
rect 115750 683040 115840 683280
rect 116080 683040 116170 683280
rect 116410 683040 116520 683280
rect 116760 683040 116850 683280
rect 117090 683040 117180 683280
rect 117420 683040 117510 683280
rect 117750 683040 117860 683280
rect 118100 683040 118190 683280
rect 118430 683040 118520 683280
rect 118760 683040 118850 683280
rect 119090 683040 119200 683280
rect 119440 683040 119530 683280
rect 119770 683040 119860 683280
rect 120100 683040 120190 683280
rect 120430 683040 120540 683280
rect 120780 683040 120870 683280
rect 121110 683040 121200 683280
rect 121440 683040 121530 683280
rect 121770 683040 122190 683280
rect 122430 683040 122540 683280
rect 122780 683040 122870 683280
rect 123110 683040 123200 683280
rect 123440 683040 123530 683280
rect 123770 683040 123880 683280
rect 124120 683040 124210 683280
rect 124450 683040 124540 683280
rect 124780 683040 124870 683280
rect 125110 683040 125220 683280
rect 125460 683040 125550 683280
rect 125790 683040 125880 683280
rect 126120 683040 126210 683280
rect 126450 683040 126560 683280
rect 126800 683040 126890 683280
rect 127130 683040 127220 683280
rect 127460 683040 127550 683280
rect 127790 683040 127900 683280
rect 128140 683040 128230 683280
rect 128470 683040 128560 683280
rect 128800 683040 128890 683280
rect 129130 683040 129240 683280
rect 129480 683040 129570 683280
rect 129810 683040 129900 683280
rect 130140 683040 130230 683280
rect 130470 683040 130580 683280
rect 130820 683040 130910 683280
rect 131150 683040 131240 683280
rect 131480 683040 131570 683280
rect 131810 683040 131920 683280
rect 132160 683040 132250 683280
rect 132490 683040 132580 683280
rect 132820 683040 132910 683280
rect 133150 683040 133570 683280
rect 133810 683040 133920 683280
rect 134160 683040 134250 683280
rect 134490 683040 134580 683280
rect 134820 683040 134910 683280
rect 135150 683040 135260 683280
rect 135500 683040 135590 683280
rect 135830 683040 135920 683280
rect 136160 683040 136250 683280
rect 136490 683040 136600 683280
rect 136840 683040 136930 683280
rect 137170 683040 137260 683280
rect 137500 683040 137590 683280
rect 137830 683040 137940 683280
rect 138180 683040 138270 683280
rect 138510 683040 138600 683280
rect 138840 683040 138930 683280
rect 139170 683040 139280 683280
rect 139520 683040 139610 683280
rect 139850 683040 139940 683280
rect 140180 683040 140270 683280
rect 140510 683040 140620 683280
rect 140860 683040 140950 683280
rect 141190 683040 141280 683280
rect 141520 683040 141610 683280
rect 141850 683040 141960 683280
rect 142200 683040 142290 683280
rect 142530 683040 142620 683280
rect 142860 683040 142950 683280
rect 143190 683040 143300 683280
rect 143540 683040 143630 683280
rect 143870 683040 143960 683280
rect 144200 683040 144290 683280
rect 144530 683040 144950 683280
rect 145190 683040 145300 683280
rect 145540 683040 145630 683280
rect 145870 683040 145960 683280
rect 146200 683040 146290 683280
rect 146530 683040 146640 683280
rect 146880 683040 146970 683280
rect 147210 683040 147300 683280
rect 147540 683040 147630 683280
rect 147870 683040 147980 683280
rect 148220 683040 148310 683280
rect 148550 683040 148640 683280
rect 148880 683040 148970 683280
rect 149210 683040 149320 683280
rect 149560 683040 149650 683280
rect 149890 683040 149980 683280
rect 150220 683040 150310 683280
rect 150550 683040 150660 683280
rect 150900 683040 150990 683280
rect 151230 683040 151320 683280
rect 151560 683040 151650 683280
rect 151890 683040 152000 683280
rect 152240 683040 152330 683280
rect 152570 683040 152660 683280
rect 152900 683040 152990 683280
rect 153230 683040 153340 683280
rect 153580 683040 153670 683280
rect 153910 683040 154000 683280
rect 154240 683040 154330 683280
rect 154570 683040 154680 683280
rect 154920 683040 155010 683280
rect 155250 683040 155340 683280
rect 155580 683040 155670 683280
rect 155910 683040 155960 683280
rect 110760 682950 155960 683040
rect 110760 682710 110810 682950
rect 111050 682710 111160 682950
rect 111400 682710 111490 682950
rect 111730 682710 111820 682950
rect 112060 682710 112150 682950
rect 112390 682710 112500 682950
rect 112740 682710 112830 682950
rect 113070 682710 113160 682950
rect 113400 682710 113490 682950
rect 113730 682710 113840 682950
rect 114080 682710 114170 682950
rect 114410 682710 114500 682950
rect 114740 682710 114830 682950
rect 115070 682710 115180 682950
rect 115420 682710 115510 682950
rect 115750 682710 115840 682950
rect 116080 682710 116170 682950
rect 116410 682710 116520 682950
rect 116760 682710 116850 682950
rect 117090 682710 117180 682950
rect 117420 682710 117510 682950
rect 117750 682710 117860 682950
rect 118100 682710 118190 682950
rect 118430 682710 118520 682950
rect 118760 682710 118850 682950
rect 119090 682710 119200 682950
rect 119440 682710 119530 682950
rect 119770 682710 119860 682950
rect 120100 682710 120190 682950
rect 120430 682710 120540 682950
rect 120780 682710 120870 682950
rect 121110 682710 121200 682950
rect 121440 682710 121530 682950
rect 121770 682710 122190 682950
rect 122430 682710 122540 682950
rect 122780 682710 122870 682950
rect 123110 682710 123200 682950
rect 123440 682710 123530 682950
rect 123770 682710 123880 682950
rect 124120 682710 124210 682950
rect 124450 682710 124540 682950
rect 124780 682710 124870 682950
rect 125110 682710 125220 682950
rect 125460 682710 125550 682950
rect 125790 682710 125880 682950
rect 126120 682710 126210 682950
rect 126450 682710 126560 682950
rect 126800 682710 126890 682950
rect 127130 682710 127220 682950
rect 127460 682710 127550 682950
rect 127790 682710 127900 682950
rect 128140 682710 128230 682950
rect 128470 682710 128560 682950
rect 128800 682710 128890 682950
rect 129130 682710 129240 682950
rect 129480 682710 129570 682950
rect 129810 682710 129900 682950
rect 130140 682710 130230 682950
rect 130470 682710 130580 682950
rect 130820 682710 130910 682950
rect 131150 682710 131240 682950
rect 131480 682710 131570 682950
rect 131810 682710 131920 682950
rect 132160 682710 132250 682950
rect 132490 682710 132580 682950
rect 132820 682710 132910 682950
rect 133150 682710 133570 682950
rect 133810 682710 133920 682950
rect 134160 682710 134250 682950
rect 134490 682710 134580 682950
rect 134820 682710 134910 682950
rect 135150 682710 135260 682950
rect 135500 682710 135590 682950
rect 135830 682710 135920 682950
rect 136160 682710 136250 682950
rect 136490 682710 136600 682950
rect 136840 682710 136930 682950
rect 137170 682710 137260 682950
rect 137500 682710 137590 682950
rect 137830 682710 137940 682950
rect 138180 682710 138270 682950
rect 138510 682710 138600 682950
rect 138840 682710 138930 682950
rect 139170 682710 139280 682950
rect 139520 682710 139610 682950
rect 139850 682710 139940 682950
rect 140180 682710 140270 682950
rect 140510 682710 140620 682950
rect 140860 682710 140950 682950
rect 141190 682710 141280 682950
rect 141520 682710 141610 682950
rect 141850 682710 141960 682950
rect 142200 682710 142290 682950
rect 142530 682710 142620 682950
rect 142860 682710 142950 682950
rect 143190 682710 143300 682950
rect 143540 682710 143630 682950
rect 143870 682710 143960 682950
rect 144200 682710 144290 682950
rect 144530 682710 144950 682950
rect 145190 682710 145300 682950
rect 145540 682710 145630 682950
rect 145870 682710 145960 682950
rect 146200 682710 146290 682950
rect 146530 682710 146640 682950
rect 146880 682710 146970 682950
rect 147210 682710 147300 682950
rect 147540 682710 147630 682950
rect 147870 682710 147980 682950
rect 148220 682710 148310 682950
rect 148550 682710 148640 682950
rect 148880 682710 148970 682950
rect 149210 682710 149320 682950
rect 149560 682710 149650 682950
rect 149890 682710 149980 682950
rect 150220 682710 150310 682950
rect 150550 682710 150660 682950
rect 150900 682710 150990 682950
rect 151230 682710 151320 682950
rect 151560 682710 151650 682950
rect 151890 682710 152000 682950
rect 152240 682710 152330 682950
rect 152570 682710 152660 682950
rect 152900 682710 152990 682950
rect 153230 682710 153340 682950
rect 153580 682710 153670 682950
rect 153910 682710 154000 682950
rect 154240 682710 154330 682950
rect 154570 682710 154680 682950
rect 154920 682710 155010 682950
rect 155250 682710 155340 682950
rect 155580 682710 155670 682950
rect 155910 682710 155960 682950
rect 110760 682620 155960 682710
rect 110760 682380 110810 682620
rect 111050 682380 111160 682620
rect 111400 682380 111490 682620
rect 111730 682380 111820 682620
rect 112060 682380 112150 682620
rect 112390 682380 112500 682620
rect 112740 682380 112830 682620
rect 113070 682380 113160 682620
rect 113400 682380 113490 682620
rect 113730 682380 113840 682620
rect 114080 682380 114170 682620
rect 114410 682380 114500 682620
rect 114740 682380 114830 682620
rect 115070 682380 115180 682620
rect 115420 682380 115510 682620
rect 115750 682380 115840 682620
rect 116080 682380 116170 682620
rect 116410 682380 116520 682620
rect 116760 682380 116850 682620
rect 117090 682380 117180 682620
rect 117420 682380 117510 682620
rect 117750 682380 117860 682620
rect 118100 682380 118190 682620
rect 118430 682380 118520 682620
rect 118760 682380 118850 682620
rect 119090 682380 119200 682620
rect 119440 682380 119530 682620
rect 119770 682380 119860 682620
rect 120100 682380 120190 682620
rect 120430 682380 120540 682620
rect 120780 682380 120870 682620
rect 121110 682380 121200 682620
rect 121440 682380 121530 682620
rect 121770 682380 122190 682620
rect 122430 682380 122540 682620
rect 122780 682380 122870 682620
rect 123110 682380 123200 682620
rect 123440 682380 123530 682620
rect 123770 682380 123880 682620
rect 124120 682380 124210 682620
rect 124450 682380 124540 682620
rect 124780 682380 124870 682620
rect 125110 682380 125220 682620
rect 125460 682380 125550 682620
rect 125790 682380 125880 682620
rect 126120 682380 126210 682620
rect 126450 682380 126560 682620
rect 126800 682380 126890 682620
rect 127130 682380 127220 682620
rect 127460 682380 127550 682620
rect 127790 682380 127900 682620
rect 128140 682380 128230 682620
rect 128470 682380 128560 682620
rect 128800 682380 128890 682620
rect 129130 682380 129240 682620
rect 129480 682380 129570 682620
rect 129810 682380 129900 682620
rect 130140 682380 130230 682620
rect 130470 682380 130580 682620
rect 130820 682380 130910 682620
rect 131150 682380 131240 682620
rect 131480 682380 131570 682620
rect 131810 682380 131920 682620
rect 132160 682380 132250 682620
rect 132490 682380 132580 682620
rect 132820 682380 132910 682620
rect 133150 682380 133570 682620
rect 133810 682380 133920 682620
rect 134160 682380 134250 682620
rect 134490 682380 134580 682620
rect 134820 682380 134910 682620
rect 135150 682380 135260 682620
rect 135500 682380 135590 682620
rect 135830 682380 135920 682620
rect 136160 682380 136250 682620
rect 136490 682380 136600 682620
rect 136840 682380 136930 682620
rect 137170 682380 137260 682620
rect 137500 682380 137590 682620
rect 137830 682380 137940 682620
rect 138180 682380 138270 682620
rect 138510 682380 138600 682620
rect 138840 682380 138930 682620
rect 139170 682380 139280 682620
rect 139520 682380 139610 682620
rect 139850 682380 139940 682620
rect 140180 682380 140270 682620
rect 140510 682380 140620 682620
rect 140860 682380 140950 682620
rect 141190 682380 141280 682620
rect 141520 682380 141610 682620
rect 141850 682380 141960 682620
rect 142200 682380 142290 682620
rect 142530 682380 142620 682620
rect 142860 682380 142950 682620
rect 143190 682380 143300 682620
rect 143540 682380 143630 682620
rect 143870 682380 143960 682620
rect 144200 682380 144290 682620
rect 144530 682380 144950 682620
rect 145190 682380 145300 682620
rect 145540 682380 145630 682620
rect 145870 682380 145960 682620
rect 146200 682380 146290 682620
rect 146530 682380 146640 682620
rect 146880 682380 146970 682620
rect 147210 682380 147300 682620
rect 147540 682380 147630 682620
rect 147870 682380 147980 682620
rect 148220 682380 148310 682620
rect 148550 682380 148640 682620
rect 148880 682380 148970 682620
rect 149210 682380 149320 682620
rect 149560 682380 149650 682620
rect 149890 682380 149980 682620
rect 150220 682380 150310 682620
rect 150550 682380 150660 682620
rect 150900 682380 150990 682620
rect 151230 682380 151320 682620
rect 151560 682380 151650 682620
rect 151890 682380 152000 682620
rect 152240 682380 152330 682620
rect 152570 682380 152660 682620
rect 152900 682380 152990 682620
rect 153230 682380 153340 682620
rect 153580 682380 153670 682620
rect 153910 682380 154000 682620
rect 154240 682380 154330 682620
rect 154570 682380 154680 682620
rect 154920 682380 155010 682620
rect 155250 682380 155340 682620
rect 155580 682380 155670 682620
rect 155910 682380 155960 682620
rect 110760 682290 155960 682380
rect 110760 682050 110810 682290
rect 111050 682050 111160 682290
rect 111400 682050 111490 682290
rect 111730 682050 111820 682290
rect 112060 682050 112150 682290
rect 112390 682050 112500 682290
rect 112740 682050 112830 682290
rect 113070 682050 113160 682290
rect 113400 682050 113490 682290
rect 113730 682050 113840 682290
rect 114080 682050 114170 682290
rect 114410 682050 114500 682290
rect 114740 682050 114830 682290
rect 115070 682050 115180 682290
rect 115420 682050 115510 682290
rect 115750 682050 115840 682290
rect 116080 682050 116170 682290
rect 116410 682050 116520 682290
rect 116760 682050 116850 682290
rect 117090 682050 117180 682290
rect 117420 682050 117510 682290
rect 117750 682050 117860 682290
rect 118100 682050 118190 682290
rect 118430 682050 118520 682290
rect 118760 682050 118850 682290
rect 119090 682050 119200 682290
rect 119440 682050 119530 682290
rect 119770 682050 119860 682290
rect 120100 682050 120190 682290
rect 120430 682050 120540 682290
rect 120780 682050 120870 682290
rect 121110 682050 121200 682290
rect 121440 682050 121530 682290
rect 121770 682050 122190 682290
rect 122430 682050 122540 682290
rect 122780 682050 122870 682290
rect 123110 682050 123200 682290
rect 123440 682050 123530 682290
rect 123770 682050 123880 682290
rect 124120 682050 124210 682290
rect 124450 682050 124540 682290
rect 124780 682050 124870 682290
rect 125110 682050 125220 682290
rect 125460 682050 125550 682290
rect 125790 682050 125880 682290
rect 126120 682050 126210 682290
rect 126450 682050 126560 682290
rect 126800 682050 126890 682290
rect 127130 682050 127220 682290
rect 127460 682050 127550 682290
rect 127790 682050 127900 682290
rect 128140 682050 128230 682290
rect 128470 682050 128560 682290
rect 128800 682050 128890 682290
rect 129130 682050 129240 682290
rect 129480 682050 129570 682290
rect 129810 682050 129900 682290
rect 130140 682050 130230 682290
rect 130470 682050 130580 682290
rect 130820 682050 130910 682290
rect 131150 682050 131240 682290
rect 131480 682050 131570 682290
rect 131810 682050 131920 682290
rect 132160 682050 132250 682290
rect 132490 682050 132580 682290
rect 132820 682050 132910 682290
rect 133150 682050 133570 682290
rect 133810 682050 133920 682290
rect 134160 682050 134250 682290
rect 134490 682050 134580 682290
rect 134820 682050 134910 682290
rect 135150 682050 135260 682290
rect 135500 682050 135590 682290
rect 135830 682050 135920 682290
rect 136160 682050 136250 682290
rect 136490 682050 136600 682290
rect 136840 682050 136930 682290
rect 137170 682050 137260 682290
rect 137500 682050 137590 682290
rect 137830 682050 137940 682290
rect 138180 682050 138270 682290
rect 138510 682050 138600 682290
rect 138840 682050 138930 682290
rect 139170 682050 139280 682290
rect 139520 682050 139610 682290
rect 139850 682050 139940 682290
rect 140180 682050 140270 682290
rect 140510 682050 140620 682290
rect 140860 682050 140950 682290
rect 141190 682050 141280 682290
rect 141520 682050 141610 682290
rect 141850 682050 141960 682290
rect 142200 682050 142290 682290
rect 142530 682050 142620 682290
rect 142860 682050 142950 682290
rect 143190 682050 143300 682290
rect 143540 682050 143630 682290
rect 143870 682050 143960 682290
rect 144200 682050 144290 682290
rect 144530 682050 144950 682290
rect 145190 682050 145300 682290
rect 145540 682050 145630 682290
rect 145870 682050 145960 682290
rect 146200 682050 146290 682290
rect 146530 682050 146640 682290
rect 146880 682050 146970 682290
rect 147210 682050 147300 682290
rect 147540 682050 147630 682290
rect 147870 682050 147980 682290
rect 148220 682050 148310 682290
rect 148550 682050 148640 682290
rect 148880 682050 148970 682290
rect 149210 682050 149320 682290
rect 149560 682050 149650 682290
rect 149890 682050 149980 682290
rect 150220 682050 150310 682290
rect 150550 682050 150660 682290
rect 150900 682050 150990 682290
rect 151230 682050 151320 682290
rect 151560 682050 151650 682290
rect 151890 682050 152000 682290
rect 152240 682050 152330 682290
rect 152570 682050 152660 682290
rect 152900 682050 152990 682290
rect 153230 682050 153340 682290
rect 153580 682050 153670 682290
rect 153910 682050 154000 682290
rect 154240 682050 154330 682290
rect 154570 682050 154680 682290
rect 154920 682050 155010 682290
rect 155250 682050 155340 682290
rect 155580 682050 155670 682290
rect 155910 682050 155960 682290
rect 110760 681940 155960 682050
rect 110760 681700 110810 681940
rect 111050 681700 111160 681940
rect 111400 681700 111490 681940
rect 111730 681700 111820 681940
rect 112060 681700 112150 681940
rect 112390 681700 112500 681940
rect 112740 681700 112830 681940
rect 113070 681700 113160 681940
rect 113400 681700 113490 681940
rect 113730 681700 113840 681940
rect 114080 681700 114170 681940
rect 114410 681700 114500 681940
rect 114740 681700 114830 681940
rect 115070 681700 115180 681940
rect 115420 681700 115510 681940
rect 115750 681700 115840 681940
rect 116080 681700 116170 681940
rect 116410 681700 116520 681940
rect 116760 681700 116850 681940
rect 117090 681700 117180 681940
rect 117420 681700 117510 681940
rect 117750 681700 117860 681940
rect 118100 681700 118190 681940
rect 118430 681700 118520 681940
rect 118760 681700 118850 681940
rect 119090 681700 119200 681940
rect 119440 681700 119530 681940
rect 119770 681700 119860 681940
rect 120100 681700 120190 681940
rect 120430 681700 120540 681940
rect 120780 681700 120870 681940
rect 121110 681700 121200 681940
rect 121440 681700 121530 681940
rect 121770 681700 122190 681940
rect 122430 681700 122540 681940
rect 122780 681700 122870 681940
rect 123110 681700 123200 681940
rect 123440 681700 123530 681940
rect 123770 681700 123880 681940
rect 124120 681700 124210 681940
rect 124450 681700 124540 681940
rect 124780 681700 124870 681940
rect 125110 681700 125220 681940
rect 125460 681700 125550 681940
rect 125790 681700 125880 681940
rect 126120 681700 126210 681940
rect 126450 681700 126560 681940
rect 126800 681700 126890 681940
rect 127130 681700 127220 681940
rect 127460 681700 127550 681940
rect 127790 681700 127900 681940
rect 128140 681700 128230 681940
rect 128470 681700 128560 681940
rect 128800 681700 128890 681940
rect 129130 681700 129240 681940
rect 129480 681700 129570 681940
rect 129810 681700 129900 681940
rect 130140 681700 130230 681940
rect 130470 681700 130580 681940
rect 130820 681700 130910 681940
rect 131150 681700 131240 681940
rect 131480 681700 131570 681940
rect 131810 681700 131920 681940
rect 132160 681700 132250 681940
rect 132490 681700 132580 681940
rect 132820 681700 132910 681940
rect 133150 681700 133570 681940
rect 133810 681700 133920 681940
rect 134160 681700 134250 681940
rect 134490 681700 134580 681940
rect 134820 681700 134910 681940
rect 135150 681700 135260 681940
rect 135500 681700 135590 681940
rect 135830 681700 135920 681940
rect 136160 681700 136250 681940
rect 136490 681700 136600 681940
rect 136840 681700 136930 681940
rect 137170 681700 137260 681940
rect 137500 681700 137590 681940
rect 137830 681700 137940 681940
rect 138180 681700 138270 681940
rect 138510 681700 138600 681940
rect 138840 681700 138930 681940
rect 139170 681700 139280 681940
rect 139520 681700 139610 681940
rect 139850 681700 139940 681940
rect 140180 681700 140270 681940
rect 140510 681700 140620 681940
rect 140860 681700 140950 681940
rect 141190 681700 141280 681940
rect 141520 681700 141610 681940
rect 141850 681700 141960 681940
rect 142200 681700 142290 681940
rect 142530 681700 142620 681940
rect 142860 681700 142950 681940
rect 143190 681700 143300 681940
rect 143540 681700 143630 681940
rect 143870 681700 143960 681940
rect 144200 681700 144290 681940
rect 144530 681700 144950 681940
rect 145190 681700 145300 681940
rect 145540 681700 145630 681940
rect 145870 681700 145960 681940
rect 146200 681700 146290 681940
rect 146530 681700 146640 681940
rect 146880 681700 146970 681940
rect 147210 681700 147300 681940
rect 147540 681700 147630 681940
rect 147870 681700 147980 681940
rect 148220 681700 148310 681940
rect 148550 681700 148640 681940
rect 148880 681700 148970 681940
rect 149210 681700 149320 681940
rect 149560 681700 149650 681940
rect 149890 681700 149980 681940
rect 150220 681700 150310 681940
rect 150550 681700 150660 681940
rect 150900 681700 150990 681940
rect 151230 681700 151320 681940
rect 151560 681700 151650 681940
rect 151890 681700 152000 681940
rect 152240 681700 152330 681940
rect 152570 681700 152660 681940
rect 152900 681700 152990 681940
rect 153230 681700 153340 681940
rect 153580 681700 153670 681940
rect 153910 681700 154000 681940
rect 154240 681700 154330 681940
rect 154570 681700 154680 681940
rect 154920 681700 155010 681940
rect 155250 681700 155340 681940
rect 155580 681700 155670 681940
rect 155910 681700 155960 681940
rect 110760 681610 155960 681700
rect 110760 681370 110810 681610
rect 111050 681370 111160 681610
rect 111400 681370 111490 681610
rect 111730 681370 111820 681610
rect 112060 681370 112150 681610
rect 112390 681370 112500 681610
rect 112740 681370 112830 681610
rect 113070 681370 113160 681610
rect 113400 681370 113490 681610
rect 113730 681370 113840 681610
rect 114080 681370 114170 681610
rect 114410 681370 114500 681610
rect 114740 681370 114830 681610
rect 115070 681370 115180 681610
rect 115420 681370 115510 681610
rect 115750 681370 115840 681610
rect 116080 681370 116170 681610
rect 116410 681370 116520 681610
rect 116760 681370 116850 681610
rect 117090 681370 117180 681610
rect 117420 681370 117510 681610
rect 117750 681370 117860 681610
rect 118100 681370 118190 681610
rect 118430 681370 118520 681610
rect 118760 681370 118850 681610
rect 119090 681370 119200 681610
rect 119440 681370 119530 681610
rect 119770 681370 119860 681610
rect 120100 681370 120190 681610
rect 120430 681370 120540 681610
rect 120780 681370 120870 681610
rect 121110 681370 121200 681610
rect 121440 681370 121530 681610
rect 121770 681370 122190 681610
rect 122430 681370 122540 681610
rect 122780 681370 122870 681610
rect 123110 681370 123200 681610
rect 123440 681370 123530 681610
rect 123770 681370 123880 681610
rect 124120 681370 124210 681610
rect 124450 681370 124540 681610
rect 124780 681370 124870 681610
rect 125110 681370 125220 681610
rect 125460 681370 125550 681610
rect 125790 681370 125880 681610
rect 126120 681370 126210 681610
rect 126450 681370 126560 681610
rect 126800 681370 126890 681610
rect 127130 681370 127220 681610
rect 127460 681370 127550 681610
rect 127790 681370 127900 681610
rect 128140 681370 128230 681610
rect 128470 681370 128560 681610
rect 128800 681370 128890 681610
rect 129130 681370 129240 681610
rect 129480 681370 129570 681610
rect 129810 681370 129900 681610
rect 130140 681370 130230 681610
rect 130470 681370 130580 681610
rect 130820 681370 130910 681610
rect 131150 681370 131240 681610
rect 131480 681370 131570 681610
rect 131810 681370 131920 681610
rect 132160 681370 132250 681610
rect 132490 681370 132580 681610
rect 132820 681370 132910 681610
rect 133150 681370 133570 681610
rect 133810 681370 133920 681610
rect 134160 681370 134250 681610
rect 134490 681370 134580 681610
rect 134820 681370 134910 681610
rect 135150 681370 135260 681610
rect 135500 681370 135590 681610
rect 135830 681370 135920 681610
rect 136160 681370 136250 681610
rect 136490 681370 136600 681610
rect 136840 681370 136930 681610
rect 137170 681370 137260 681610
rect 137500 681370 137590 681610
rect 137830 681370 137940 681610
rect 138180 681370 138270 681610
rect 138510 681370 138600 681610
rect 138840 681370 138930 681610
rect 139170 681370 139280 681610
rect 139520 681370 139610 681610
rect 139850 681370 139940 681610
rect 140180 681370 140270 681610
rect 140510 681370 140620 681610
rect 140860 681370 140950 681610
rect 141190 681370 141280 681610
rect 141520 681370 141610 681610
rect 141850 681370 141960 681610
rect 142200 681370 142290 681610
rect 142530 681370 142620 681610
rect 142860 681370 142950 681610
rect 143190 681370 143300 681610
rect 143540 681370 143630 681610
rect 143870 681370 143960 681610
rect 144200 681370 144290 681610
rect 144530 681370 144950 681610
rect 145190 681370 145300 681610
rect 145540 681370 145630 681610
rect 145870 681370 145960 681610
rect 146200 681370 146290 681610
rect 146530 681370 146640 681610
rect 146880 681370 146970 681610
rect 147210 681370 147300 681610
rect 147540 681370 147630 681610
rect 147870 681370 147980 681610
rect 148220 681370 148310 681610
rect 148550 681370 148640 681610
rect 148880 681370 148970 681610
rect 149210 681370 149320 681610
rect 149560 681370 149650 681610
rect 149890 681370 149980 681610
rect 150220 681370 150310 681610
rect 150550 681370 150660 681610
rect 150900 681370 150990 681610
rect 151230 681370 151320 681610
rect 151560 681370 151650 681610
rect 151890 681370 152000 681610
rect 152240 681370 152330 681610
rect 152570 681370 152660 681610
rect 152900 681370 152990 681610
rect 153230 681370 153340 681610
rect 153580 681370 153670 681610
rect 153910 681370 154000 681610
rect 154240 681370 154330 681610
rect 154570 681370 154680 681610
rect 154920 681370 155010 681610
rect 155250 681370 155340 681610
rect 155580 681370 155670 681610
rect 155910 681370 155960 681610
rect 110760 681280 155960 681370
rect 110760 681040 110810 681280
rect 111050 681040 111160 681280
rect 111400 681040 111490 681280
rect 111730 681040 111820 681280
rect 112060 681040 112150 681280
rect 112390 681040 112500 681280
rect 112740 681040 112830 681280
rect 113070 681040 113160 681280
rect 113400 681040 113490 681280
rect 113730 681040 113840 681280
rect 114080 681040 114170 681280
rect 114410 681040 114500 681280
rect 114740 681040 114830 681280
rect 115070 681040 115180 681280
rect 115420 681040 115510 681280
rect 115750 681040 115840 681280
rect 116080 681040 116170 681280
rect 116410 681040 116520 681280
rect 116760 681040 116850 681280
rect 117090 681040 117180 681280
rect 117420 681040 117510 681280
rect 117750 681040 117860 681280
rect 118100 681040 118190 681280
rect 118430 681040 118520 681280
rect 118760 681040 118850 681280
rect 119090 681040 119200 681280
rect 119440 681040 119530 681280
rect 119770 681040 119860 681280
rect 120100 681040 120190 681280
rect 120430 681040 120540 681280
rect 120780 681040 120870 681280
rect 121110 681040 121200 681280
rect 121440 681040 121530 681280
rect 121770 681040 122190 681280
rect 122430 681040 122540 681280
rect 122780 681040 122870 681280
rect 123110 681040 123200 681280
rect 123440 681040 123530 681280
rect 123770 681040 123880 681280
rect 124120 681040 124210 681280
rect 124450 681040 124540 681280
rect 124780 681040 124870 681280
rect 125110 681040 125220 681280
rect 125460 681040 125550 681280
rect 125790 681040 125880 681280
rect 126120 681040 126210 681280
rect 126450 681040 126560 681280
rect 126800 681040 126890 681280
rect 127130 681040 127220 681280
rect 127460 681040 127550 681280
rect 127790 681040 127900 681280
rect 128140 681040 128230 681280
rect 128470 681040 128560 681280
rect 128800 681040 128890 681280
rect 129130 681040 129240 681280
rect 129480 681040 129570 681280
rect 129810 681040 129900 681280
rect 130140 681040 130230 681280
rect 130470 681040 130580 681280
rect 130820 681040 130910 681280
rect 131150 681040 131240 681280
rect 131480 681040 131570 681280
rect 131810 681040 131920 681280
rect 132160 681040 132250 681280
rect 132490 681040 132580 681280
rect 132820 681040 132910 681280
rect 133150 681040 133570 681280
rect 133810 681040 133920 681280
rect 134160 681040 134250 681280
rect 134490 681040 134580 681280
rect 134820 681040 134910 681280
rect 135150 681040 135260 681280
rect 135500 681040 135590 681280
rect 135830 681040 135920 681280
rect 136160 681040 136250 681280
rect 136490 681040 136600 681280
rect 136840 681040 136930 681280
rect 137170 681040 137260 681280
rect 137500 681040 137590 681280
rect 137830 681040 137940 681280
rect 138180 681040 138270 681280
rect 138510 681040 138600 681280
rect 138840 681040 138930 681280
rect 139170 681040 139280 681280
rect 139520 681040 139610 681280
rect 139850 681040 139940 681280
rect 140180 681040 140270 681280
rect 140510 681040 140620 681280
rect 140860 681040 140950 681280
rect 141190 681040 141280 681280
rect 141520 681040 141610 681280
rect 141850 681040 141960 681280
rect 142200 681040 142290 681280
rect 142530 681040 142620 681280
rect 142860 681040 142950 681280
rect 143190 681040 143300 681280
rect 143540 681040 143630 681280
rect 143870 681040 143960 681280
rect 144200 681040 144290 681280
rect 144530 681040 144950 681280
rect 145190 681040 145300 681280
rect 145540 681040 145630 681280
rect 145870 681040 145960 681280
rect 146200 681040 146290 681280
rect 146530 681040 146640 681280
rect 146880 681040 146970 681280
rect 147210 681040 147300 681280
rect 147540 681040 147630 681280
rect 147870 681040 147980 681280
rect 148220 681040 148310 681280
rect 148550 681040 148640 681280
rect 148880 681040 148970 681280
rect 149210 681040 149320 681280
rect 149560 681040 149650 681280
rect 149890 681040 149980 681280
rect 150220 681040 150310 681280
rect 150550 681040 150660 681280
rect 150900 681040 150990 681280
rect 151230 681040 151320 681280
rect 151560 681040 151650 681280
rect 151890 681040 152000 681280
rect 152240 681040 152330 681280
rect 152570 681040 152660 681280
rect 152900 681040 152990 681280
rect 153230 681040 153340 681280
rect 153580 681040 153670 681280
rect 153910 681040 154000 681280
rect 154240 681040 154330 681280
rect 154570 681040 154680 681280
rect 154920 681040 155010 681280
rect 155250 681040 155340 681280
rect 155580 681040 155670 681280
rect 155910 681040 155960 681280
rect 110760 680950 155960 681040
rect 110760 680710 110810 680950
rect 111050 680710 111160 680950
rect 111400 680710 111490 680950
rect 111730 680710 111820 680950
rect 112060 680710 112150 680950
rect 112390 680710 112500 680950
rect 112740 680710 112830 680950
rect 113070 680710 113160 680950
rect 113400 680710 113490 680950
rect 113730 680710 113840 680950
rect 114080 680710 114170 680950
rect 114410 680710 114500 680950
rect 114740 680710 114830 680950
rect 115070 680710 115180 680950
rect 115420 680710 115510 680950
rect 115750 680710 115840 680950
rect 116080 680710 116170 680950
rect 116410 680710 116520 680950
rect 116760 680710 116850 680950
rect 117090 680710 117180 680950
rect 117420 680710 117510 680950
rect 117750 680710 117860 680950
rect 118100 680710 118190 680950
rect 118430 680710 118520 680950
rect 118760 680710 118850 680950
rect 119090 680710 119200 680950
rect 119440 680710 119530 680950
rect 119770 680710 119860 680950
rect 120100 680710 120190 680950
rect 120430 680710 120540 680950
rect 120780 680710 120870 680950
rect 121110 680710 121200 680950
rect 121440 680710 121530 680950
rect 121770 680710 122190 680950
rect 122430 680710 122540 680950
rect 122780 680710 122870 680950
rect 123110 680710 123200 680950
rect 123440 680710 123530 680950
rect 123770 680710 123880 680950
rect 124120 680710 124210 680950
rect 124450 680710 124540 680950
rect 124780 680710 124870 680950
rect 125110 680710 125220 680950
rect 125460 680710 125550 680950
rect 125790 680710 125880 680950
rect 126120 680710 126210 680950
rect 126450 680710 126560 680950
rect 126800 680710 126890 680950
rect 127130 680710 127220 680950
rect 127460 680710 127550 680950
rect 127790 680710 127900 680950
rect 128140 680710 128230 680950
rect 128470 680710 128560 680950
rect 128800 680710 128890 680950
rect 129130 680710 129240 680950
rect 129480 680710 129570 680950
rect 129810 680710 129900 680950
rect 130140 680710 130230 680950
rect 130470 680710 130580 680950
rect 130820 680710 130910 680950
rect 131150 680710 131240 680950
rect 131480 680710 131570 680950
rect 131810 680710 131920 680950
rect 132160 680710 132250 680950
rect 132490 680710 132580 680950
rect 132820 680710 132910 680950
rect 133150 680710 133570 680950
rect 133810 680710 133920 680950
rect 134160 680710 134250 680950
rect 134490 680710 134580 680950
rect 134820 680710 134910 680950
rect 135150 680710 135260 680950
rect 135500 680710 135590 680950
rect 135830 680710 135920 680950
rect 136160 680710 136250 680950
rect 136490 680710 136600 680950
rect 136840 680710 136930 680950
rect 137170 680710 137260 680950
rect 137500 680710 137590 680950
rect 137830 680710 137940 680950
rect 138180 680710 138270 680950
rect 138510 680710 138600 680950
rect 138840 680710 138930 680950
rect 139170 680710 139280 680950
rect 139520 680710 139610 680950
rect 139850 680710 139940 680950
rect 140180 680710 140270 680950
rect 140510 680710 140620 680950
rect 140860 680710 140950 680950
rect 141190 680710 141280 680950
rect 141520 680710 141610 680950
rect 141850 680710 141960 680950
rect 142200 680710 142290 680950
rect 142530 680710 142620 680950
rect 142860 680710 142950 680950
rect 143190 680710 143300 680950
rect 143540 680710 143630 680950
rect 143870 680710 143960 680950
rect 144200 680710 144290 680950
rect 144530 680710 144950 680950
rect 145190 680710 145300 680950
rect 145540 680710 145630 680950
rect 145870 680710 145960 680950
rect 146200 680710 146290 680950
rect 146530 680710 146640 680950
rect 146880 680710 146970 680950
rect 147210 680710 147300 680950
rect 147540 680710 147630 680950
rect 147870 680710 147980 680950
rect 148220 680710 148310 680950
rect 148550 680710 148640 680950
rect 148880 680710 148970 680950
rect 149210 680710 149320 680950
rect 149560 680710 149650 680950
rect 149890 680710 149980 680950
rect 150220 680710 150310 680950
rect 150550 680710 150660 680950
rect 150900 680710 150990 680950
rect 151230 680710 151320 680950
rect 151560 680710 151650 680950
rect 151890 680710 152000 680950
rect 152240 680710 152330 680950
rect 152570 680710 152660 680950
rect 152900 680710 152990 680950
rect 153230 680710 153340 680950
rect 153580 680710 153670 680950
rect 153910 680710 154000 680950
rect 154240 680710 154330 680950
rect 154570 680710 154680 680950
rect 154920 680710 155010 680950
rect 155250 680710 155340 680950
rect 155580 680710 155670 680950
rect 155910 680710 155960 680950
rect 110760 680600 155960 680710
rect 110760 680360 110810 680600
rect 111050 680360 111160 680600
rect 111400 680360 111490 680600
rect 111730 680360 111820 680600
rect 112060 680360 112150 680600
rect 112390 680360 112500 680600
rect 112740 680360 112830 680600
rect 113070 680360 113160 680600
rect 113400 680360 113490 680600
rect 113730 680360 113840 680600
rect 114080 680360 114170 680600
rect 114410 680360 114500 680600
rect 114740 680360 114830 680600
rect 115070 680360 115180 680600
rect 115420 680360 115510 680600
rect 115750 680360 115840 680600
rect 116080 680360 116170 680600
rect 116410 680360 116520 680600
rect 116760 680360 116850 680600
rect 117090 680360 117180 680600
rect 117420 680360 117510 680600
rect 117750 680360 117860 680600
rect 118100 680360 118190 680600
rect 118430 680360 118520 680600
rect 118760 680360 118850 680600
rect 119090 680360 119200 680600
rect 119440 680360 119530 680600
rect 119770 680360 119860 680600
rect 120100 680360 120190 680600
rect 120430 680360 120540 680600
rect 120780 680360 120870 680600
rect 121110 680360 121200 680600
rect 121440 680360 121530 680600
rect 121770 680360 122190 680600
rect 122430 680360 122540 680600
rect 122780 680360 122870 680600
rect 123110 680360 123200 680600
rect 123440 680360 123530 680600
rect 123770 680360 123880 680600
rect 124120 680360 124210 680600
rect 124450 680360 124540 680600
rect 124780 680360 124870 680600
rect 125110 680360 125220 680600
rect 125460 680360 125550 680600
rect 125790 680360 125880 680600
rect 126120 680360 126210 680600
rect 126450 680360 126560 680600
rect 126800 680360 126890 680600
rect 127130 680360 127220 680600
rect 127460 680360 127550 680600
rect 127790 680360 127900 680600
rect 128140 680360 128230 680600
rect 128470 680360 128560 680600
rect 128800 680360 128890 680600
rect 129130 680360 129240 680600
rect 129480 680360 129570 680600
rect 129810 680360 129900 680600
rect 130140 680360 130230 680600
rect 130470 680360 130580 680600
rect 130820 680360 130910 680600
rect 131150 680360 131240 680600
rect 131480 680360 131570 680600
rect 131810 680360 131920 680600
rect 132160 680360 132250 680600
rect 132490 680360 132580 680600
rect 132820 680360 132910 680600
rect 133150 680360 133570 680600
rect 133810 680360 133920 680600
rect 134160 680360 134250 680600
rect 134490 680360 134580 680600
rect 134820 680360 134910 680600
rect 135150 680360 135260 680600
rect 135500 680360 135590 680600
rect 135830 680360 135920 680600
rect 136160 680360 136250 680600
rect 136490 680360 136600 680600
rect 136840 680360 136930 680600
rect 137170 680360 137260 680600
rect 137500 680360 137590 680600
rect 137830 680360 137940 680600
rect 138180 680360 138270 680600
rect 138510 680360 138600 680600
rect 138840 680360 138930 680600
rect 139170 680360 139280 680600
rect 139520 680360 139610 680600
rect 139850 680360 139940 680600
rect 140180 680360 140270 680600
rect 140510 680360 140620 680600
rect 140860 680360 140950 680600
rect 141190 680360 141280 680600
rect 141520 680360 141610 680600
rect 141850 680360 141960 680600
rect 142200 680360 142290 680600
rect 142530 680360 142620 680600
rect 142860 680360 142950 680600
rect 143190 680360 143300 680600
rect 143540 680360 143630 680600
rect 143870 680360 143960 680600
rect 144200 680360 144290 680600
rect 144530 680360 144950 680600
rect 145190 680360 145300 680600
rect 145540 680360 145630 680600
rect 145870 680360 145960 680600
rect 146200 680360 146290 680600
rect 146530 680360 146640 680600
rect 146880 680360 146970 680600
rect 147210 680360 147300 680600
rect 147540 680360 147630 680600
rect 147870 680360 147980 680600
rect 148220 680360 148310 680600
rect 148550 680360 148640 680600
rect 148880 680360 148970 680600
rect 149210 680360 149320 680600
rect 149560 680360 149650 680600
rect 149890 680360 149980 680600
rect 150220 680360 150310 680600
rect 150550 680360 150660 680600
rect 150900 680360 150990 680600
rect 151230 680360 151320 680600
rect 151560 680360 151650 680600
rect 151890 680360 152000 680600
rect 152240 680360 152330 680600
rect 152570 680360 152660 680600
rect 152900 680360 152990 680600
rect 153230 680360 153340 680600
rect 153580 680360 153670 680600
rect 153910 680360 154000 680600
rect 154240 680360 154330 680600
rect 154570 680360 154680 680600
rect 154920 680360 155010 680600
rect 155250 680360 155340 680600
rect 155580 680360 155670 680600
rect 155910 680360 155960 680600
rect 110760 680270 155960 680360
rect 110760 680030 110810 680270
rect 111050 680030 111160 680270
rect 111400 680030 111490 680270
rect 111730 680030 111820 680270
rect 112060 680030 112150 680270
rect 112390 680030 112500 680270
rect 112740 680030 112830 680270
rect 113070 680030 113160 680270
rect 113400 680030 113490 680270
rect 113730 680030 113840 680270
rect 114080 680030 114170 680270
rect 114410 680030 114500 680270
rect 114740 680030 114830 680270
rect 115070 680030 115180 680270
rect 115420 680030 115510 680270
rect 115750 680030 115840 680270
rect 116080 680030 116170 680270
rect 116410 680030 116520 680270
rect 116760 680030 116850 680270
rect 117090 680030 117180 680270
rect 117420 680030 117510 680270
rect 117750 680030 117860 680270
rect 118100 680030 118190 680270
rect 118430 680030 118520 680270
rect 118760 680030 118850 680270
rect 119090 680030 119200 680270
rect 119440 680030 119530 680270
rect 119770 680030 119860 680270
rect 120100 680030 120190 680270
rect 120430 680030 120540 680270
rect 120780 680030 120870 680270
rect 121110 680030 121200 680270
rect 121440 680030 121530 680270
rect 121770 680030 122190 680270
rect 122430 680030 122540 680270
rect 122780 680030 122870 680270
rect 123110 680030 123200 680270
rect 123440 680030 123530 680270
rect 123770 680030 123880 680270
rect 124120 680030 124210 680270
rect 124450 680030 124540 680270
rect 124780 680030 124870 680270
rect 125110 680030 125220 680270
rect 125460 680030 125550 680270
rect 125790 680030 125880 680270
rect 126120 680030 126210 680270
rect 126450 680030 126560 680270
rect 126800 680030 126890 680270
rect 127130 680030 127220 680270
rect 127460 680030 127550 680270
rect 127790 680030 127900 680270
rect 128140 680030 128230 680270
rect 128470 680030 128560 680270
rect 128800 680030 128890 680270
rect 129130 680030 129240 680270
rect 129480 680030 129570 680270
rect 129810 680030 129900 680270
rect 130140 680030 130230 680270
rect 130470 680030 130580 680270
rect 130820 680030 130910 680270
rect 131150 680030 131240 680270
rect 131480 680030 131570 680270
rect 131810 680030 131920 680270
rect 132160 680030 132250 680270
rect 132490 680030 132580 680270
rect 132820 680030 132910 680270
rect 133150 680030 133570 680270
rect 133810 680030 133920 680270
rect 134160 680030 134250 680270
rect 134490 680030 134580 680270
rect 134820 680030 134910 680270
rect 135150 680030 135260 680270
rect 135500 680030 135590 680270
rect 135830 680030 135920 680270
rect 136160 680030 136250 680270
rect 136490 680030 136600 680270
rect 136840 680030 136930 680270
rect 137170 680030 137260 680270
rect 137500 680030 137590 680270
rect 137830 680030 137940 680270
rect 138180 680030 138270 680270
rect 138510 680030 138600 680270
rect 138840 680030 138930 680270
rect 139170 680030 139280 680270
rect 139520 680030 139610 680270
rect 139850 680030 139940 680270
rect 140180 680030 140270 680270
rect 140510 680030 140620 680270
rect 140860 680030 140950 680270
rect 141190 680030 141280 680270
rect 141520 680030 141610 680270
rect 141850 680030 141960 680270
rect 142200 680030 142290 680270
rect 142530 680030 142620 680270
rect 142860 680030 142950 680270
rect 143190 680030 143300 680270
rect 143540 680030 143630 680270
rect 143870 680030 143960 680270
rect 144200 680030 144290 680270
rect 144530 680030 144950 680270
rect 145190 680030 145300 680270
rect 145540 680030 145630 680270
rect 145870 680030 145960 680270
rect 146200 680030 146290 680270
rect 146530 680030 146640 680270
rect 146880 680030 146970 680270
rect 147210 680030 147300 680270
rect 147540 680030 147630 680270
rect 147870 680030 147980 680270
rect 148220 680030 148310 680270
rect 148550 680030 148640 680270
rect 148880 680030 148970 680270
rect 149210 680030 149320 680270
rect 149560 680030 149650 680270
rect 149890 680030 149980 680270
rect 150220 680030 150310 680270
rect 150550 680030 150660 680270
rect 150900 680030 150990 680270
rect 151230 680030 151320 680270
rect 151560 680030 151650 680270
rect 151890 680030 152000 680270
rect 152240 680030 152330 680270
rect 152570 680030 152660 680270
rect 152900 680030 152990 680270
rect 153230 680030 153340 680270
rect 153580 680030 153670 680270
rect 153910 680030 154000 680270
rect 154240 680030 154330 680270
rect 154570 680030 154680 680270
rect 154920 680030 155010 680270
rect 155250 680030 155340 680270
rect 155580 680030 155670 680270
rect 155910 680030 155960 680270
rect 110760 679940 155960 680030
rect 110760 679700 110810 679940
rect 111050 679700 111160 679940
rect 111400 679700 111490 679940
rect 111730 679700 111820 679940
rect 112060 679700 112150 679940
rect 112390 679700 112500 679940
rect 112740 679700 112830 679940
rect 113070 679700 113160 679940
rect 113400 679700 113490 679940
rect 113730 679700 113840 679940
rect 114080 679700 114170 679940
rect 114410 679700 114500 679940
rect 114740 679700 114830 679940
rect 115070 679700 115180 679940
rect 115420 679700 115510 679940
rect 115750 679700 115840 679940
rect 116080 679700 116170 679940
rect 116410 679700 116520 679940
rect 116760 679700 116850 679940
rect 117090 679700 117180 679940
rect 117420 679700 117510 679940
rect 117750 679700 117860 679940
rect 118100 679700 118190 679940
rect 118430 679700 118520 679940
rect 118760 679700 118850 679940
rect 119090 679700 119200 679940
rect 119440 679700 119530 679940
rect 119770 679700 119860 679940
rect 120100 679700 120190 679940
rect 120430 679700 120540 679940
rect 120780 679700 120870 679940
rect 121110 679700 121200 679940
rect 121440 679700 121530 679940
rect 121770 679700 122190 679940
rect 122430 679700 122540 679940
rect 122780 679700 122870 679940
rect 123110 679700 123200 679940
rect 123440 679700 123530 679940
rect 123770 679700 123880 679940
rect 124120 679700 124210 679940
rect 124450 679700 124540 679940
rect 124780 679700 124870 679940
rect 125110 679700 125220 679940
rect 125460 679700 125550 679940
rect 125790 679700 125880 679940
rect 126120 679700 126210 679940
rect 126450 679700 126560 679940
rect 126800 679700 126890 679940
rect 127130 679700 127220 679940
rect 127460 679700 127550 679940
rect 127790 679700 127900 679940
rect 128140 679700 128230 679940
rect 128470 679700 128560 679940
rect 128800 679700 128890 679940
rect 129130 679700 129240 679940
rect 129480 679700 129570 679940
rect 129810 679700 129900 679940
rect 130140 679700 130230 679940
rect 130470 679700 130580 679940
rect 130820 679700 130910 679940
rect 131150 679700 131240 679940
rect 131480 679700 131570 679940
rect 131810 679700 131920 679940
rect 132160 679700 132250 679940
rect 132490 679700 132580 679940
rect 132820 679700 132910 679940
rect 133150 679700 133570 679940
rect 133810 679700 133920 679940
rect 134160 679700 134250 679940
rect 134490 679700 134580 679940
rect 134820 679700 134910 679940
rect 135150 679700 135260 679940
rect 135500 679700 135590 679940
rect 135830 679700 135920 679940
rect 136160 679700 136250 679940
rect 136490 679700 136600 679940
rect 136840 679700 136930 679940
rect 137170 679700 137260 679940
rect 137500 679700 137590 679940
rect 137830 679700 137940 679940
rect 138180 679700 138270 679940
rect 138510 679700 138600 679940
rect 138840 679700 138930 679940
rect 139170 679700 139280 679940
rect 139520 679700 139610 679940
rect 139850 679700 139940 679940
rect 140180 679700 140270 679940
rect 140510 679700 140620 679940
rect 140860 679700 140950 679940
rect 141190 679700 141280 679940
rect 141520 679700 141610 679940
rect 141850 679700 141960 679940
rect 142200 679700 142290 679940
rect 142530 679700 142620 679940
rect 142860 679700 142950 679940
rect 143190 679700 143300 679940
rect 143540 679700 143630 679940
rect 143870 679700 143960 679940
rect 144200 679700 144290 679940
rect 144530 679700 144950 679940
rect 145190 679700 145300 679940
rect 145540 679700 145630 679940
rect 145870 679700 145960 679940
rect 146200 679700 146290 679940
rect 146530 679700 146640 679940
rect 146880 679700 146970 679940
rect 147210 679700 147300 679940
rect 147540 679700 147630 679940
rect 147870 679700 147980 679940
rect 148220 679700 148310 679940
rect 148550 679700 148640 679940
rect 148880 679700 148970 679940
rect 149210 679700 149320 679940
rect 149560 679700 149650 679940
rect 149890 679700 149980 679940
rect 150220 679700 150310 679940
rect 150550 679700 150660 679940
rect 150900 679700 150990 679940
rect 151230 679700 151320 679940
rect 151560 679700 151650 679940
rect 151890 679700 152000 679940
rect 152240 679700 152330 679940
rect 152570 679700 152660 679940
rect 152900 679700 152990 679940
rect 153230 679700 153340 679940
rect 153580 679700 153670 679940
rect 153910 679700 154000 679940
rect 154240 679700 154330 679940
rect 154570 679700 154680 679940
rect 154920 679700 155010 679940
rect 155250 679700 155340 679940
rect 155580 679700 155670 679940
rect 155910 679700 155960 679940
rect 110760 679610 155960 679700
rect 110760 679370 110810 679610
rect 111050 679370 111160 679610
rect 111400 679370 111490 679610
rect 111730 679370 111820 679610
rect 112060 679370 112150 679610
rect 112390 679370 112500 679610
rect 112740 679370 112830 679610
rect 113070 679370 113160 679610
rect 113400 679370 113490 679610
rect 113730 679370 113840 679610
rect 114080 679370 114170 679610
rect 114410 679370 114500 679610
rect 114740 679370 114830 679610
rect 115070 679370 115180 679610
rect 115420 679370 115510 679610
rect 115750 679370 115840 679610
rect 116080 679370 116170 679610
rect 116410 679370 116520 679610
rect 116760 679370 116850 679610
rect 117090 679370 117180 679610
rect 117420 679370 117510 679610
rect 117750 679370 117860 679610
rect 118100 679370 118190 679610
rect 118430 679370 118520 679610
rect 118760 679370 118850 679610
rect 119090 679370 119200 679610
rect 119440 679370 119530 679610
rect 119770 679370 119860 679610
rect 120100 679370 120190 679610
rect 120430 679370 120540 679610
rect 120780 679370 120870 679610
rect 121110 679370 121200 679610
rect 121440 679370 121530 679610
rect 121770 679370 122190 679610
rect 122430 679370 122540 679610
rect 122780 679370 122870 679610
rect 123110 679370 123200 679610
rect 123440 679370 123530 679610
rect 123770 679370 123880 679610
rect 124120 679370 124210 679610
rect 124450 679370 124540 679610
rect 124780 679370 124870 679610
rect 125110 679370 125220 679610
rect 125460 679370 125550 679610
rect 125790 679370 125880 679610
rect 126120 679370 126210 679610
rect 126450 679370 126560 679610
rect 126800 679370 126890 679610
rect 127130 679370 127220 679610
rect 127460 679370 127550 679610
rect 127790 679370 127900 679610
rect 128140 679370 128230 679610
rect 128470 679370 128560 679610
rect 128800 679370 128890 679610
rect 129130 679370 129240 679610
rect 129480 679370 129570 679610
rect 129810 679370 129900 679610
rect 130140 679370 130230 679610
rect 130470 679370 130580 679610
rect 130820 679370 130910 679610
rect 131150 679370 131240 679610
rect 131480 679370 131570 679610
rect 131810 679370 131920 679610
rect 132160 679370 132250 679610
rect 132490 679370 132580 679610
rect 132820 679370 132910 679610
rect 133150 679370 133570 679610
rect 133810 679370 133920 679610
rect 134160 679370 134250 679610
rect 134490 679370 134580 679610
rect 134820 679370 134910 679610
rect 135150 679370 135260 679610
rect 135500 679370 135590 679610
rect 135830 679370 135920 679610
rect 136160 679370 136250 679610
rect 136490 679370 136600 679610
rect 136840 679370 136930 679610
rect 137170 679370 137260 679610
rect 137500 679370 137590 679610
rect 137830 679370 137940 679610
rect 138180 679370 138270 679610
rect 138510 679370 138600 679610
rect 138840 679370 138930 679610
rect 139170 679370 139280 679610
rect 139520 679370 139610 679610
rect 139850 679370 139940 679610
rect 140180 679370 140270 679610
rect 140510 679370 140620 679610
rect 140860 679370 140950 679610
rect 141190 679370 141280 679610
rect 141520 679370 141610 679610
rect 141850 679370 141960 679610
rect 142200 679370 142290 679610
rect 142530 679370 142620 679610
rect 142860 679370 142950 679610
rect 143190 679370 143300 679610
rect 143540 679370 143630 679610
rect 143870 679370 143960 679610
rect 144200 679370 144290 679610
rect 144530 679370 144950 679610
rect 145190 679370 145300 679610
rect 145540 679370 145630 679610
rect 145870 679370 145960 679610
rect 146200 679370 146290 679610
rect 146530 679370 146640 679610
rect 146880 679370 146970 679610
rect 147210 679370 147300 679610
rect 147540 679370 147630 679610
rect 147870 679370 147980 679610
rect 148220 679370 148310 679610
rect 148550 679370 148640 679610
rect 148880 679370 148970 679610
rect 149210 679370 149320 679610
rect 149560 679370 149650 679610
rect 149890 679370 149980 679610
rect 150220 679370 150310 679610
rect 150550 679370 150660 679610
rect 150900 679370 150990 679610
rect 151230 679370 151320 679610
rect 151560 679370 151650 679610
rect 151890 679370 152000 679610
rect 152240 679370 152330 679610
rect 152570 679370 152660 679610
rect 152900 679370 152990 679610
rect 153230 679370 153340 679610
rect 153580 679370 153670 679610
rect 153910 679370 154000 679610
rect 154240 679370 154330 679610
rect 154570 679370 154680 679610
rect 154920 679370 155010 679610
rect 155250 679370 155340 679610
rect 155580 679370 155670 679610
rect 155910 679370 155960 679610
rect 110760 679260 155960 679370
rect 110760 679147 110810 679260
rect 103643 679020 110810 679147
rect 111050 679020 111160 679260
rect 111400 679020 111490 679260
rect 111730 679020 111820 679260
rect 112060 679020 112150 679260
rect 112390 679020 112500 679260
rect 112740 679020 112830 679260
rect 113070 679020 113160 679260
rect 113400 679020 113490 679260
rect 113730 679020 113840 679260
rect 114080 679020 114170 679260
rect 114410 679020 114500 679260
rect 114740 679020 114830 679260
rect 115070 679020 115180 679260
rect 115420 679020 115510 679260
rect 115750 679020 115840 679260
rect 116080 679020 116170 679260
rect 116410 679020 116520 679260
rect 116760 679020 116850 679260
rect 117090 679020 117180 679260
rect 117420 679020 117510 679260
rect 117750 679020 117860 679260
rect 118100 679020 118190 679260
rect 118430 679020 118520 679260
rect 118760 679020 118850 679260
rect 119090 679020 119200 679260
rect 119440 679020 119530 679260
rect 119770 679020 119860 679260
rect 120100 679020 120190 679260
rect 120430 679020 120540 679260
rect 120780 679020 120870 679260
rect 121110 679020 121200 679260
rect 121440 679020 121530 679260
rect 121770 679020 122190 679260
rect 122430 679020 122540 679260
rect 122780 679020 122870 679260
rect 123110 679020 123200 679260
rect 123440 679020 123530 679260
rect 123770 679020 123880 679260
rect 124120 679020 124210 679260
rect 124450 679020 124540 679260
rect 124780 679020 124870 679260
rect 125110 679020 125220 679260
rect 125460 679020 125550 679260
rect 125790 679020 125880 679260
rect 126120 679020 126210 679260
rect 126450 679020 126560 679260
rect 126800 679020 126890 679260
rect 127130 679020 127220 679260
rect 127460 679020 127550 679260
rect 127790 679020 127900 679260
rect 128140 679020 128230 679260
rect 128470 679020 128560 679260
rect 128800 679020 128890 679260
rect 129130 679020 129240 679260
rect 129480 679020 129570 679260
rect 129810 679020 129900 679260
rect 130140 679020 130230 679260
rect 130470 679020 130580 679260
rect 130820 679020 130910 679260
rect 131150 679020 131240 679260
rect 131480 679020 131570 679260
rect 131810 679020 131920 679260
rect 132160 679020 132250 679260
rect 132490 679020 132580 679260
rect 132820 679020 132910 679260
rect 133150 679020 133570 679260
rect 133810 679020 133920 679260
rect 134160 679020 134250 679260
rect 134490 679020 134580 679260
rect 134820 679020 134910 679260
rect 135150 679020 135260 679260
rect 135500 679020 135590 679260
rect 135830 679020 135920 679260
rect 136160 679020 136250 679260
rect 136490 679020 136600 679260
rect 136840 679020 136930 679260
rect 137170 679020 137260 679260
rect 137500 679020 137590 679260
rect 137830 679020 137940 679260
rect 138180 679020 138270 679260
rect 138510 679020 138600 679260
rect 138840 679020 138930 679260
rect 139170 679020 139280 679260
rect 139520 679020 139610 679260
rect 139850 679020 139940 679260
rect 140180 679020 140270 679260
rect 140510 679020 140620 679260
rect 140860 679020 140950 679260
rect 141190 679020 141280 679260
rect 141520 679020 141610 679260
rect 141850 679020 141960 679260
rect 142200 679020 142290 679260
rect 142530 679020 142620 679260
rect 142860 679020 142950 679260
rect 143190 679020 143300 679260
rect 143540 679020 143630 679260
rect 143870 679020 143960 679260
rect 144200 679020 144290 679260
rect 144530 679020 144950 679260
rect 145190 679020 145300 679260
rect 145540 679020 145630 679260
rect 145870 679020 145960 679260
rect 146200 679020 146290 679260
rect 146530 679020 146640 679260
rect 146880 679020 146970 679260
rect 147210 679020 147300 679260
rect 147540 679020 147630 679260
rect 147870 679020 147980 679260
rect 148220 679020 148310 679260
rect 148550 679020 148640 679260
rect 148880 679020 148970 679260
rect 149210 679020 149320 679260
rect 149560 679020 149650 679260
rect 149890 679020 149980 679260
rect 150220 679020 150310 679260
rect 150550 679020 150660 679260
rect 150900 679020 150990 679260
rect 151230 679020 151320 679260
rect 151560 679020 151650 679260
rect 151890 679020 152000 679260
rect 152240 679020 152330 679260
rect 152570 679020 152660 679260
rect 152900 679020 152990 679260
rect 153230 679020 153340 679260
rect 153580 679020 153670 679260
rect 153910 679020 154000 679260
rect 154240 679020 154330 679260
rect 154570 679020 154680 679260
rect 154920 679020 155010 679260
rect 155250 679020 155340 679260
rect 155580 679020 155670 679260
rect 155910 679147 155960 679260
rect 157440 679147 162436 686032
rect 321017 681560 321497 702300
rect 212764 681080 321497 681560
rect 212764 680040 212924 681080
rect 415740 679850 416220 702680
rect 230810 679370 416220 679850
rect 467200 703150 467220 703220
rect 467290 703150 467320 703220
rect 467390 703150 467420 703220
rect 467490 703150 467520 703220
rect 467200 703130 467520 703150
rect 467200 703060 467220 703130
rect 467290 703060 467320 703130
rect 467390 703060 467420 703130
rect 467490 703060 467520 703130
rect 155910 679020 162436 679147
rect 103643 678980 162436 679020
rect 103643 678740 107220 678980
rect 107480 678740 107580 678980
rect 107840 678740 107940 678980
rect 108200 678740 108300 678980
rect 108560 678979 162436 678980
rect 108560 678930 157520 678979
rect 108560 678740 110810 678930
rect 103643 678690 110810 678740
rect 111050 678690 111160 678930
rect 111400 678690 111490 678930
rect 111730 678690 111820 678930
rect 112060 678690 112150 678930
rect 112390 678690 112500 678930
rect 112740 678690 112830 678930
rect 113070 678690 113160 678930
rect 113400 678690 113490 678930
rect 113730 678690 113840 678930
rect 114080 678690 114170 678930
rect 114410 678690 114500 678930
rect 114740 678690 114830 678930
rect 115070 678690 115180 678930
rect 115420 678690 115510 678930
rect 115750 678690 115840 678930
rect 116080 678690 116170 678930
rect 116410 678690 116520 678930
rect 116760 678690 116850 678930
rect 117090 678690 117180 678930
rect 117420 678690 117510 678930
rect 117750 678690 117860 678930
rect 118100 678690 118190 678930
rect 118430 678690 118520 678930
rect 118760 678690 118850 678930
rect 119090 678690 119200 678930
rect 119440 678690 119530 678930
rect 119770 678690 119860 678930
rect 120100 678690 120190 678930
rect 120430 678690 120540 678930
rect 120780 678690 120870 678930
rect 121110 678690 121200 678930
rect 121440 678690 121530 678930
rect 121770 678690 122190 678930
rect 122430 678690 122540 678930
rect 122780 678690 122870 678930
rect 123110 678690 123200 678930
rect 123440 678690 123530 678930
rect 123770 678690 123880 678930
rect 124120 678690 124210 678930
rect 124450 678690 124540 678930
rect 124780 678690 124870 678930
rect 125110 678690 125220 678930
rect 125460 678690 125550 678930
rect 125790 678690 125880 678930
rect 126120 678690 126210 678930
rect 126450 678690 126560 678930
rect 126800 678690 126890 678930
rect 127130 678690 127220 678930
rect 127460 678690 127550 678930
rect 127790 678690 127900 678930
rect 128140 678690 128230 678930
rect 128470 678690 128560 678930
rect 128800 678690 128890 678930
rect 129130 678690 129240 678930
rect 129480 678690 129570 678930
rect 129810 678690 129900 678930
rect 130140 678690 130230 678930
rect 130470 678690 130580 678930
rect 130820 678690 130910 678930
rect 131150 678690 131240 678930
rect 131480 678690 131570 678930
rect 131810 678690 131920 678930
rect 132160 678690 132250 678930
rect 132490 678690 132580 678930
rect 132820 678690 132910 678930
rect 133150 678690 133570 678930
rect 133810 678690 133920 678930
rect 134160 678690 134250 678930
rect 134490 678690 134580 678930
rect 134820 678690 134910 678930
rect 135150 678690 135260 678930
rect 135500 678690 135590 678930
rect 135830 678690 135920 678930
rect 136160 678690 136250 678930
rect 136490 678690 136600 678930
rect 136840 678690 136930 678930
rect 137170 678690 137260 678930
rect 137500 678690 137590 678930
rect 137830 678690 137940 678930
rect 138180 678690 138270 678930
rect 138510 678690 138600 678930
rect 138840 678690 138930 678930
rect 139170 678690 139280 678930
rect 139520 678690 139610 678930
rect 139850 678690 139940 678930
rect 140180 678690 140270 678930
rect 140510 678690 140620 678930
rect 140860 678690 140950 678930
rect 141190 678690 141280 678930
rect 141520 678690 141610 678930
rect 141850 678690 141960 678930
rect 142200 678690 142290 678930
rect 142530 678690 142620 678930
rect 142860 678690 142950 678930
rect 143190 678690 143300 678930
rect 143540 678690 143630 678930
rect 143870 678690 143960 678930
rect 144200 678690 144290 678930
rect 144530 678690 144950 678930
rect 145190 678690 145300 678930
rect 145540 678690 145630 678930
rect 145870 678690 145960 678930
rect 146200 678690 146290 678930
rect 146530 678690 146640 678930
rect 146880 678690 146970 678930
rect 147210 678690 147300 678930
rect 147540 678690 147630 678930
rect 147870 678690 147980 678930
rect 148220 678690 148310 678930
rect 148550 678690 148640 678930
rect 148880 678690 148970 678930
rect 149210 678690 149320 678930
rect 149560 678690 149650 678930
rect 149890 678690 149980 678930
rect 150220 678690 150310 678930
rect 150550 678690 150660 678930
rect 150900 678690 150990 678930
rect 151230 678690 151320 678930
rect 151560 678690 151650 678930
rect 151890 678690 152000 678930
rect 152240 678690 152330 678930
rect 152570 678690 152660 678930
rect 152900 678690 152990 678930
rect 153230 678690 153340 678930
rect 153580 678690 153670 678930
rect 153910 678690 154000 678930
rect 154240 678690 154330 678930
rect 154570 678690 154680 678930
rect 154920 678690 155010 678930
rect 155250 678690 155340 678930
rect 155580 678690 155670 678930
rect 155910 678739 157520 678930
rect 157780 678739 157880 678979
rect 158140 678739 158240 678979
rect 158500 678739 158600 678979
rect 158860 678739 162436 678979
rect 155910 678690 162436 678739
rect 103643 678640 162436 678690
rect 103643 678400 107220 678640
rect 107480 678400 107580 678640
rect 107840 678400 107940 678640
rect 108200 678400 108300 678640
rect 108560 678639 162436 678640
rect 108560 678600 157520 678639
rect 108560 678400 110810 678600
rect 103643 678360 110810 678400
rect 111050 678360 111160 678600
rect 111400 678360 111490 678600
rect 111730 678360 111820 678600
rect 112060 678360 112150 678600
rect 112390 678360 112500 678600
rect 112740 678360 112830 678600
rect 113070 678360 113160 678600
rect 113400 678360 113490 678600
rect 113730 678360 113840 678600
rect 114080 678360 114170 678600
rect 114410 678360 114500 678600
rect 114740 678360 114830 678600
rect 115070 678360 115180 678600
rect 115420 678360 115510 678600
rect 115750 678360 115840 678600
rect 116080 678360 116170 678600
rect 116410 678360 116520 678600
rect 116760 678360 116850 678600
rect 117090 678360 117180 678600
rect 117420 678360 117510 678600
rect 117750 678360 117860 678600
rect 118100 678360 118190 678600
rect 118430 678360 118520 678600
rect 118760 678360 118850 678600
rect 119090 678360 119200 678600
rect 119440 678360 119530 678600
rect 119770 678360 119860 678600
rect 120100 678360 120190 678600
rect 120430 678360 120540 678600
rect 120780 678360 120870 678600
rect 121110 678360 121200 678600
rect 121440 678360 121530 678600
rect 121770 678360 122190 678600
rect 122430 678360 122540 678600
rect 122780 678360 122870 678600
rect 123110 678360 123200 678600
rect 123440 678360 123530 678600
rect 123770 678360 123880 678600
rect 124120 678360 124210 678600
rect 124450 678360 124540 678600
rect 124780 678360 124870 678600
rect 125110 678360 125220 678600
rect 125460 678360 125550 678600
rect 125790 678360 125880 678600
rect 126120 678360 126210 678600
rect 126450 678360 126560 678600
rect 126800 678360 126890 678600
rect 127130 678360 127220 678600
rect 127460 678360 127550 678600
rect 127790 678360 127900 678600
rect 128140 678360 128230 678600
rect 128470 678360 128560 678600
rect 128800 678360 128890 678600
rect 129130 678360 129240 678600
rect 129480 678360 129570 678600
rect 129810 678360 129900 678600
rect 130140 678360 130230 678600
rect 130470 678360 130580 678600
rect 130820 678360 130910 678600
rect 131150 678360 131240 678600
rect 131480 678360 131570 678600
rect 131810 678360 131920 678600
rect 132160 678360 132250 678600
rect 132490 678360 132580 678600
rect 132820 678360 132910 678600
rect 133150 678360 133570 678600
rect 133810 678360 133920 678600
rect 134160 678360 134250 678600
rect 134490 678360 134580 678600
rect 134820 678360 134910 678600
rect 135150 678360 135260 678600
rect 135500 678360 135590 678600
rect 135830 678360 135920 678600
rect 136160 678360 136250 678600
rect 136490 678360 136600 678600
rect 136840 678360 136930 678600
rect 137170 678360 137260 678600
rect 137500 678360 137590 678600
rect 137830 678360 137940 678600
rect 138180 678360 138270 678600
rect 138510 678360 138600 678600
rect 138840 678360 138930 678600
rect 139170 678360 139280 678600
rect 139520 678360 139610 678600
rect 139850 678360 139940 678600
rect 140180 678360 140270 678600
rect 140510 678360 140620 678600
rect 140860 678360 140950 678600
rect 141190 678360 141280 678600
rect 141520 678360 141610 678600
rect 141850 678360 141960 678600
rect 142200 678360 142290 678600
rect 142530 678360 142620 678600
rect 142860 678360 142950 678600
rect 143190 678360 143300 678600
rect 143540 678360 143630 678600
rect 143870 678360 143960 678600
rect 144200 678360 144290 678600
rect 144530 678360 144950 678600
rect 145190 678360 145300 678600
rect 145540 678360 145630 678600
rect 145870 678360 145960 678600
rect 146200 678360 146290 678600
rect 146530 678360 146640 678600
rect 146880 678360 146970 678600
rect 147210 678360 147300 678600
rect 147540 678360 147630 678600
rect 147870 678360 147980 678600
rect 148220 678360 148310 678600
rect 148550 678360 148640 678600
rect 148880 678360 148970 678600
rect 149210 678360 149320 678600
rect 149560 678360 149650 678600
rect 149890 678360 149980 678600
rect 150220 678360 150310 678600
rect 150550 678360 150660 678600
rect 150900 678360 150990 678600
rect 151230 678360 151320 678600
rect 151560 678360 151650 678600
rect 151890 678360 152000 678600
rect 152240 678360 152330 678600
rect 152570 678360 152660 678600
rect 152900 678360 152990 678600
rect 153230 678360 153340 678600
rect 153580 678360 153670 678600
rect 153910 678360 154000 678600
rect 154240 678360 154330 678600
rect 154570 678360 154680 678600
rect 154920 678360 155010 678600
rect 155250 678360 155340 678600
rect 155580 678360 155670 678600
rect 155910 678399 157520 678600
rect 157780 678399 157880 678639
rect 158140 678399 158240 678639
rect 158500 678399 158600 678639
rect 158860 678399 162436 678639
rect 155910 678360 162436 678399
rect 103643 678300 162436 678360
rect 103643 678060 107220 678300
rect 107480 678060 107580 678300
rect 107840 678060 107940 678300
rect 108200 678060 108300 678300
rect 108560 678299 162436 678300
rect 108560 678270 157520 678299
rect 108560 678060 110810 678270
rect 103643 678030 110810 678060
rect 111050 678030 111160 678270
rect 111400 678030 111490 678270
rect 111730 678030 111820 678270
rect 112060 678030 112150 678270
rect 112390 678030 112500 678270
rect 112740 678030 112830 678270
rect 113070 678030 113160 678270
rect 113400 678030 113490 678270
rect 113730 678030 113840 678270
rect 114080 678030 114170 678270
rect 114410 678030 114500 678270
rect 114740 678030 114830 678270
rect 115070 678030 115180 678270
rect 115420 678030 115510 678270
rect 115750 678030 115840 678270
rect 116080 678030 116170 678270
rect 116410 678030 116520 678270
rect 116760 678030 116850 678270
rect 117090 678030 117180 678270
rect 117420 678030 117510 678270
rect 117750 678030 117860 678270
rect 118100 678030 118190 678270
rect 118430 678030 118520 678270
rect 118760 678030 118850 678270
rect 119090 678030 119200 678270
rect 119440 678030 119530 678270
rect 119770 678030 119860 678270
rect 120100 678030 120190 678270
rect 120430 678030 120540 678270
rect 120780 678030 120870 678270
rect 121110 678030 121200 678270
rect 121440 678030 121530 678270
rect 121770 678030 122190 678270
rect 122430 678030 122540 678270
rect 122780 678030 122870 678270
rect 123110 678030 123200 678270
rect 123440 678030 123530 678270
rect 123770 678030 123880 678270
rect 124120 678030 124210 678270
rect 124450 678030 124540 678270
rect 124780 678030 124870 678270
rect 125110 678030 125220 678270
rect 125460 678030 125550 678270
rect 125790 678030 125880 678270
rect 126120 678030 126210 678270
rect 126450 678030 126560 678270
rect 126800 678030 126890 678270
rect 127130 678030 127220 678270
rect 127460 678030 127550 678270
rect 127790 678030 127900 678270
rect 128140 678030 128230 678270
rect 128470 678030 128560 678270
rect 128800 678030 128890 678270
rect 129130 678030 129240 678270
rect 129480 678030 129570 678270
rect 129810 678030 129900 678270
rect 130140 678030 130230 678270
rect 130470 678030 130580 678270
rect 130820 678030 130910 678270
rect 131150 678030 131240 678270
rect 131480 678030 131570 678270
rect 131810 678030 131920 678270
rect 132160 678030 132250 678270
rect 132490 678030 132580 678270
rect 132820 678030 132910 678270
rect 133150 678030 133570 678270
rect 133810 678030 133920 678270
rect 134160 678030 134250 678270
rect 134490 678030 134580 678270
rect 134820 678030 134910 678270
rect 135150 678030 135260 678270
rect 135500 678030 135590 678270
rect 135830 678030 135920 678270
rect 136160 678030 136250 678270
rect 136490 678030 136600 678270
rect 136840 678030 136930 678270
rect 137170 678030 137260 678270
rect 137500 678030 137590 678270
rect 137830 678030 137940 678270
rect 138180 678030 138270 678270
rect 138510 678030 138600 678270
rect 138840 678030 138930 678270
rect 139170 678030 139280 678270
rect 139520 678030 139610 678270
rect 139850 678030 139940 678270
rect 140180 678030 140270 678270
rect 140510 678030 140620 678270
rect 140860 678030 140950 678270
rect 141190 678030 141280 678270
rect 141520 678030 141610 678270
rect 141850 678030 141960 678270
rect 142200 678030 142290 678270
rect 142530 678030 142620 678270
rect 142860 678030 142950 678270
rect 143190 678030 143300 678270
rect 143540 678030 143630 678270
rect 143870 678030 143960 678270
rect 144200 678030 144290 678270
rect 144530 678030 144950 678270
rect 145190 678030 145300 678270
rect 145540 678030 145630 678270
rect 145870 678030 145960 678270
rect 146200 678030 146290 678270
rect 146530 678030 146640 678270
rect 146880 678030 146970 678270
rect 147210 678030 147300 678270
rect 147540 678030 147630 678270
rect 147870 678030 147980 678270
rect 148220 678030 148310 678270
rect 148550 678030 148640 678270
rect 148880 678030 148970 678270
rect 149210 678030 149320 678270
rect 149560 678030 149650 678270
rect 149890 678030 149980 678270
rect 150220 678030 150310 678270
rect 150550 678030 150660 678270
rect 150900 678030 150990 678270
rect 151230 678030 151320 678270
rect 151560 678030 151650 678270
rect 151890 678030 152000 678270
rect 152240 678030 152330 678270
rect 152570 678030 152660 678270
rect 152900 678030 152990 678270
rect 153230 678030 153340 678270
rect 153580 678030 153670 678270
rect 153910 678030 154000 678270
rect 154240 678030 154330 678270
rect 154570 678030 154680 678270
rect 154920 678030 155010 678270
rect 155250 678030 155340 678270
rect 155580 678030 155670 678270
rect 155910 678059 157520 678270
rect 157780 678059 157880 678299
rect 158140 678059 158240 678299
rect 158500 678059 158600 678299
rect 158860 678059 162436 678299
rect 155910 678030 162436 678059
rect 103643 677960 162436 678030
rect 103643 677720 107220 677960
rect 107480 677720 107580 677960
rect 107840 677720 107940 677960
rect 108200 677720 108300 677960
rect 108560 677959 162436 677960
rect 108560 677920 157520 677959
rect 108560 677720 110810 677920
rect 103643 677680 110810 677720
rect 111050 677680 111160 677920
rect 111400 677680 111490 677920
rect 111730 677680 111820 677920
rect 112060 677680 112150 677920
rect 112390 677680 112500 677920
rect 112740 677680 112830 677920
rect 113070 677680 113160 677920
rect 113400 677680 113490 677920
rect 113730 677680 113840 677920
rect 114080 677680 114170 677920
rect 114410 677680 114500 677920
rect 114740 677680 114830 677920
rect 115070 677680 115180 677920
rect 115420 677680 115510 677920
rect 115750 677680 115840 677920
rect 116080 677680 116170 677920
rect 116410 677680 116520 677920
rect 116760 677680 116850 677920
rect 117090 677680 117180 677920
rect 117420 677680 117510 677920
rect 117750 677680 117860 677920
rect 118100 677680 118190 677920
rect 118430 677680 118520 677920
rect 118760 677680 118850 677920
rect 119090 677680 119200 677920
rect 119440 677680 119530 677920
rect 119770 677680 119860 677920
rect 120100 677680 120190 677920
rect 120430 677680 120540 677920
rect 120780 677680 120870 677920
rect 121110 677680 121200 677920
rect 121440 677680 121530 677920
rect 121770 677680 122190 677920
rect 122430 677680 122540 677920
rect 122780 677680 122870 677920
rect 123110 677680 123200 677920
rect 123440 677680 123530 677920
rect 123770 677680 123880 677920
rect 124120 677680 124210 677920
rect 124450 677680 124540 677920
rect 124780 677680 124870 677920
rect 125110 677680 125220 677920
rect 125460 677680 125550 677920
rect 125790 677680 125880 677920
rect 126120 677680 126210 677920
rect 126450 677680 126560 677920
rect 126800 677680 126890 677920
rect 127130 677680 127220 677920
rect 127460 677680 127550 677920
rect 127790 677680 127900 677920
rect 128140 677680 128230 677920
rect 128470 677680 128560 677920
rect 128800 677680 128890 677920
rect 129130 677680 129240 677920
rect 129480 677680 129570 677920
rect 129810 677680 129900 677920
rect 130140 677680 130230 677920
rect 130470 677680 130580 677920
rect 130820 677680 130910 677920
rect 131150 677680 131240 677920
rect 131480 677680 131570 677920
rect 131810 677680 131920 677920
rect 132160 677680 132250 677920
rect 132490 677680 132580 677920
rect 132820 677680 132910 677920
rect 133150 677680 133570 677920
rect 133810 677680 133920 677920
rect 134160 677680 134250 677920
rect 134490 677680 134580 677920
rect 134820 677680 134910 677920
rect 135150 677680 135260 677920
rect 135500 677680 135590 677920
rect 135830 677680 135920 677920
rect 136160 677680 136250 677920
rect 136490 677680 136600 677920
rect 136840 677680 136930 677920
rect 137170 677680 137260 677920
rect 137500 677680 137590 677920
rect 137830 677680 137940 677920
rect 138180 677680 138270 677920
rect 138510 677680 138600 677920
rect 138840 677680 138930 677920
rect 139170 677680 139280 677920
rect 139520 677680 139610 677920
rect 139850 677680 139940 677920
rect 140180 677680 140270 677920
rect 140510 677680 140620 677920
rect 140860 677680 140950 677920
rect 141190 677680 141280 677920
rect 141520 677680 141610 677920
rect 141850 677680 141960 677920
rect 142200 677680 142290 677920
rect 142530 677680 142620 677920
rect 142860 677680 142950 677920
rect 143190 677680 143300 677920
rect 143540 677680 143630 677920
rect 143870 677680 143960 677920
rect 144200 677680 144290 677920
rect 144530 677680 144950 677920
rect 145190 677680 145300 677920
rect 145540 677680 145630 677920
rect 145870 677680 145960 677920
rect 146200 677680 146290 677920
rect 146530 677680 146640 677920
rect 146880 677680 146970 677920
rect 147210 677680 147300 677920
rect 147540 677680 147630 677920
rect 147870 677680 147980 677920
rect 148220 677680 148310 677920
rect 148550 677680 148640 677920
rect 148880 677680 148970 677920
rect 149210 677680 149320 677920
rect 149560 677680 149650 677920
rect 149890 677680 149980 677920
rect 150220 677680 150310 677920
rect 150550 677680 150660 677920
rect 150900 677680 150990 677920
rect 151230 677680 151320 677920
rect 151560 677680 151650 677920
rect 151890 677680 152000 677920
rect 152240 677680 152330 677920
rect 152570 677680 152660 677920
rect 152900 677680 152990 677920
rect 153230 677680 153340 677920
rect 153580 677680 153670 677920
rect 153910 677680 154000 677920
rect 154240 677680 154330 677920
rect 154570 677680 154680 677920
rect 154920 677680 155010 677920
rect 155250 677680 155340 677920
rect 155580 677680 155670 677920
rect 155910 677719 157520 677920
rect 157780 677719 157880 677959
rect 158140 677719 158240 677959
rect 158500 677719 158600 677959
rect 158860 677719 162436 677959
rect 155910 677680 162436 677719
rect 103643 677620 162436 677680
rect 103643 677380 107220 677620
rect 107480 677380 107580 677620
rect 107840 677380 107940 677620
rect 108200 677380 108300 677620
rect 108560 677619 162436 677620
rect 108560 677590 157520 677619
rect 108560 677380 110810 677590
rect 103643 677350 110810 677380
rect 111050 677350 111160 677590
rect 111400 677350 111490 677590
rect 111730 677350 111820 677590
rect 112060 677350 112150 677590
rect 112390 677350 112500 677590
rect 112740 677350 112830 677590
rect 113070 677350 113160 677590
rect 113400 677350 113490 677590
rect 113730 677350 113840 677590
rect 114080 677350 114170 677590
rect 114410 677350 114500 677590
rect 114740 677350 114830 677590
rect 115070 677350 115180 677590
rect 115420 677350 115510 677590
rect 115750 677350 115840 677590
rect 116080 677350 116170 677590
rect 116410 677350 116520 677590
rect 116760 677350 116850 677590
rect 117090 677350 117180 677590
rect 117420 677350 117510 677590
rect 117750 677350 117860 677590
rect 118100 677350 118190 677590
rect 118430 677350 118520 677590
rect 118760 677350 118850 677590
rect 119090 677350 119200 677590
rect 119440 677350 119530 677590
rect 119770 677350 119860 677590
rect 120100 677350 120190 677590
rect 120430 677350 120540 677590
rect 120780 677350 120870 677590
rect 121110 677350 121200 677590
rect 121440 677350 121530 677590
rect 121770 677350 122190 677590
rect 122430 677350 122540 677590
rect 122780 677350 122870 677590
rect 123110 677350 123200 677590
rect 123440 677350 123530 677590
rect 123770 677350 123880 677590
rect 124120 677350 124210 677590
rect 124450 677350 124540 677590
rect 124780 677350 124870 677590
rect 125110 677350 125220 677590
rect 125460 677350 125550 677590
rect 125790 677350 125880 677590
rect 126120 677350 126210 677590
rect 126450 677350 126560 677590
rect 126800 677350 126890 677590
rect 127130 677350 127220 677590
rect 127460 677350 127550 677590
rect 127790 677350 127900 677590
rect 128140 677350 128230 677590
rect 128470 677350 128560 677590
rect 128800 677350 128890 677590
rect 129130 677350 129240 677590
rect 129480 677350 129570 677590
rect 129810 677350 129900 677590
rect 130140 677350 130230 677590
rect 130470 677350 130580 677590
rect 130820 677350 130910 677590
rect 131150 677350 131240 677590
rect 131480 677350 131570 677590
rect 131810 677350 131920 677590
rect 132160 677350 132250 677590
rect 132490 677350 132580 677590
rect 132820 677350 132910 677590
rect 133150 677350 133570 677590
rect 133810 677350 133920 677590
rect 134160 677350 134250 677590
rect 134490 677350 134580 677590
rect 134820 677350 134910 677590
rect 135150 677350 135260 677590
rect 135500 677350 135590 677590
rect 135830 677350 135920 677590
rect 136160 677350 136250 677590
rect 136490 677350 136600 677590
rect 136840 677350 136930 677590
rect 137170 677350 137260 677590
rect 137500 677350 137590 677590
rect 137830 677350 137940 677590
rect 138180 677350 138270 677590
rect 138510 677350 138600 677590
rect 138840 677350 138930 677590
rect 139170 677350 139280 677590
rect 139520 677350 139610 677590
rect 139850 677350 139940 677590
rect 140180 677350 140270 677590
rect 140510 677350 140620 677590
rect 140860 677350 140950 677590
rect 141190 677350 141280 677590
rect 141520 677350 141610 677590
rect 141850 677350 141960 677590
rect 142200 677350 142290 677590
rect 142530 677350 142620 677590
rect 142860 677350 142950 677590
rect 143190 677350 143300 677590
rect 143540 677350 143630 677590
rect 143870 677350 143960 677590
rect 144200 677350 144290 677590
rect 144530 677350 144950 677590
rect 145190 677350 145300 677590
rect 145540 677350 145630 677590
rect 145870 677350 145960 677590
rect 146200 677350 146290 677590
rect 146530 677350 146640 677590
rect 146880 677350 146970 677590
rect 147210 677350 147300 677590
rect 147540 677350 147630 677590
rect 147870 677350 147980 677590
rect 148220 677350 148310 677590
rect 148550 677350 148640 677590
rect 148880 677350 148970 677590
rect 149210 677350 149320 677590
rect 149560 677350 149650 677590
rect 149890 677350 149980 677590
rect 150220 677350 150310 677590
rect 150550 677350 150660 677590
rect 150900 677350 150990 677590
rect 151230 677350 151320 677590
rect 151560 677350 151650 677590
rect 151890 677350 152000 677590
rect 152240 677350 152330 677590
rect 152570 677350 152660 677590
rect 152900 677350 152990 677590
rect 153230 677350 153340 677590
rect 153580 677350 153670 677590
rect 153910 677350 154000 677590
rect 154240 677350 154330 677590
rect 154570 677350 154680 677590
rect 154920 677350 155010 677590
rect 155250 677350 155340 677590
rect 155580 677350 155670 677590
rect 155910 677379 157520 677590
rect 157780 677379 157880 677619
rect 158140 677379 158240 677619
rect 158500 677379 158600 677619
rect 158860 677379 162436 677619
rect 155910 677350 162436 677379
rect 103643 677280 162436 677350
rect 103643 677040 107220 677280
rect 107480 677040 107580 677280
rect 107840 677040 107940 677280
rect 108200 677040 108300 677280
rect 108560 677279 162436 677280
rect 108560 677260 157520 677279
rect 108560 677040 110810 677260
rect 103643 677020 110810 677040
rect 111050 677020 111160 677260
rect 111400 677020 111490 677260
rect 111730 677020 111820 677260
rect 112060 677020 112150 677260
rect 112390 677020 112500 677260
rect 112740 677020 112830 677260
rect 113070 677020 113160 677260
rect 113400 677020 113490 677260
rect 113730 677020 113840 677260
rect 114080 677020 114170 677260
rect 114410 677020 114500 677260
rect 114740 677020 114830 677260
rect 115070 677020 115180 677260
rect 115420 677020 115510 677260
rect 115750 677020 115840 677260
rect 116080 677020 116170 677260
rect 116410 677020 116520 677260
rect 116760 677020 116850 677260
rect 117090 677020 117180 677260
rect 117420 677020 117510 677260
rect 117750 677020 117860 677260
rect 118100 677020 118190 677260
rect 118430 677020 118520 677260
rect 118760 677020 118850 677260
rect 119090 677020 119200 677260
rect 119440 677020 119530 677260
rect 119770 677020 119860 677260
rect 120100 677020 120190 677260
rect 120430 677020 120540 677260
rect 120780 677020 120870 677260
rect 121110 677020 121200 677260
rect 121440 677020 121530 677260
rect 121770 677020 122190 677260
rect 122430 677020 122540 677260
rect 122780 677020 122870 677260
rect 123110 677020 123200 677260
rect 123440 677020 123530 677260
rect 123770 677020 123880 677260
rect 124120 677020 124210 677260
rect 124450 677020 124540 677260
rect 124780 677020 124870 677260
rect 125110 677020 125220 677260
rect 125460 677020 125550 677260
rect 125790 677020 125880 677260
rect 126120 677020 126210 677260
rect 126450 677020 126560 677260
rect 126800 677020 126890 677260
rect 127130 677020 127220 677260
rect 127460 677020 127550 677260
rect 127790 677020 127900 677260
rect 128140 677020 128230 677260
rect 128470 677020 128560 677260
rect 128800 677020 128890 677260
rect 129130 677020 129240 677260
rect 129480 677020 129570 677260
rect 129810 677020 129900 677260
rect 130140 677020 130230 677260
rect 130470 677020 130580 677260
rect 130820 677020 130910 677260
rect 131150 677020 131240 677260
rect 131480 677020 131570 677260
rect 131810 677020 131920 677260
rect 132160 677020 132250 677260
rect 132490 677020 132580 677260
rect 132820 677020 132910 677260
rect 133150 677020 133570 677260
rect 133810 677020 133920 677260
rect 134160 677020 134250 677260
rect 134490 677020 134580 677260
rect 134820 677020 134910 677260
rect 135150 677020 135260 677260
rect 135500 677020 135590 677260
rect 135830 677020 135920 677260
rect 136160 677020 136250 677260
rect 136490 677020 136600 677260
rect 136840 677020 136930 677260
rect 137170 677020 137260 677260
rect 137500 677020 137590 677260
rect 137830 677020 137940 677260
rect 138180 677020 138270 677260
rect 138510 677020 138600 677260
rect 138840 677020 138930 677260
rect 139170 677020 139280 677260
rect 139520 677020 139610 677260
rect 139850 677020 139940 677260
rect 140180 677020 140270 677260
rect 140510 677020 140620 677260
rect 140860 677020 140950 677260
rect 141190 677020 141280 677260
rect 141520 677020 141610 677260
rect 141850 677020 141960 677260
rect 142200 677020 142290 677260
rect 142530 677020 142620 677260
rect 142860 677020 142950 677260
rect 143190 677020 143300 677260
rect 143540 677020 143630 677260
rect 143870 677020 143960 677260
rect 144200 677020 144290 677260
rect 144530 677020 144950 677260
rect 145190 677020 145300 677260
rect 145540 677020 145630 677260
rect 145870 677020 145960 677260
rect 146200 677020 146290 677260
rect 146530 677020 146640 677260
rect 146880 677020 146970 677260
rect 147210 677020 147300 677260
rect 147540 677020 147630 677260
rect 147870 677020 147980 677260
rect 148220 677020 148310 677260
rect 148550 677020 148640 677260
rect 148880 677020 148970 677260
rect 149210 677020 149320 677260
rect 149560 677020 149650 677260
rect 149890 677020 149980 677260
rect 150220 677020 150310 677260
rect 150550 677020 150660 677260
rect 150900 677020 150990 677260
rect 151230 677020 151320 677260
rect 151560 677020 151650 677260
rect 151890 677020 152000 677260
rect 152240 677020 152330 677260
rect 152570 677020 152660 677260
rect 152900 677020 152990 677260
rect 153230 677020 153340 677260
rect 153580 677020 153670 677260
rect 153910 677020 154000 677260
rect 154240 677020 154330 677260
rect 154570 677020 154680 677260
rect 154920 677020 155010 677260
rect 155250 677020 155340 677260
rect 155580 677020 155670 677260
rect 155910 677039 157520 677260
rect 157780 677039 157880 677279
rect 158140 677039 158240 677279
rect 158500 677039 158600 677279
rect 158860 677039 162436 677279
rect 155910 677020 162436 677039
rect 103643 676940 162436 677020
rect 103643 676700 107220 676940
rect 107480 676700 107580 676940
rect 107840 676700 107940 676940
rect 108200 676700 108300 676940
rect 108560 676939 162436 676940
rect 108560 676930 157520 676939
rect 108560 676700 110810 676930
rect 103643 676690 110810 676700
rect 111050 676690 111160 676930
rect 111400 676690 111490 676930
rect 111730 676690 111820 676930
rect 112060 676690 112150 676930
rect 112390 676690 112500 676930
rect 112740 676690 112830 676930
rect 113070 676690 113160 676930
rect 113400 676690 113490 676930
rect 113730 676690 113840 676930
rect 114080 676690 114170 676930
rect 114410 676690 114500 676930
rect 114740 676690 114830 676930
rect 115070 676690 115180 676930
rect 115420 676690 115510 676930
rect 115750 676690 115840 676930
rect 116080 676690 116170 676930
rect 116410 676690 116520 676930
rect 116760 676690 116850 676930
rect 117090 676690 117180 676930
rect 117420 676690 117510 676930
rect 117750 676690 117860 676930
rect 118100 676690 118190 676930
rect 118430 676690 118520 676930
rect 118760 676690 118850 676930
rect 119090 676690 119200 676930
rect 119440 676690 119530 676930
rect 119770 676690 119860 676930
rect 120100 676690 120190 676930
rect 120430 676690 120540 676930
rect 120780 676690 120870 676930
rect 121110 676690 121200 676930
rect 121440 676690 121530 676930
rect 121770 676690 122190 676930
rect 122430 676690 122540 676930
rect 122780 676690 122870 676930
rect 123110 676690 123200 676930
rect 123440 676690 123530 676930
rect 123770 676690 123880 676930
rect 124120 676690 124210 676930
rect 124450 676690 124540 676930
rect 124780 676690 124870 676930
rect 125110 676690 125220 676930
rect 125460 676690 125550 676930
rect 125790 676690 125880 676930
rect 126120 676690 126210 676930
rect 126450 676690 126560 676930
rect 126800 676690 126890 676930
rect 127130 676690 127220 676930
rect 127460 676690 127550 676930
rect 127790 676690 127900 676930
rect 128140 676690 128230 676930
rect 128470 676690 128560 676930
rect 128800 676690 128890 676930
rect 129130 676690 129240 676930
rect 129480 676690 129570 676930
rect 129810 676690 129900 676930
rect 130140 676690 130230 676930
rect 130470 676690 130580 676930
rect 130820 676690 130910 676930
rect 131150 676690 131240 676930
rect 131480 676690 131570 676930
rect 131810 676690 131920 676930
rect 132160 676690 132250 676930
rect 132490 676690 132580 676930
rect 132820 676690 132910 676930
rect 133150 676690 133570 676930
rect 133810 676690 133920 676930
rect 134160 676690 134250 676930
rect 134490 676690 134580 676930
rect 134820 676690 134910 676930
rect 135150 676690 135260 676930
rect 135500 676690 135590 676930
rect 135830 676690 135920 676930
rect 136160 676690 136250 676930
rect 136490 676690 136600 676930
rect 136840 676690 136930 676930
rect 137170 676690 137260 676930
rect 137500 676690 137590 676930
rect 137830 676690 137940 676930
rect 138180 676690 138270 676930
rect 138510 676690 138600 676930
rect 138840 676690 138930 676930
rect 139170 676690 139280 676930
rect 139520 676690 139610 676930
rect 139850 676690 139940 676930
rect 140180 676690 140270 676930
rect 140510 676690 140620 676930
rect 140860 676690 140950 676930
rect 141190 676690 141280 676930
rect 141520 676690 141610 676930
rect 141850 676690 141960 676930
rect 142200 676690 142290 676930
rect 142530 676690 142620 676930
rect 142860 676690 142950 676930
rect 143190 676690 143300 676930
rect 143540 676690 143630 676930
rect 143870 676690 143960 676930
rect 144200 676690 144290 676930
rect 144530 676690 144950 676930
rect 145190 676690 145300 676930
rect 145540 676690 145630 676930
rect 145870 676690 145960 676930
rect 146200 676690 146290 676930
rect 146530 676690 146640 676930
rect 146880 676690 146970 676930
rect 147210 676690 147300 676930
rect 147540 676690 147630 676930
rect 147870 676690 147980 676930
rect 148220 676690 148310 676930
rect 148550 676690 148640 676930
rect 148880 676690 148970 676930
rect 149210 676690 149320 676930
rect 149560 676690 149650 676930
rect 149890 676690 149980 676930
rect 150220 676690 150310 676930
rect 150550 676690 150660 676930
rect 150900 676690 150990 676930
rect 151230 676690 151320 676930
rect 151560 676690 151650 676930
rect 151890 676690 152000 676930
rect 152240 676690 152330 676930
rect 152570 676690 152660 676930
rect 152900 676690 152990 676930
rect 153230 676690 153340 676930
rect 153580 676690 153670 676930
rect 153910 676690 154000 676930
rect 154240 676690 154330 676930
rect 154570 676690 154680 676930
rect 154920 676690 155010 676930
rect 155250 676690 155340 676930
rect 155580 676690 155670 676930
rect 155910 676699 157520 676930
rect 157780 676699 157880 676939
rect 158140 676699 158240 676939
rect 158500 676699 158600 676939
rect 158860 676699 162436 676939
rect 155910 676690 162436 676699
rect 103643 676600 162436 676690
rect 103643 676360 107220 676600
rect 107480 676360 107580 676600
rect 107840 676360 107940 676600
rect 108200 676360 108300 676600
rect 108560 676599 162436 676600
rect 108560 676580 157520 676599
rect 108560 676360 110810 676580
rect 103643 676340 110810 676360
rect 111050 676340 111160 676580
rect 111400 676340 111490 676580
rect 111730 676340 111820 676580
rect 112060 676340 112150 676580
rect 112390 676340 112500 676580
rect 112740 676340 112830 676580
rect 113070 676340 113160 676580
rect 113400 676340 113490 676580
rect 113730 676340 113840 676580
rect 114080 676340 114170 676580
rect 114410 676340 114500 676580
rect 114740 676340 114830 676580
rect 115070 676340 115180 676580
rect 115420 676340 115510 676580
rect 115750 676340 115840 676580
rect 116080 676340 116170 676580
rect 116410 676340 116520 676580
rect 116760 676340 116850 676580
rect 117090 676340 117180 676580
rect 117420 676340 117510 676580
rect 117750 676340 117860 676580
rect 118100 676340 118190 676580
rect 118430 676340 118520 676580
rect 118760 676340 118850 676580
rect 119090 676340 119200 676580
rect 119440 676340 119530 676580
rect 119770 676340 119860 676580
rect 120100 676340 120190 676580
rect 120430 676340 120540 676580
rect 120780 676340 120870 676580
rect 121110 676340 121200 676580
rect 121440 676340 121530 676580
rect 121770 676340 122190 676580
rect 122430 676340 122540 676580
rect 122780 676340 122870 676580
rect 123110 676340 123200 676580
rect 123440 676340 123530 676580
rect 123770 676340 123880 676580
rect 124120 676340 124210 676580
rect 124450 676340 124540 676580
rect 124780 676340 124870 676580
rect 125110 676340 125220 676580
rect 125460 676340 125550 676580
rect 125790 676340 125880 676580
rect 126120 676340 126210 676580
rect 126450 676340 126560 676580
rect 126800 676340 126890 676580
rect 127130 676340 127220 676580
rect 127460 676340 127550 676580
rect 127790 676340 127900 676580
rect 128140 676340 128230 676580
rect 128470 676340 128560 676580
rect 128800 676340 128890 676580
rect 129130 676340 129240 676580
rect 129480 676340 129570 676580
rect 129810 676340 129900 676580
rect 130140 676340 130230 676580
rect 130470 676340 130580 676580
rect 130820 676340 130910 676580
rect 131150 676340 131240 676580
rect 131480 676340 131570 676580
rect 131810 676340 131920 676580
rect 132160 676340 132250 676580
rect 132490 676340 132580 676580
rect 132820 676340 132910 676580
rect 133150 676340 133570 676580
rect 133810 676340 133920 676580
rect 134160 676340 134250 676580
rect 134490 676340 134580 676580
rect 134820 676340 134910 676580
rect 135150 676340 135260 676580
rect 135500 676340 135590 676580
rect 135830 676340 135920 676580
rect 136160 676340 136250 676580
rect 136490 676340 136600 676580
rect 136840 676340 136930 676580
rect 137170 676340 137260 676580
rect 137500 676340 137590 676580
rect 137830 676340 137940 676580
rect 138180 676340 138270 676580
rect 138510 676340 138600 676580
rect 138840 676340 138930 676580
rect 139170 676340 139280 676580
rect 139520 676340 139610 676580
rect 139850 676340 139940 676580
rect 140180 676340 140270 676580
rect 140510 676340 140620 676580
rect 140860 676340 140950 676580
rect 141190 676340 141280 676580
rect 141520 676340 141610 676580
rect 141850 676340 141960 676580
rect 142200 676340 142290 676580
rect 142530 676340 142620 676580
rect 142860 676340 142950 676580
rect 143190 676340 143300 676580
rect 143540 676340 143630 676580
rect 143870 676340 143960 676580
rect 144200 676340 144290 676580
rect 144530 676340 144950 676580
rect 145190 676340 145300 676580
rect 145540 676340 145630 676580
rect 145870 676340 145960 676580
rect 146200 676340 146290 676580
rect 146530 676340 146640 676580
rect 146880 676340 146970 676580
rect 147210 676340 147300 676580
rect 147540 676340 147630 676580
rect 147870 676340 147980 676580
rect 148220 676340 148310 676580
rect 148550 676340 148640 676580
rect 148880 676340 148970 676580
rect 149210 676340 149320 676580
rect 149560 676340 149650 676580
rect 149890 676340 149980 676580
rect 150220 676340 150310 676580
rect 150550 676340 150660 676580
rect 150900 676340 150990 676580
rect 151230 676340 151320 676580
rect 151560 676340 151650 676580
rect 151890 676340 152000 676580
rect 152240 676340 152330 676580
rect 152570 676340 152660 676580
rect 152900 676340 152990 676580
rect 153230 676340 153340 676580
rect 153580 676340 153670 676580
rect 153910 676340 154000 676580
rect 154240 676340 154330 676580
rect 154570 676340 154680 676580
rect 154920 676340 155010 676580
rect 155250 676340 155340 676580
rect 155580 676340 155670 676580
rect 155910 676359 157520 676580
rect 157780 676359 157880 676599
rect 158140 676359 158240 676599
rect 158500 676359 158600 676599
rect 158860 676359 162436 676599
rect 155910 676340 162436 676359
rect 103643 676260 162436 676340
rect 103643 676020 107220 676260
rect 107480 676020 107580 676260
rect 107840 676020 107940 676260
rect 108200 676020 108300 676260
rect 108560 676259 162436 676260
rect 108560 676250 157520 676259
rect 108560 676020 110810 676250
rect 103643 676010 110810 676020
rect 111050 676010 111160 676250
rect 111400 676010 111490 676250
rect 111730 676010 111820 676250
rect 112060 676010 112150 676250
rect 112390 676010 112500 676250
rect 112740 676010 112830 676250
rect 113070 676010 113160 676250
rect 113400 676010 113490 676250
rect 113730 676010 113840 676250
rect 114080 676010 114170 676250
rect 114410 676010 114500 676250
rect 114740 676010 114830 676250
rect 115070 676010 115180 676250
rect 115420 676010 115510 676250
rect 115750 676010 115840 676250
rect 116080 676010 116170 676250
rect 116410 676010 116520 676250
rect 116760 676010 116850 676250
rect 117090 676010 117180 676250
rect 117420 676010 117510 676250
rect 117750 676010 117860 676250
rect 118100 676010 118190 676250
rect 118430 676010 118520 676250
rect 118760 676010 118850 676250
rect 119090 676010 119200 676250
rect 119440 676010 119530 676250
rect 119770 676010 119860 676250
rect 120100 676010 120190 676250
rect 120430 676010 120540 676250
rect 120780 676010 120870 676250
rect 121110 676010 121200 676250
rect 121440 676010 121530 676250
rect 121770 676010 122190 676250
rect 122430 676010 122540 676250
rect 122780 676010 122870 676250
rect 123110 676010 123200 676250
rect 123440 676010 123530 676250
rect 123770 676010 123880 676250
rect 124120 676010 124210 676250
rect 124450 676010 124540 676250
rect 124780 676010 124870 676250
rect 125110 676010 125220 676250
rect 125460 676010 125550 676250
rect 125790 676010 125880 676250
rect 126120 676010 126210 676250
rect 126450 676010 126560 676250
rect 126800 676010 126890 676250
rect 127130 676010 127220 676250
rect 127460 676010 127550 676250
rect 127790 676010 127900 676250
rect 128140 676010 128230 676250
rect 128470 676010 128560 676250
rect 128800 676010 128890 676250
rect 129130 676010 129240 676250
rect 129480 676010 129570 676250
rect 129810 676010 129900 676250
rect 130140 676010 130230 676250
rect 130470 676010 130580 676250
rect 130820 676010 130910 676250
rect 131150 676010 131240 676250
rect 131480 676010 131570 676250
rect 131810 676010 131920 676250
rect 132160 676010 132250 676250
rect 132490 676010 132580 676250
rect 132820 676010 132910 676250
rect 133150 676010 133570 676250
rect 133810 676010 133920 676250
rect 134160 676010 134250 676250
rect 134490 676010 134580 676250
rect 134820 676010 134910 676250
rect 135150 676010 135260 676250
rect 135500 676010 135590 676250
rect 135830 676010 135920 676250
rect 136160 676010 136250 676250
rect 136490 676010 136600 676250
rect 136840 676010 136930 676250
rect 137170 676010 137260 676250
rect 137500 676010 137590 676250
rect 137830 676010 137940 676250
rect 138180 676010 138270 676250
rect 138510 676010 138600 676250
rect 138840 676010 138930 676250
rect 139170 676010 139280 676250
rect 139520 676010 139610 676250
rect 139850 676010 139940 676250
rect 140180 676010 140270 676250
rect 140510 676010 140620 676250
rect 140860 676010 140950 676250
rect 141190 676010 141280 676250
rect 141520 676010 141610 676250
rect 141850 676010 141960 676250
rect 142200 676010 142290 676250
rect 142530 676010 142620 676250
rect 142860 676010 142950 676250
rect 143190 676010 143300 676250
rect 143540 676010 143630 676250
rect 143870 676010 143960 676250
rect 144200 676010 144290 676250
rect 144530 676010 144950 676250
rect 145190 676010 145300 676250
rect 145540 676010 145630 676250
rect 145870 676010 145960 676250
rect 146200 676010 146290 676250
rect 146530 676010 146640 676250
rect 146880 676010 146970 676250
rect 147210 676010 147300 676250
rect 147540 676010 147630 676250
rect 147870 676010 147980 676250
rect 148220 676010 148310 676250
rect 148550 676010 148640 676250
rect 148880 676010 148970 676250
rect 149210 676010 149320 676250
rect 149560 676010 149650 676250
rect 149890 676010 149980 676250
rect 150220 676010 150310 676250
rect 150550 676010 150660 676250
rect 150900 676010 150990 676250
rect 151230 676010 151320 676250
rect 151560 676010 151650 676250
rect 151890 676010 152000 676250
rect 152240 676010 152330 676250
rect 152570 676010 152660 676250
rect 152900 676010 152990 676250
rect 153230 676010 153340 676250
rect 153580 676010 153670 676250
rect 153910 676010 154000 676250
rect 154240 676010 154330 676250
rect 154570 676010 154680 676250
rect 154920 676010 155010 676250
rect 155250 676010 155340 676250
rect 155580 676010 155670 676250
rect 155910 676019 157520 676250
rect 157780 676019 157880 676259
rect 158140 676019 158240 676259
rect 158500 676019 158600 676259
rect 158860 676019 162436 676259
rect 155910 676010 162436 676019
rect 103643 675920 162436 676010
rect 103643 675680 107220 675920
rect 107480 675680 107580 675920
rect 107840 675680 107940 675920
rect 108200 675680 108300 675920
rect 108560 675680 110810 675920
rect 111050 675680 111160 675920
rect 111400 675680 111490 675920
rect 111730 675680 111820 675920
rect 112060 675680 112150 675920
rect 112390 675680 112500 675920
rect 112740 675680 112830 675920
rect 113070 675680 113160 675920
rect 113400 675680 113490 675920
rect 113730 675680 113840 675920
rect 114080 675680 114170 675920
rect 114410 675680 114500 675920
rect 114740 675680 114830 675920
rect 115070 675680 115180 675920
rect 115420 675680 115510 675920
rect 115750 675680 115840 675920
rect 116080 675680 116170 675920
rect 116410 675680 116520 675920
rect 116760 675680 116850 675920
rect 117090 675680 117180 675920
rect 117420 675680 117510 675920
rect 117750 675680 117860 675920
rect 118100 675680 118190 675920
rect 118430 675680 118520 675920
rect 118760 675680 118850 675920
rect 119090 675680 119200 675920
rect 119440 675680 119530 675920
rect 119770 675680 119860 675920
rect 120100 675680 120190 675920
rect 120430 675680 120540 675920
rect 120780 675680 120870 675920
rect 121110 675680 121200 675920
rect 121440 675680 121530 675920
rect 121770 675680 122190 675920
rect 122430 675680 122540 675920
rect 122780 675680 122870 675920
rect 123110 675680 123200 675920
rect 123440 675680 123530 675920
rect 123770 675680 123880 675920
rect 124120 675680 124210 675920
rect 124450 675680 124540 675920
rect 124780 675680 124870 675920
rect 125110 675680 125220 675920
rect 125460 675680 125550 675920
rect 125790 675680 125880 675920
rect 126120 675680 126210 675920
rect 126450 675680 126560 675920
rect 126800 675680 126890 675920
rect 127130 675680 127220 675920
rect 127460 675680 127550 675920
rect 127790 675680 127900 675920
rect 128140 675680 128230 675920
rect 128470 675680 128560 675920
rect 128800 675680 128890 675920
rect 129130 675680 129240 675920
rect 129480 675680 129570 675920
rect 129810 675680 129900 675920
rect 130140 675680 130230 675920
rect 130470 675680 130580 675920
rect 130820 675680 130910 675920
rect 131150 675680 131240 675920
rect 131480 675680 131570 675920
rect 131810 675680 131920 675920
rect 132160 675680 132250 675920
rect 132490 675680 132580 675920
rect 132820 675680 132910 675920
rect 133150 675680 133570 675920
rect 133810 675680 133920 675920
rect 134160 675680 134250 675920
rect 134490 675680 134580 675920
rect 134820 675680 134910 675920
rect 135150 675680 135260 675920
rect 135500 675680 135590 675920
rect 135830 675680 135920 675920
rect 136160 675680 136250 675920
rect 136490 675680 136600 675920
rect 136840 675680 136930 675920
rect 137170 675680 137260 675920
rect 137500 675680 137590 675920
rect 137830 675680 137940 675920
rect 138180 675680 138270 675920
rect 138510 675680 138600 675920
rect 138840 675680 138930 675920
rect 139170 675680 139280 675920
rect 139520 675680 139610 675920
rect 139850 675680 139940 675920
rect 140180 675680 140270 675920
rect 140510 675680 140620 675920
rect 140860 675680 140950 675920
rect 141190 675680 141280 675920
rect 141520 675680 141610 675920
rect 141850 675680 141960 675920
rect 142200 675680 142290 675920
rect 142530 675680 142620 675920
rect 142860 675680 142950 675920
rect 143190 675680 143300 675920
rect 143540 675680 143630 675920
rect 143870 675680 143960 675920
rect 144200 675680 144290 675920
rect 144530 675680 144950 675920
rect 145190 675680 145300 675920
rect 145540 675680 145630 675920
rect 145870 675680 145960 675920
rect 146200 675680 146290 675920
rect 146530 675680 146640 675920
rect 146880 675680 146970 675920
rect 147210 675680 147300 675920
rect 147540 675680 147630 675920
rect 147870 675680 147980 675920
rect 148220 675680 148310 675920
rect 148550 675680 148640 675920
rect 148880 675680 148970 675920
rect 149210 675680 149320 675920
rect 149560 675680 149650 675920
rect 149890 675680 149980 675920
rect 150220 675680 150310 675920
rect 150550 675680 150660 675920
rect 150900 675680 150990 675920
rect 151230 675680 151320 675920
rect 151560 675680 151650 675920
rect 151890 675680 152000 675920
rect 152240 675680 152330 675920
rect 152570 675680 152660 675920
rect 152900 675680 152990 675920
rect 153230 675680 153340 675920
rect 153580 675680 153670 675920
rect 153910 675680 154000 675920
rect 154240 675680 154330 675920
rect 154570 675680 154680 675920
rect 154920 675680 155010 675920
rect 155250 675680 155340 675920
rect 155580 675680 155670 675920
rect 155910 675919 162436 675920
rect 155910 675680 157520 675919
rect 103643 675679 157520 675680
rect 157780 675679 157880 675919
rect 158140 675679 158240 675919
rect 158500 675679 158600 675919
rect 158860 675679 162436 675919
rect 103643 675590 162436 675679
rect 103643 675580 110810 675590
rect 103643 675340 107220 675580
rect 107480 675340 107580 675580
rect 107840 675340 107940 675580
rect 108200 675340 108300 675580
rect 108560 675350 110810 675580
rect 111050 675350 111160 675590
rect 111400 675350 111490 675590
rect 111730 675350 111820 675590
rect 112060 675350 112150 675590
rect 112390 675350 112500 675590
rect 112740 675350 112830 675590
rect 113070 675350 113160 675590
rect 113400 675350 113490 675590
rect 113730 675350 113840 675590
rect 114080 675350 114170 675590
rect 114410 675350 114500 675590
rect 114740 675350 114830 675590
rect 115070 675350 115180 675590
rect 115420 675350 115510 675590
rect 115750 675350 115840 675590
rect 116080 675350 116170 675590
rect 116410 675350 116520 675590
rect 116760 675350 116850 675590
rect 117090 675350 117180 675590
rect 117420 675350 117510 675590
rect 117750 675350 117860 675590
rect 118100 675350 118190 675590
rect 118430 675350 118520 675590
rect 118760 675350 118850 675590
rect 119090 675350 119200 675590
rect 119440 675350 119530 675590
rect 119770 675350 119860 675590
rect 120100 675350 120190 675590
rect 120430 675350 120540 675590
rect 120780 675350 120870 675590
rect 121110 675350 121200 675590
rect 121440 675350 121530 675590
rect 121770 675350 122190 675590
rect 122430 675350 122540 675590
rect 122780 675350 122870 675590
rect 123110 675350 123200 675590
rect 123440 675350 123530 675590
rect 123770 675350 123880 675590
rect 124120 675350 124210 675590
rect 124450 675350 124540 675590
rect 124780 675350 124870 675590
rect 125110 675350 125220 675590
rect 125460 675350 125550 675590
rect 125790 675350 125880 675590
rect 126120 675350 126210 675590
rect 126450 675350 126560 675590
rect 126800 675350 126890 675590
rect 127130 675350 127220 675590
rect 127460 675350 127550 675590
rect 127790 675350 127900 675590
rect 128140 675350 128230 675590
rect 128470 675350 128560 675590
rect 128800 675350 128890 675590
rect 129130 675350 129240 675590
rect 129480 675350 129570 675590
rect 129810 675350 129900 675590
rect 130140 675350 130230 675590
rect 130470 675350 130580 675590
rect 130820 675350 130910 675590
rect 131150 675350 131240 675590
rect 131480 675350 131570 675590
rect 131810 675350 131920 675590
rect 132160 675350 132250 675590
rect 132490 675350 132580 675590
rect 132820 675350 132910 675590
rect 133150 675350 133570 675590
rect 133810 675350 133920 675590
rect 134160 675350 134250 675590
rect 134490 675350 134580 675590
rect 134820 675350 134910 675590
rect 135150 675350 135260 675590
rect 135500 675350 135590 675590
rect 135830 675350 135920 675590
rect 136160 675350 136250 675590
rect 136490 675350 136600 675590
rect 136840 675350 136930 675590
rect 137170 675350 137260 675590
rect 137500 675350 137590 675590
rect 137830 675350 137940 675590
rect 138180 675350 138270 675590
rect 138510 675350 138600 675590
rect 138840 675350 138930 675590
rect 139170 675350 139280 675590
rect 139520 675350 139610 675590
rect 139850 675350 139940 675590
rect 140180 675350 140270 675590
rect 140510 675350 140620 675590
rect 140860 675350 140950 675590
rect 141190 675350 141280 675590
rect 141520 675350 141610 675590
rect 141850 675350 141960 675590
rect 142200 675350 142290 675590
rect 142530 675350 142620 675590
rect 142860 675350 142950 675590
rect 143190 675350 143300 675590
rect 143540 675350 143630 675590
rect 143870 675350 143960 675590
rect 144200 675350 144290 675590
rect 144530 675350 144950 675590
rect 145190 675350 145300 675590
rect 145540 675350 145630 675590
rect 145870 675350 145960 675590
rect 146200 675350 146290 675590
rect 146530 675350 146640 675590
rect 146880 675350 146970 675590
rect 147210 675350 147300 675590
rect 147540 675350 147630 675590
rect 147870 675350 147980 675590
rect 148220 675350 148310 675590
rect 148550 675350 148640 675590
rect 148880 675350 148970 675590
rect 149210 675350 149320 675590
rect 149560 675350 149650 675590
rect 149890 675350 149980 675590
rect 150220 675350 150310 675590
rect 150550 675350 150660 675590
rect 150900 675350 150990 675590
rect 151230 675350 151320 675590
rect 151560 675350 151650 675590
rect 151890 675350 152000 675590
rect 152240 675350 152330 675590
rect 152570 675350 152660 675590
rect 152900 675350 152990 675590
rect 153230 675350 153340 675590
rect 153580 675350 153670 675590
rect 153910 675350 154000 675590
rect 154240 675350 154330 675590
rect 154570 675350 154680 675590
rect 154920 675350 155010 675590
rect 155250 675350 155340 675590
rect 155580 675350 155670 675590
rect 155910 675579 162436 675590
rect 155910 675350 157520 675579
rect 108560 675340 157520 675350
rect 103643 675339 157520 675340
rect 157780 675339 157880 675579
rect 158140 675339 158240 675579
rect 158500 675339 158600 675579
rect 158860 675339 162436 675579
rect 103643 675240 162436 675339
rect 103643 675000 107220 675240
rect 107480 675000 107580 675240
rect 107840 675000 107940 675240
rect 108200 675000 108300 675240
rect 108560 675000 110810 675240
rect 111050 675000 111160 675240
rect 111400 675000 111490 675240
rect 111730 675000 111820 675240
rect 112060 675000 112150 675240
rect 112390 675000 112500 675240
rect 112740 675000 112830 675240
rect 113070 675000 113160 675240
rect 113400 675000 113490 675240
rect 113730 675000 113840 675240
rect 114080 675000 114170 675240
rect 114410 675000 114500 675240
rect 114740 675000 114830 675240
rect 115070 675000 115180 675240
rect 115420 675000 115510 675240
rect 115750 675000 115840 675240
rect 116080 675000 116170 675240
rect 116410 675000 116520 675240
rect 116760 675000 116850 675240
rect 117090 675000 117180 675240
rect 117420 675000 117510 675240
rect 117750 675000 117860 675240
rect 118100 675000 118190 675240
rect 118430 675000 118520 675240
rect 118760 675000 118850 675240
rect 119090 675000 119200 675240
rect 119440 675000 119530 675240
rect 119770 675000 119860 675240
rect 120100 675000 120190 675240
rect 120430 675000 120540 675240
rect 120780 675000 120870 675240
rect 121110 675000 121200 675240
rect 121440 675000 121530 675240
rect 121770 675000 122190 675240
rect 122430 675000 122540 675240
rect 122780 675000 122870 675240
rect 123110 675000 123200 675240
rect 123440 675000 123530 675240
rect 123770 675000 123880 675240
rect 124120 675000 124210 675240
rect 124450 675000 124540 675240
rect 124780 675000 124870 675240
rect 125110 675000 125220 675240
rect 125460 675000 125550 675240
rect 125790 675000 125880 675240
rect 126120 675000 126210 675240
rect 126450 675000 126560 675240
rect 126800 675000 126890 675240
rect 127130 675000 127220 675240
rect 127460 675000 127550 675240
rect 127790 675000 127900 675240
rect 128140 675000 128230 675240
rect 128470 675000 128560 675240
rect 128800 675000 128890 675240
rect 129130 675000 129240 675240
rect 129480 675000 129570 675240
rect 129810 675000 129900 675240
rect 130140 675000 130230 675240
rect 130470 675000 130580 675240
rect 130820 675000 130910 675240
rect 131150 675000 131240 675240
rect 131480 675000 131570 675240
rect 131810 675000 131920 675240
rect 132160 675000 132250 675240
rect 132490 675000 132580 675240
rect 132820 675000 132910 675240
rect 133150 675000 133570 675240
rect 133810 675000 133920 675240
rect 134160 675000 134250 675240
rect 134490 675000 134580 675240
rect 134820 675000 134910 675240
rect 135150 675000 135260 675240
rect 135500 675000 135590 675240
rect 135830 675000 135920 675240
rect 136160 675000 136250 675240
rect 136490 675000 136600 675240
rect 136840 675000 136930 675240
rect 137170 675000 137260 675240
rect 137500 675000 137590 675240
rect 137830 675000 137940 675240
rect 138180 675000 138270 675240
rect 138510 675000 138600 675240
rect 138840 675000 138930 675240
rect 139170 675000 139280 675240
rect 139520 675000 139610 675240
rect 139850 675000 139940 675240
rect 140180 675000 140270 675240
rect 140510 675000 140620 675240
rect 140860 675000 140950 675240
rect 141190 675000 141280 675240
rect 141520 675000 141610 675240
rect 141850 675000 141960 675240
rect 142200 675000 142290 675240
rect 142530 675000 142620 675240
rect 142860 675000 142950 675240
rect 143190 675000 143300 675240
rect 143540 675000 143630 675240
rect 143870 675000 143960 675240
rect 144200 675000 144290 675240
rect 144530 675000 144950 675240
rect 145190 675000 145300 675240
rect 145540 675000 145630 675240
rect 145870 675000 145960 675240
rect 146200 675000 146290 675240
rect 146530 675000 146640 675240
rect 146880 675000 146970 675240
rect 147210 675000 147300 675240
rect 147540 675000 147630 675240
rect 147870 675000 147980 675240
rect 148220 675000 148310 675240
rect 148550 675000 148640 675240
rect 148880 675000 148970 675240
rect 149210 675000 149320 675240
rect 149560 675000 149650 675240
rect 149890 675000 149980 675240
rect 150220 675000 150310 675240
rect 150550 675000 150660 675240
rect 150900 675000 150990 675240
rect 151230 675000 151320 675240
rect 151560 675000 151650 675240
rect 151890 675000 152000 675240
rect 152240 675000 152330 675240
rect 152570 675000 152660 675240
rect 152900 675000 152990 675240
rect 153230 675000 153340 675240
rect 153580 675000 153670 675240
rect 153910 675000 154000 675240
rect 154240 675000 154330 675240
rect 154570 675000 154680 675240
rect 154920 675000 155010 675240
rect 155250 675000 155340 675240
rect 155580 675000 155670 675240
rect 155910 675239 162436 675240
rect 155910 675000 157520 675239
rect 103643 674999 157520 675000
rect 157780 674999 157880 675239
rect 158140 674999 158240 675239
rect 158500 674999 158600 675239
rect 158860 674999 162436 675239
rect 103643 674910 162436 674999
rect 103643 674900 110810 674910
rect 103643 674660 107220 674900
rect 107480 674660 107580 674900
rect 107840 674660 107940 674900
rect 108200 674660 108300 674900
rect 108560 674670 110810 674900
rect 111050 674670 111160 674910
rect 111400 674670 111490 674910
rect 111730 674670 111820 674910
rect 112060 674670 112150 674910
rect 112390 674670 112500 674910
rect 112740 674670 112830 674910
rect 113070 674670 113160 674910
rect 113400 674670 113490 674910
rect 113730 674670 113840 674910
rect 114080 674670 114170 674910
rect 114410 674670 114500 674910
rect 114740 674670 114830 674910
rect 115070 674670 115180 674910
rect 115420 674670 115510 674910
rect 115750 674670 115840 674910
rect 116080 674670 116170 674910
rect 116410 674670 116520 674910
rect 116760 674670 116850 674910
rect 117090 674670 117180 674910
rect 117420 674670 117510 674910
rect 117750 674670 117860 674910
rect 118100 674670 118190 674910
rect 118430 674670 118520 674910
rect 118760 674670 118850 674910
rect 119090 674670 119200 674910
rect 119440 674670 119530 674910
rect 119770 674670 119860 674910
rect 120100 674670 120190 674910
rect 120430 674670 120540 674910
rect 120780 674670 120870 674910
rect 121110 674670 121200 674910
rect 121440 674670 121530 674910
rect 121770 674670 122190 674910
rect 122430 674670 122540 674910
rect 122780 674670 122870 674910
rect 123110 674670 123200 674910
rect 123440 674670 123530 674910
rect 123770 674670 123880 674910
rect 124120 674670 124210 674910
rect 124450 674670 124540 674910
rect 124780 674670 124870 674910
rect 125110 674670 125220 674910
rect 125460 674670 125550 674910
rect 125790 674670 125880 674910
rect 126120 674670 126210 674910
rect 126450 674670 126560 674910
rect 126800 674670 126890 674910
rect 127130 674670 127220 674910
rect 127460 674670 127550 674910
rect 127790 674670 127900 674910
rect 128140 674670 128230 674910
rect 128470 674670 128560 674910
rect 128800 674670 128890 674910
rect 129130 674670 129240 674910
rect 129480 674670 129570 674910
rect 129810 674670 129900 674910
rect 130140 674670 130230 674910
rect 130470 674670 130580 674910
rect 130820 674670 130910 674910
rect 131150 674670 131240 674910
rect 131480 674670 131570 674910
rect 131810 674670 131920 674910
rect 132160 674670 132250 674910
rect 132490 674670 132580 674910
rect 132820 674670 132910 674910
rect 133150 674670 133570 674910
rect 133810 674670 133920 674910
rect 134160 674670 134250 674910
rect 134490 674670 134580 674910
rect 134820 674670 134910 674910
rect 135150 674670 135260 674910
rect 135500 674670 135590 674910
rect 135830 674670 135920 674910
rect 136160 674670 136250 674910
rect 136490 674670 136600 674910
rect 136840 674670 136930 674910
rect 137170 674670 137260 674910
rect 137500 674670 137590 674910
rect 137830 674670 137940 674910
rect 138180 674670 138270 674910
rect 138510 674670 138600 674910
rect 138840 674670 138930 674910
rect 139170 674670 139280 674910
rect 139520 674670 139610 674910
rect 139850 674670 139940 674910
rect 140180 674670 140270 674910
rect 140510 674670 140620 674910
rect 140860 674670 140950 674910
rect 141190 674670 141280 674910
rect 141520 674670 141610 674910
rect 141850 674670 141960 674910
rect 142200 674670 142290 674910
rect 142530 674670 142620 674910
rect 142860 674670 142950 674910
rect 143190 674670 143300 674910
rect 143540 674670 143630 674910
rect 143870 674670 143960 674910
rect 144200 674670 144290 674910
rect 144530 674670 144950 674910
rect 145190 674670 145300 674910
rect 145540 674670 145630 674910
rect 145870 674670 145960 674910
rect 146200 674670 146290 674910
rect 146530 674670 146640 674910
rect 146880 674670 146970 674910
rect 147210 674670 147300 674910
rect 147540 674670 147630 674910
rect 147870 674670 147980 674910
rect 148220 674670 148310 674910
rect 148550 674670 148640 674910
rect 148880 674670 148970 674910
rect 149210 674670 149320 674910
rect 149560 674670 149650 674910
rect 149890 674670 149980 674910
rect 150220 674670 150310 674910
rect 150550 674670 150660 674910
rect 150900 674670 150990 674910
rect 151230 674670 151320 674910
rect 151560 674670 151650 674910
rect 151890 674670 152000 674910
rect 152240 674670 152330 674910
rect 152570 674670 152660 674910
rect 152900 674670 152990 674910
rect 153230 674670 153340 674910
rect 153580 674670 153670 674910
rect 153910 674670 154000 674910
rect 154240 674670 154330 674910
rect 154570 674670 154680 674910
rect 154920 674670 155010 674910
rect 155250 674670 155340 674910
rect 155580 674670 155670 674910
rect 155910 674899 162436 674910
rect 155910 674670 157520 674899
rect 108560 674660 157520 674670
rect 103643 674659 157520 674660
rect 157780 674659 157880 674899
rect 158140 674659 158240 674899
rect 158500 674659 158600 674899
rect 158860 674659 162436 674899
rect 103643 674580 162436 674659
rect 103643 674560 110810 674580
rect 103643 674320 107220 674560
rect 107480 674320 107580 674560
rect 107840 674320 107940 674560
rect 108200 674320 108300 674560
rect 108560 674340 110810 674560
rect 111050 674340 111160 674580
rect 111400 674340 111490 674580
rect 111730 674340 111820 674580
rect 112060 674340 112150 674580
rect 112390 674340 112500 674580
rect 112740 674340 112830 674580
rect 113070 674340 113160 674580
rect 113400 674340 113490 674580
rect 113730 674340 113840 674580
rect 114080 674340 114170 674580
rect 114410 674340 114500 674580
rect 114740 674340 114830 674580
rect 115070 674340 115180 674580
rect 115420 674340 115510 674580
rect 115750 674340 115840 674580
rect 116080 674340 116170 674580
rect 116410 674340 116520 674580
rect 116760 674340 116850 674580
rect 117090 674340 117180 674580
rect 117420 674340 117510 674580
rect 117750 674340 117860 674580
rect 118100 674340 118190 674580
rect 118430 674340 118520 674580
rect 118760 674340 118850 674580
rect 119090 674340 119200 674580
rect 119440 674340 119530 674580
rect 119770 674340 119860 674580
rect 120100 674340 120190 674580
rect 120430 674340 120540 674580
rect 120780 674340 120870 674580
rect 121110 674340 121200 674580
rect 121440 674340 121530 674580
rect 121770 674340 122190 674580
rect 122430 674340 122540 674580
rect 122780 674340 122870 674580
rect 123110 674340 123200 674580
rect 123440 674340 123530 674580
rect 123770 674340 123880 674580
rect 124120 674340 124210 674580
rect 124450 674340 124540 674580
rect 124780 674340 124870 674580
rect 125110 674340 125220 674580
rect 125460 674340 125550 674580
rect 125790 674340 125880 674580
rect 126120 674340 126210 674580
rect 126450 674340 126560 674580
rect 126800 674340 126890 674580
rect 127130 674340 127220 674580
rect 127460 674340 127550 674580
rect 127790 674340 127900 674580
rect 128140 674340 128230 674580
rect 128470 674340 128560 674580
rect 128800 674340 128890 674580
rect 129130 674340 129240 674580
rect 129480 674340 129570 674580
rect 129810 674340 129900 674580
rect 130140 674340 130230 674580
rect 130470 674340 130580 674580
rect 130820 674340 130910 674580
rect 131150 674340 131240 674580
rect 131480 674340 131570 674580
rect 131810 674340 131920 674580
rect 132160 674340 132250 674580
rect 132490 674340 132580 674580
rect 132820 674340 132910 674580
rect 133150 674340 133570 674580
rect 133810 674340 133920 674580
rect 134160 674340 134250 674580
rect 134490 674340 134580 674580
rect 134820 674340 134910 674580
rect 135150 674340 135260 674580
rect 135500 674340 135590 674580
rect 135830 674340 135920 674580
rect 136160 674340 136250 674580
rect 136490 674340 136600 674580
rect 136840 674340 136930 674580
rect 137170 674340 137260 674580
rect 137500 674340 137590 674580
rect 137830 674340 137940 674580
rect 138180 674340 138270 674580
rect 138510 674340 138600 674580
rect 138840 674340 138930 674580
rect 139170 674340 139280 674580
rect 139520 674340 139610 674580
rect 139850 674340 139940 674580
rect 140180 674340 140270 674580
rect 140510 674340 140620 674580
rect 140860 674340 140950 674580
rect 141190 674340 141280 674580
rect 141520 674340 141610 674580
rect 141850 674340 141960 674580
rect 142200 674340 142290 674580
rect 142530 674340 142620 674580
rect 142860 674340 142950 674580
rect 143190 674340 143300 674580
rect 143540 674340 143630 674580
rect 143870 674340 143960 674580
rect 144200 674340 144290 674580
rect 144530 674340 144950 674580
rect 145190 674340 145300 674580
rect 145540 674340 145630 674580
rect 145870 674340 145960 674580
rect 146200 674340 146290 674580
rect 146530 674340 146640 674580
rect 146880 674340 146970 674580
rect 147210 674340 147300 674580
rect 147540 674340 147630 674580
rect 147870 674340 147980 674580
rect 148220 674340 148310 674580
rect 148550 674340 148640 674580
rect 148880 674340 148970 674580
rect 149210 674340 149320 674580
rect 149560 674340 149650 674580
rect 149890 674340 149980 674580
rect 150220 674340 150310 674580
rect 150550 674340 150660 674580
rect 150900 674340 150990 674580
rect 151230 674340 151320 674580
rect 151560 674340 151650 674580
rect 151890 674340 152000 674580
rect 152240 674340 152330 674580
rect 152570 674340 152660 674580
rect 152900 674340 152990 674580
rect 153230 674340 153340 674580
rect 153580 674340 153670 674580
rect 153910 674340 154000 674580
rect 154240 674340 154330 674580
rect 154570 674340 154680 674580
rect 154920 674340 155010 674580
rect 155250 674340 155340 674580
rect 155580 674340 155670 674580
rect 155910 674559 162436 674580
rect 155910 674340 157520 674559
rect 108560 674320 157520 674340
rect 103643 674319 157520 674320
rect 157780 674319 157880 674559
rect 158140 674319 158240 674559
rect 158500 674319 158600 674559
rect 158860 674319 162436 674559
rect 103643 674250 162436 674319
rect 103643 674152 110810 674250
rect 103643 657627 108640 674152
rect 110760 674010 110810 674152
rect 111050 674010 111160 674250
rect 111400 674010 111490 674250
rect 111730 674010 111820 674250
rect 112060 674010 112150 674250
rect 112390 674010 112500 674250
rect 112740 674010 112830 674250
rect 113070 674010 113160 674250
rect 113400 674010 113490 674250
rect 113730 674010 113840 674250
rect 114080 674010 114170 674250
rect 114410 674010 114500 674250
rect 114740 674010 114830 674250
rect 115070 674010 115180 674250
rect 115420 674010 115510 674250
rect 115750 674010 115840 674250
rect 116080 674010 116170 674250
rect 116410 674010 116520 674250
rect 116760 674010 116850 674250
rect 117090 674010 117180 674250
rect 117420 674010 117510 674250
rect 117750 674010 117860 674250
rect 118100 674010 118190 674250
rect 118430 674010 118520 674250
rect 118760 674010 118850 674250
rect 119090 674010 119200 674250
rect 119440 674010 119530 674250
rect 119770 674010 119860 674250
rect 120100 674010 120190 674250
rect 120430 674010 120540 674250
rect 120780 674010 120870 674250
rect 121110 674010 121200 674250
rect 121440 674010 121530 674250
rect 121770 674010 122190 674250
rect 122430 674010 122540 674250
rect 122780 674010 122870 674250
rect 123110 674010 123200 674250
rect 123440 674010 123530 674250
rect 123770 674010 123880 674250
rect 124120 674010 124210 674250
rect 124450 674010 124540 674250
rect 124780 674010 124870 674250
rect 125110 674010 125220 674250
rect 125460 674010 125550 674250
rect 125790 674010 125880 674250
rect 126120 674010 126210 674250
rect 126450 674010 126560 674250
rect 126800 674010 126890 674250
rect 127130 674010 127220 674250
rect 127460 674010 127550 674250
rect 127790 674010 127900 674250
rect 128140 674010 128230 674250
rect 128470 674010 128560 674250
rect 128800 674010 128890 674250
rect 129130 674010 129240 674250
rect 129480 674010 129570 674250
rect 129810 674010 129900 674250
rect 130140 674010 130230 674250
rect 130470 674010 130580 674250
rect 130820 674010 130910 674250
rect 131150 674010 131240 674250
rect 131480 674010 131570 674250
rect 131810 674010 131920 674250
rect 132160 674010 132250 674250
rect 132490 674010 132580 674250
rect 132820 674010 132910 674250
rect 133150 674010 133570 674250
rect 133810 674010 133920 674250
rect 134160 674010 134250 674250
rect 134490 674010 134580 674250
rect 134820 674010 134910 674250
rect 135150 674010 135260 674250
rect 135500 674010 135590 674250
rect 135830 674010 135920 674250
rect 136160 674010 136250 674250
rect 136490 674010 136600 674250
rect 136840 674010 136930 674250
rect 137170 674010 137260 674250
rect 137500 674010 137590 674250
rect 137830 674010 137940 674250
rect 138180 674010 138270 674250
rect 138510 674010 138600 674250
rect 138840 674010 138930 674250
rect 139170 674010 139280 674250
rect 139520 674010 139610 674250
rect 139850 674010 139940 674250
rect 140180 674010 140270 674250
rect 140510 674010 140620 674250
rect 140860 674010 140950 674250
rect 141190 674010 141280 674250
rect 141520 674010 141610 674250
rect 141850 674010 141960 674250
rect 142200 674010 142290 674250
rect 142530 674010 142620 674250
rect 142860 674010 142950 674250
rect 143190 674010 143300 674250
rect 143540 674010 143630 674250
rect 143870 674010 143960 674250
rect 144200 674010 144290 674250
rect 144530 674010 144950 674250
rect 145190 674010 145300 674250
rect 145540 674010 145630 674250
rect 145870 674010 145960 674250
rect 146200 674010 146290 674250
rect 146530 674010 146640 674250
rect 146880 674010 146970 674250
rect 147210 674010 147300 674250
rect 147540 674010 147630 674250
rect 147870 674010 147980 674250
rect 148220 674010 148310 674250
rect 148550 674010 148640 674250
rect 148880 674010 148970 674250
rect 149210 674010 149320 674250
rect 149560 674010 149650 674250
rect 149890 674010 149980 674250
rect 150220 674010 150310 674250
rect 150550 674010 150660 674250
rect 150900 674010 150990 674250
rect 151230 674010 151320 674250
rect 151560 674010 151650 674250
rect 151890 674010 152000 674250
rect 152240 674010 152330 674250
rect 152570 674010 152660 674250
rect 152900 674010 152990 674250
rect 153230 674010 153340 674250
rect 153580 674010 153670 674250
rect 153910 674010 154000 674250
rect 154240 674010 154330 674250
rect 154570 674010 154680 674250
rect 154920 674010 155010 674250
rect 155250 674010 155340 674250
rect 155580 674010 155670 674250
rect 155910 674152 162436 674250
rect 155910 674010 155960 674152
rect 110760 673900 155960 674010
rect 110760 673660 110810 673900
rect 111050 673660 111160 673900
rect 111400 673660 111490 673900
rect 111730 673660 111820 673900
rect 112060 673660 112150 673900
rect 112390 673660 112500 673900
rect 112740 673660 112830 673900
rect 113070 673660 113160 673900
rect 113400 673660 113490 673900
rect 113730 673660 113840 673900
rect 114080 673660 114170 673900
rect 114410 673660 114500 673900
rect 114740 673660 114830 673900
rect 115070 673660 115180 673900
rect 115420 673660 115510 673900
rect 115750 673660 115840 673900
rect 116080 673660 116170 673900
rect 116410 673660 116520 673900
rect 116760 673660 116850 673900
rect 117090 673660 117180 673900
rect 117420 673660 117510 673900
rect 117750 673660 117860 673900
rect 118100 673660 118190 673900
rect 118430 673660 118520 673900
rect 118760 673660 118850 673900
rect 119090 673660 119200 673900
rect 119440 673660 119530 673900
rect 119770 673660 119860 673900
rect 120100 673660 120190 673900
rect 120430 673660 120540 673900
rect 120780 673660 120870 673900
rect 121110 673660 121200 673900
rect 121440 673660 121530 673900
rect 121770 673660 122190 673900
rect 122430 673660 122540 673900
rect 122780 673660 122870 673900
rect 123110 673660 123200 673900
rect 123440 673660 123530 673900
rect 123770 673660 123880 673900
rect 124120 673660 124210 673900
rect 124450 673660 124540 673900
rect 124780 673660 124870 673900
rect 125110 673660 125220 673900
rect 125460 673660 125550 673900
rect 125790 673660 125880 673900
rect 126120 673660 126210 673900
rect 126450 673660 126560 673900
rect 126800 673660 126890 673900
rect 127130 673660 127220 673900
rect 127460 673660 127550 673900
rect 127790 673660 127900 673900
rect 128140 673660 128230 673900
rect 128470 673660 128560 673900
rect 128800 673660 128890 673900
rect 129130 673660 129240 673900
rect 129480 673660 129570 673900
rect 129810 673660 129900 673900
rect 130140 673660 130230 673900
rect 130470 673660 130580 673900
rect 130820 673660 130910 673900
rect 131150 673660 131240 673900
rect 131480 673660 131570 673900
rect 131810 673660 131920 673900
rect 132160 673660 132250 673900
rect 132490 673660 132580 673900
rect 132820 673660 132910 673900
rect 133150 673660 133570 673900
rect 133810 673660 133920 673900
rect 134160 673660 134250 673900
rect 134490 673660 134580 673900
rect 134820 673660 134910 673900
rect 135150 673660 135260 673900
rect 135500 673660 135590 673900
rect 135830 673660 135920 673900
rect 136160 673660 136250 673900
rect 136490 673660 136600 673900
rect 136840 673660 136930 673900
rect 137170 673660 137260 673900
rect 137500 673660 137590 673900
rect 137830 673660 137940 673900
rect 138180 673660 138270 673900
rect 138510 673660 138600 673900
rect 138840 673660 138930 673900
rect 139170 673660 139280 673900
rect 139520 673660 139610 673900
rect 139850 673660 139940 673900
rect 140180 673660 140270 673900
rect 140510 673660 140620 673900
rect 140860 673660 140950 673900
rect 141190 673660 141280 673900
rect 141520 673660 141610 673900
rect 141850 673660 141960 673900
rect 142200 673660 142290 673900
rect 142530 673660 142620 673900
rect 142860 673660 142950 673900
rect 143190 673660 143300 673900
rect 143540 673660 143630 673900
rect 143870 673660 143960 673900
rect 144200 673660 144290 673900
rect 144530 673660 144950 673900
rect 145190 673660 145300 673900
rect 145540 673660 145630 673900
rect 145870 673660 145960 673900
rect 146200 673660 146290 673900
rect 146530 673660 146640 673900
rect 146880 673660 146970 673900
rect 147210 673660 147300 673900
rect 147540 673660 147630 673900
rect 147870 673660 147980 673900
rect 148220 673660 148310 673900
rect 148550 673660 148640 673900
rect 148880 673660 148970 673900
rect 149210 673660 149320 673900
rect 149560 673660 149650 673900
rect 149890 673660 149980 673900
rect 150220 673660 150310 673900
rect 150550 673660 150660 673900
rect 150900 673660 150990 673900
rect 151230 673660 151320 673900
rect 151560 673660 151650 673900
rect 151890 673660 152000 673900
rect 152240 673660 152330 673900
rect 152570 673660 152660 673900
rect 152900 673660 152990 673900
rect 153230 673660 153340 673900
rect 153580 673660 153670 673900
rect 153910 673660 154000 673900
rect 154240 673660 154330 673900
rect 154570 673660 154680 673900
rect 154920 673660 155010 673900
rect 155250 673660 155340 673900
rect 155580 673660 155670 673900
rect 155910 673660 155960 673900
rect 110760 673570 155960 673660
rect 110760 673330 110810 673570
rect 111050 673330 111160 673570
rect 111400 673330 111490 673570
rect 111730 673330 111820 673570
rect 112060 673330 112150 673570
rect 112390 673330 112500 673570
rect 112740 673330 112830 673570
rect 113070 673330 113160 673570
rect 113400 673330 113490 673570
rect 113730 673330 113840 673570
rect 114080 673330 114170 673570
rect 114410 673330 114500 673570
rect 114740 673330 114830 673570
rect 115070 673330 115180 673570
rect 115420 673330 115510 673570
rect 115750 673330 115840 673570
rect 116080 673330 116170 673570
rect 116410 673330 116520 673570
rect 116760 673330 116850 673570
rect 117090 673330 117180 673570
rect 117420 673330 117510 673570
rect 117750 673330 117860 673570
rect 118100 673330 118190 673570
rect 118430 673330 118520 673570
rect 118760 673330 118850 673570
rect 119090 673330 119200 673570
rect 119440 673330 119530 673570
rect 119770 673330 119860 673570
rect 120100 673330 120190 673570
rect 120430 673330 120540 673570
rect 120780 673330 120870 673570
rect 121110 673330 121200 673570
rect 121440 673330 121530 673570
rect 121770 673330 122190 673570
rect 122430 673330 122540 673570
rect 122780 673330 122870 673570
rect 123110 673330 123200 673570
rect 123440 673330 123530 673570
rect 123770 673330 123880 673570
rect 124120 673330 124210 673570
rect 124450 673330 124540 673570
rect 124780 673330 124870 673570
rect 125110 673330 125220 673570
rect 125460 673330 125550 673570
rect 125790 673330 125880 673570
rect 126120 673330 126210 673570
rect 126450 673330 126560 673570
rect 126800 673330 126890 673570
rect 127130 673330 127220 673570
rect 127460 673330 127550 673570
rect 127790 673330 127900 673570
rect 128140 673330 128230 673570
rect 128470 673330 128560 673570
rect 128800 673330 128890 673570
rect 129130 673330 129240 673570
rect 129480 673330 129570 673570
rect 129810 673330 129900 673570
rect 130140 673330 130230 673570
rect 130470 673330 130580 673570
rect 130820 673330 130910 673570
rect 131150 673330 131240 673570
rect 131480 673330 131570 673570
rect 131810 673330 131920 673570
rect 132160 673330 132250 673570
rect 132490 673330 132580 673570
rect 132820 673330 132910 673570
rect 133150 673330 133570 673570
rect 133810 673330 133920 673570
rect 134160 673330 134250 673570
rect 134490 673330 134580 673570
rect 134820 673330 134910 673570
rect 135150 673330 135260 673570
rect 135500 673330 135590 673570
rect 135830 673330 135920 673570
rect 136160 673330 136250 673570
rect 136490 673330 136600 673570
rect 136840 673330 136930 673570
rect 137170 673330 137260 673570
rect 137500 673330 137590 673570
rect 137830 673330 137940 673570
rect 138180 673330 138270 673570
rect 138510 673330 138600 673570
rect 138840 673330 138930 673570
rect 139170 673330 139280 673570
rect 139520 673330 139610 673570
rect 139850 673330 139940 673570
rect 140180 673330 140270 673570
rect 140510 673330 140620 673570
rect 140860 673330 140950 673570
rect 141190 673330 141280 673570
rect 141520 673330 141610 673570
rect 141850 673330 141960 673570
rect 142200 673330 142290 673570
rect 142530 673330 142620 673570
rect 142860 673330 142950 673570
rect 143190 673330 143300 673570
rect 143540 673330 143630 673570
rect 143870 673330 143960 673570
rect 144200 673330 144290 673570
rect 144530 673330 144950 673570
rect 145190 673330 145300 673570
rect 145540 673330 145630 673570
rect 145870 673330 145960 673570
rect 146200 673330 146290 673570
rect 146530 673330 146640 673570
rect 146880 673330 146970 673570
rect 147210 673330 147300 673570
rect 147540 673330 147630 673570
rect 147870 673330 147980 673570
rect 148220 673330 148310 673570
rect 148550 673330 148640 673570
rect 148880 673330 148970 673570
rect 149210 673330 149320 673570
rect 149560 673330 149650 673570
rect 149890 673330 149980 673570
rect 150220 673330 150310 673570
rect 150550 673330 150660 673570
rect 150900 673330 150990 673570
rect 151230 673330 151320 673570
rect 151560 673330 151650 673570
rect 151890 673330 152000 673570
rect 152240 673330 152330 673570
rect 152570 673330 152660 673570
rect 152900 673330 152990 673570
rect 153230 673330 153340 673570
rect 153580 673330 153670 673570
rect 153910 673330 154000 673570
rect 154240 673330 154330 673570
rect 154570 673330 154680 673570
rect 154920 673330 155010 673570
rect 155250 673330 155340 673570
rect 155580 673330 155670 673570
rect 155910 673330 155960 673570
rect 110760 673240 155960 673330
rect 110760 673000 110810 673240
rect 111050 673000 111160 673240
rect 111400 673000 111490 673240
rect 111730 673000 111820 673240
rect 112060 673000 112150 673240
rect 112390 673000 112500 673240
rect 112740 673000 112830 673240
rect 113070 673000 113160 673240
rect 113400 673000 113490 673240
rect 113730 673000 113840 673240
rect 114080 673000 114170 673240
rect 114410 673000 114500 673240
rect 114740 673000 114830 673240
rect 115070 673000 115180 673240
rect 115420 673000 115510 673240
rect 115750 673000 115840 673240
rect 116080 673000 116170 673240
rect 116410 673000 116520 673240
rect 116760 673000 116850 673240
rect 117090 673000 117180 673240
rect 117420 673000 117510 673240
rect 117750 673000 117860 673240
rect 118100 673000 118190 673240
rect 118430 673000 118520 673240
rect 118760 673000 118850 673240
rect 119090 673000 119200 673240
rect 119440 673000 119530 673240
rect 119770 673000 119860 673240
rect 120100 673000 120190 673240
rect 120430 673000 120540 673240
rect 120780 673000 120870 673240
rect 121110 673000 121200 673240
rect 121440 673000 121530 673240
rect 121770 673000 122190 673240
rect 122430 673000 122540 673240
rect 122780 673000 122870 673240
rect 123110 673000 123200 673240
rect 123440 673000 123530 673240
rect 123770 673000 123880 673240
rect 124120 673000 124210 673240
rect 124450 673000 124540 673240
rect 124780 673000 124870 673240
rect 125110 673000 125220 673240
rect 125460 673000 125550 673240
rect 125790 673000 125880 673240
rect 126120 673000 126210 673240
rect 126450 673000 126560 673240
rect 126800 673000 126890 673240
rect 127130 673000 127220 673240
rect 127460 673000 127550 673240
rect 127790 673000 127900 673240
rect 128140 673000 128230 673240
rect 128470 673000 128560 673240
rect 128800 673000 128890 673240
rect 129130 673000 129240 673240
rect 129480 673000 129570 673240
rect 129810 673000 129900 673240
rect 130140 673000 130230 673240
rect 130470 673000 130580 673240
rect 130820 673000 130910 673240
rect 131150 673000 131240 673240
rect 131480 673000 131570 673240
rect 131810 673000 131920 673240
rect 132160 673000 132250 673240
rect 132490 673000 132580 673240
rect 132820 673000 132910 673240
rect 133150 673000 133570 673240
rect 133810 673000 133920 673240
rect 134160 673000 134250 673240
rect 134490 673000 134580 673240
rect 134820 673000 134910 673240
rect 135150 673000 135260 673240
rect 135500 673000 135590 673240
rect 135830 673000 135920 673240
rect 136160 673000 136250 673240
rect 136490 673000 136600 673240
rect 136840 673000 136930 673240
rect 137170 673000 137260 673240
rect 137500 673000 137590 673240
rect 137830 673000 137940 673240
rect 138180 673000 138270 673240
rect 138510 673000 138600 673240
rect 138840 673000 138930 673240
rect 139170 673000 139280 673240
rect 139520 673000 139610 673240
rect 139850 673000 139940 673240
rect 140180 673000 140270 673240
rect 140510 673000 140620 673240
rect 140860 673000 140950 673240
rect 141190 673000 141280 673240
rect 141520 673000 141610 673240
rect 141850 673000 141960 673240
rect 142200 673000 142290 673240
rect 142530 673000 142620 673240
rect 142860 673000 142950 673240
rect 143190 673000 143300 673240
rect 143540 673000 143630 673240
rect 143870 673000 143960 673240
rect 144200 673000 144290 673240
rect 144530 673000 144950 673240
rect 145190 673000 145300 673240
rect 145540 673000 145630 673240
rect 145870 673000 145960 673240
rect 146200 673000 146290 673240
rect 146530 673000 146640 673240
rect 146880 673000 146970 673240
rect 147210 673000 147300 673240
rect 147540 673000 147630 673240
rect 147870 673000 147980 673240
rect 148220 673000 148310 673240
rect 148550 673000 148640 673240
rect 148880 673000 148970 673240
rect 149210 673000 149320 673240
rect 149560 673000 149650 673240
rect 149890 673000 149980 673240
rect 150220 673000 150310 673240
rect 150550 673000 150660 673240
rect 150900 673000 150990 673240
rect 151230 673000 151320 673240
rect 151560 673000 151650 673240
rect 151890 673000 152000 673240
rect 152240 673000 152330 673240
rect 152570 673000 152660 673240
rect 152900 673000 152990 673240
rect 153230 673000 153340 673240
rect 153580 673000 153670 673240
rect 153910 673000 154000 673240
rect 154240 673000 154330 673240
rect 154570 673000 154680 673240
rect 154920 673000 155010 673240
rect 155250 673000 155340 673240
rect 155580 673000 155670 673240
rect 155910 673000 155960 673240
rect 110760 672910 155960 673000
rect 110760 672670 110810 672910
rect 111050 672670 111160 672910
rect 111400 672670 111490 672910
rect 111730 672670 111820 672910
rect 112060 672670 112150 672910
rect 112390 672670 112500 672910
rect 112740 672670 112830 672910
rect 113070 672670 113160 672910
rect 113400 672670 113490 672910
rect 113730 672670 113840 672910
rect 114080 672670 114170 672910
rect 114410 672670 114500 672910
rect 114740 672670 114830 672910
rect 115070 672670 115180 672910
rect 115420 672670 115510 672910
rect 115750 672670 115840 672910
rect 116080 672670 116170 672910
rect 116410 672670 116520 672910
rect 116760 672670 116850 672910
rect 117090 672670 117180 672910
rect 117420 672670 117510 672910
rect 117750 672670 117860 672910
rect 118100 672670 118190 672910
rect 118430 672670 118520 672910
rect 118760 672670 118850 672910
rect 119090 672670 119200 672910
rect 119440 672670 119530 672910
rect 119770 672670 119860 672910
rect 120100 672670 120190 672910
rect 120430 672670 120540 672910
rect 120780 672670 120870 672910
rect 121110 672670 121200 672910
rect 121440 672670 121530 672910
rect 121770 672670 122190 672910
rect 122430 672670 122540 672910
rect 122780 672670 122870 672910
rect 123110 672670 123200 672910
rect 123440 672670 123530 672910
rect 123770 672670 123880 672910
rect 124120 672670 124210 672910
rect 124450 672670 124540 672910
rect 124780 672670 124870 672910
rect 125110 672670 125220 672910
rect 125460 672670 125550 672910
rect 125790 672670 125880 672910
rect 126120 672670 126210 672910
rect 126450 672670 126560 672910
rect 126800 672670 126890 672910
rect 127130 672670 127220 672910
rect 127460 672670 127550 672910
rect 127790 672670 127900 672910
rect 128140 672670 128230 672910
rect 128470 672670 128560 672910
rect 128800 672670 128890 672910
rect 129130 672670 129240 672910
rect 129480 672670 129570 672910
rect 129810 672670 129900 672910
rect 130140 672670 130230 672910
rect 130470 672670 130580 672910
rect 130820 672670 130910 672910
rect 131150 672670 131240 672910
rect 131480 672670 131570 672910
rect 131810 672670 131920 672910
rect 132160 672670 132250 672910
rect 132490 672670 132580 672910
rect 132820 672670 132910 672910
rect 133150 672670 133570 672910
rect 133810 672670 133920 672910
rect 134160 672670 134250 672910
rect 134490 672670 134580 672910
rect 134820 672670 134910 672910
rect 135150 672670 135260 672910
rect 135500 672670 135590 672910
rect 135830 672670 135920 672910
rect 136160 672670 136250 672910
rect 136490 672670 136600 672910
rect 136840 672670 136930 672910
rect 137170 672670 137260 672910
rect 137500 672670 137590 672910
rect 137830 672670 137940 672910
rect 138180 672670 138270 672910
rect 138510 672670 138600 672910
rect 138840 672670 138930 672910
rect 139170 672670 139280 672910
rect 139520 672670 139610 672910
rect 139850 672670 139940 672910
rect 140180 672670 140270 672910
rect 140510 672670 140620 672910
rect 140860 672670 140950 672910
rect 141190 672670 141280 672910
rect 141520 672670 141610 672910
rect 141850 672670 141960 672910
rect 142200 672670 142290 672910
rect 142530 672670 142620 672910
rect 142860 672670 142950 672910
rect 143190 672670 143300 672910
rect 143540 672670 143630 672910
rect 143870 672670 143960 672910
rect 144200 672670 144290 672910
rect 144530 672670 144950 672910
rect 145190 672670 145300 672910
rect 145540 672670 145630 672910
rect 145870 672670 145960 672910
rect 146200 672670 146290 672910
rect 146530 672670 146640 672910
rect 146880 672670 146970 672910
rect 147210 672670 147300 672910
rect 147540 672670 147630 672910
rect 147870 672670 147980 672910
rect 148220 672670 148310 672910
rect 148550 672670 148640 672910
rect 148880 672670 148970 672910
rect 149210 672670 149320 672910
rect 149560 672670 149650 672910
rect 149890 672670 149980 672910
rect 150220 672670 150310 672910
rect 150550 672670 150660 672910
rect 150900 672670 150990 672910
rect 151230 672670 151320 672910
rect 151560 672670 151650 672910
rect 151890 672670 152000 672910
rect 152240 672670 152330 672910
rect 152570 672670 152660 672910
rect 152900 672670 152990 672910
rect 153230 672670 153340 672910
rect 153580 672670 153670 672910
rect 153910 672670 154000 672910
rect 154240 672670 154330 672910
rect 154570 672670 154680 672910
rect 154920 672670 155010 672910
rect 155250 672670 155340 672910
rect 155580 672670 155670 672910
rect 155910 672670 155960 672910
rect 110760 672560 155960 672670
rect 110760 672320 110810 672560
rect 111050 672320 111160 672560
rect 111400 672320 111490 672560
rect 111730 672320 111820 672560
rect 112060 672320 112150 672560
rect 112390 672320 112500 672560
rect 112740 672320 112830 672560
rect 113070 672320 113160 672560
rect 113400 672320 113490 672560
rect 113730 672320 113840 672560
rect 114080 672320 114170 672560
rect 114410 672320 114500 672560
rect 114740 672320 114830 672560
rect 115070 672320 115180 672560
rect 115420 672320 115510 672560
rect 115750 672320 115840 672560
rect 116080 672320 116170 672560
rect 116410 672320 116520 672560
rect 116760 672320 116850 672560
rect 117090 672320 117180 672560
rect 117420 672320 117510 672560
rect 117750 672320 117860 672560
rect 118100 672320 118190 672560
rect 118430 672320 118520 672560
rect 118760 672320 118850 672560
rect 119090 672320 119200 672560
rect 119440 672320 119530 672560
rect 119770 672320 119860 672560
rect 120100 672320 120190 672560
rect 120430 672320 120540 672560
rect 120780 672320 120870 672560
rect 121110 672320 121200 672560
rect 121440 672320 121530 672560
rect 121770 672320 122190 672560
rect 122430 672320 122540 672560
rect 122780 672320 122870 672560
rect 123110 672320 123200 672560
rect 123440 672320 123530 672560
rect 123770 672320 123880 672560
rect 124120 672320 124210 672560
rect 124450 672320 124540 672560
rect 124780 672320 124870 672560
rect 125110 672320 125220 672560
rect 125460 672320 125550 672560
rect 125790 672320 125880 672560
rect 126120 672320 126210 672560
rect 126450 672320 126560 672560
rect 126800 672320 126890 672560
rect 127130 672320 127220 672560
rect 127460 672320 127550 672560
rect 127790 672320 127900 672560
rect 128140 672320 128230 672560
rect 128470 672320 128560 672560
rect 128800 672320 128890 672560
rect 129130 672320 129240 672560
rect 129480 672320 129570 672560
rect 129810 672320 129900 672560
rect 130140 672320 130230 672560
rect 130470 672320 130580 672560
rect 130820 672320 130910 672560
rect 131150 672320 131240 672560
rect 131480 672320 131570 672560
rect 131810 672320 131920 672560
rect 132160 672320 132250 672560
rect 132490 672320 132580 672560
rect 132820 672320 132910 672560
rect 133150 672320 133570 672560
rect 133810 672320 133920 672560
rect 134160 672320 134250 672560
rect 134490 672320 134580 672560
rect 134820 672320 134910 672560
rect 135150 672320 135260 672560
rect 135500 672320 135590 672560
rect 135830 672320 135920 672560
rect 136160 672320 136250 672560
rect 136490 672320 136600 672560
rect 136840 672320 136930 672560
rect 137170 672320 137260 672560
rect 137500 672320 137590 672560
rect 137830 672320 137940 672560
rect 138180 672320 138270 672560
rect 138510 672320 138600 672560
rect 138840 672320 138930 672560
rect 139170 672320 139280 672560
rect 139520 672320 139610 672560
rect 139850 672320 139940 672560
rect 140180 672320 140270 672560
rect 140510 672320 140620 672560
rect 140860 672320 140950 672560
rect 141190 672320 141280 672560
rect 141520 672320 141610 672560
rect 141850 672320 141960 672560
rect 142200 672320 142290 672560
rect 142530 672320 142620 672560
rect 142860 672320 142950 672560
rect 143190 672320 143300 672560
rect 143540 672320 143630 672560
rect 143870 672320 143960 672560
rect 144200 672320 144290 672560
rect 144530 672320 144950 672560
rect 145190 672320 145300 672560
rect 145540 672320 145630 672560
rect 145870 672320 145960 672560
rect 146200 672320 146290 672560
rect 146530 672320 146640 672560
rect 146880 672320 146970 672560
rect 147210 672320 147300 672560
rect 147540 672320 147630 672560
rect 147870 672320 147980 672560
rect 148220 672320 148310 672560
rect 148550 672320 148640 672560
rect 148880 672320 148970 672560
rect 149210 672320 149320 672560
rect 149560 672320 149650 672560
rect 149890 672320 149980 672560
rect 150220 672320 150310 672560
rect 150550 672320 150660 672560
rect 150900 672320 150990 672560
rect 151230 672320 151320 672560
rect 151560 672320 151650 672560
rect 151890 672320 152000 672560
rect 152240 672320 152330 672560
rect 152570 672320 152660 672560
rect 152900 672320 152990 672560
rect 153230 672320 153340 672560
rect 153580 672320 153670 672560
rect 153910 672320 154000 672560
rect 154240 672320 154330 672560
rect 154570 672320 154680 672560
rect 154920 672320 155010 672560
rect 155250 672320 155340 672560
rect 155580 672320 155670 672560
rect 155910 672320 155960 672560
rect 110760 671900 155960 672320
rect 110760 671660 110810 671900
rect 111050 671660 111140 671900
rect 111380 671660 111470 671900
rect 111710 671660 111800 671900
rect 112040 671660 112150 671900
rect 112390 671660 112480 671900
rect 112720 671660 112810 671900
rect 113050 671660 113140 671900
rect 113380 671660 113490 671900
rect 113730 671660 113820 671900
rect 114060 671660 114150 671900
rect 114390 671660 114480 671900
rect 114720 671660 114830 671900
rect 115070 671660 115160 671900
rect 115400 671660 115490 671900
rect 115730 671660 115820 671900
rect 116060 671660 116170 671900
rect 116410 671660 116500 671900
rect 116740 671660 116830 671900
rect 117070 671660 117160 671900
rect 117400 671660 117510 671900
rect 117750 671660 117840 671900
rect 118080 671660 118170 671900
rect 118410 671660 118500 671900
rect 118740 671660 118850 671900
rect 119090 671660 119180 671900
rect 119420 671660 119510 671900
rect 119750 671660 119840 671900
rect 120080 671660 120190 671900
rect 120430 671660 120520 671900
rect 120760 671660 120850 671900
rect 121090 671660 121180 671900
rect 121420 671660 121530 671900
rect 121770 671660 122190 671900
rect 122430 671660 122520 671900
rect 122760 671660 122850 671900
rect 123090 671660 123180 671900
rect 123420 671660 123530 671900
rect 123770 671660 123860 671900
rect 124100 671660 124190 671900
rect 124430 671660 124520 671900
rect 124760 671660 124870 671900
rect 125110 671660 125200 671900
rect 125440 671660 125530 671900
rect 125770 671660 125860 671900
rect 126100 671660 126210 671900
rect 126450 671660 126540 671900
rect 126780 671660 126870 671900
rect 127110 671660 127200 671900
rect 127440 671660 127550 671900
rect 127790 671660 127880 671900
rect 128120 671660 128210 671900
rect 128450 671660 128540 671900
rect 128780 671660 128890 671900
rect 129130 671660 129220 671900
rect 129460 671660 129550 671900
rect 129790 671660 129880 671900
rect 130120 671660 130230 671900
rect 130470 671660 130560 671900
rect 130800 671660 130890 671900
rect 131130 671660 131220 671900
rect 131460 671660 131570 671900
rect 131810 671660 131900 671900
rect 132140 671660 132230 671900
rect 132470 671660 132560 671900
rect 132800 671660 132910 671900
rect 133150 671660 133570 671900
rect 133810 671660 133900 671900
rect 134140 671660 134230 671900
rect 134470 671660 134560 671900
rect 134800 671660 134910 671900
rect 135150 671660 135240 671900
rect 135480 671660 135570 671900
rect 135810 671660 135900 671900
rect 136140 671660 136250 671900
rect 136490 671660 136580 671900
rect 136820 671660 136910 671900
rect 137150 671660 137240 671900
rect 137480 671660 137590 671900
rect 137830 671660 137920 671900
rect 138160 671660 138250 671900
rect 138490 671660 138580 671900
rect 138820 671660 138930 671900
rect 139170 671660 139260 671900
rect 139500 671660 139590 671900
rect 139830 671660 139920 671900
rect 140160 671660 140270 671900
rect 140510 671660 140600 671900
rect 140840 671660 140930 671900
rect 141170 671660 141260 671900
rect 141500 671660 141610 671900
rect 141850 671660 141940 671900
rect 142180 671660 142270 671900
rect 142510 671660 142600 671900
rect 142840 671660 142950 671900
rect 143190 671660 143280 671900
rect 143520 671660 143610 671900
rect 143850 671660 143940 671900
rect 144180 671660 144290 671900
rect 144530 671660 144950 671900
rect 145190 671660 145280 671900
rect 145520 671660 145610 671900
rect 145850 671660 145940 671900
rect 146180 671660 146290 671900
rect 146530 671660 146620 671900
rect 146860 671660 146950 671900
rect 147190 671660 147280 671900
rect 147520 671660 147630 671900
rect 147870 671660 147960 671900
rect 148200 671660 148290 671900
rect 148530 671660 148620 671900
rect 148860 671660 148970 671900
rect 149210 671660 149300 671900
rect 149540 671660 149630 671900
rect 149870 671660 149960 671900
rect 150200 671660 150310 671900
rect 150550 671660 150640 671900
rect 150880 671660 150970 671900
rect 151210 671660 151300 671900
rect 151540 671660 151650 671900
rect 151890 671660 151980 671900
rect 152220 671660 152310 671900
rect 152550 671660 152640 671900
rect 152880 671660 152990 671900
rect 153230 671660 153320 671900
rect 153560 671660 153650 671900
rect 153890 671660 153980 671900
rect 154220 671660 154330 671900
rect 154570 671660 154660 671900
rect 154900 671660 154990 671900
rect 155230 671660 155320 671900
rect 155560 671660 155670 671900
rect 155910 671660 155960 671900
rect 110760 671550 155960 671660
rect 110760 671310 110810 671550
rect 111050 671310 111140 671550
rect 111380 671310 111470 671550
rect 111710 671310 111800 671550
rect 112040 671310 112150 671550
rect 112390 671310 112480 671550
rect 112720 671310 112810 671550
rect 113050 671310 113140 671550
rect 113380 671310 113490 671550
rect 113730 671310 113820 671550
rect 114060 671310 114150 671550
rect 114390 671310 114480 671550
rect 114720 671310 114830 671550
rect 115070 671310 115160 671550
rect 115400 671310 115490 671550
rect 115730 671310 115820 671550
rect 116060 671310 116170 671550
rect 116410 671310 116500 671550
rect 116740 671310 116830 671550
rect 117070 671310 117160 671550
rect 117400 671310 117510 671550
rect 117750 671310 117840 671550
rect 118080 671310 118170 671550
rect 118410 671310 118500 671550
rect 118740 671310 118850 671550
rect 119090 671310 119180 671550
rect 119420 671310 119510 671550
rect 119750 671310 119840 671550
rect 120080 671310 120190 671550
rect 120430 671310 120520 671550
rect 120760 671310 120850 671550
rect 121090 671310 121180 671550
rect 121420 671310 121530 671550
rect 121770 671310 122190 671550
rect 122430 671310 122520 671550
rect 122760 671310 122850 671550
rect 123090 671310 123180 671550
rect 123420 671310 123530 671550
rect 123770 671310 123860 671550
rect 124100 671310 124190 671550
rect 124430 671310 124520 671550
rect 124760 671310 124870 671550
rect 125110 671310 125200 671550
rect 125440 671310 125530 671550
rect 125770 671310 125860 671550
rect 126100 671310 126210 671550
rect 126450 671310 126540 671550
rect 126780 671310 126870 671550
rect 127110 671310 127200 671550
rect 127440 671310 127550 671550
rect 127790 671310 127880 671550
rect 128120 671310 128210 671550
rect 128450 671310 128540 671550
rect 128780 671310 128890 671550
rect 129130 671310 129220 671550
rect 129460 671310 129550 671550
rect 129790 671310 129880 671550
rect 130120 671310 130230 671550
rect 130470 671310 130560 671550
rect 130800 671310 130890 671550
rect 131130 671310 131220 671550
rect 131460 671310 131570 671550
rect 131810 671310 131900 671550
rect 132140 671310 132230 671550
rect 132470 671310 132560 671550
rect 132800 671310 132910 671550
rect 133150 671310 133570 671550
rect 133810 671310 133900 671550
rect 134140 671310 134230 671550
rect 134470 671310 134560 671550
rect 134800 671310 134910 671550
rect 135150 671310 135240 671550
rect 135480 671310 135570 671550
rect 135810 671310 135900 671550
rect 136140 671310 136250 671550
rect 136490 671310 136580 671550
rect 136820 671310 136910 671550
rect 137150 671310 137240 671550
rect 137480 671310 137590 671550
rect 137830 671310 137920 671550
rect 138160 671310 138250 671550
rect 138490 671310 138580 671550
rect 138820 671310 138930 671550
rect 139170 671310 139260 671550
rect 139500 671310 139590 671550
rect 139830 671310 139920 671550
rect 140160 671310 140270 671550
rect 140510 671310 140600 671550
rect 140840 671310 140930 671550
rect 141170 671310 141260 671550
rect 141500 671310 141610 671550
rect 141850 671310 141940 671550
rect 142180 671310 142270 671550
rect 142510 671310 142600 671550
rect 142840 671310 142950 671550
rect 143190 671310 143280 671550
rect 143520 671310 143610 671550
rect 143850 671310 143940 671550
rect 144180 671310 144290 671550
rect 144530 671310 144950 671550
rect 145190 671310 145280 671550
rect 145520 671310 145610 671550
rect 145850 671310 145940 671550
rect 146180 671310 146290 671550
rect 146530 671310 146620 671550
rect 146860 671310 146950 671550
rect 147190 671310 147280 671550
rect 147520 671310 147630 671550
rect 147870 671310 147960 671550
rect 148200 671310 148290 671550
rect 148530 671310 148620 671550
rect 148860 671310 148970 671550
rect 149210 671310 149300 671550
rect 149540 671310 149630 671550
rect 149870 671310 149960 671550
rect 150200 671310 150310 671550
rect 150550 671310 150640 671550
rect 150880 671310 150970 671550
rect 151210 671310 151300 671550
rect 151540 671310 151650 671550
rect 151890 671310 151980 671550
rect 152220 671310 152310 671550
rect 152550 671310 152640 671550
rect 152880 671310 152990 671550
rect 153230 671310 153320 671550
rect 153560 671310 153650 671550
rect 153890 671310 153980 671550
rect 154220 671310 154330 671550
rect 154570 671310 154660 671550
rect 154900 671310 154990 671550
rect 155230 671310 155320 671550
rect 155560 671310 155670 671550
rect 155910 671310 155960 671550
rect 110760 671220 155960 671310
rect 110760 670980 110810 671220
rect 111050 670980 111140 671220
rect 111380 670980 111470 671220
rect 111710 670980 111800 671220
rect 112040 670980 112150 671220
rect 112390 670980 112480 671220
rect 112720 670980 112810 671220
rect 113050 670980 113140 671220
rect 113380 670980 113490 671220
rect 113730 670980 113820 671220
rect 114060 670980 114150 671220
rect 114390 670980 114480 671220
rect 114720 670980 114830 671220
rect 115070 670980 115160 671220
rect 115400 670980 115490 671220
rect 115730 670980 115820 671220
rect 116060 670980 116170 671220
rect 116410 670980 116500 671220
rect 116740 670980 116830 671220
rect 117070 670980 117160 671220
rect 117400 670980 117510 671220
rect 117750 670980 117840 671220
rect 118080 670980 118170 671220
rect 118410 670980 118500 671220
rect 118740 670980 118850 671220
rect 119090 670980 119180 671220
rect 119420 670980 119510 671220
rect 119750 670980 119840 671220
rect 120080 670980 120190 671220
rect 120430 670980 120520 671220
rect 120760 670980 120850 671220
rect 121090 670980 121180 671220
rect 121420 670980 121530 671220
rect 121770 670980 122190 671220
rect 122430 670980 122520 671220
rect 122760 670980 122850 671220
rect 123090 670980 123180 671220
rect 123420 670980 123530 671220
rect 123770 670980 123860 671220
rect 124100 670980 124190 671220
rect 124430 670980 124520 671220
rect 124760 670980 124870 671220
rect 125110 670980 125200 671220
rect 125440 670980 125530 671220
rect 125770 670980 125860 671220
rect 126100 670980 126210 671220
rect 126450 670980 126540 671220
rect 126780 670980 126870 671220
rect 127110 670980 127200 671220
rect 127440 670980 127550 671220
rect 127790 670980 127880 671220
rect 128120 670980 128210 671220
rect 128450 670980 128540 671220
rect 128780 670980 128890 671220
rect 129130 670980 129220 671220
rect 129460 670980 129550 671220
rect 129790 670980 129880 671220
rect 130120 670980 130230 671220
rect 130470 670980 130560 671220
rect 130800 670980 130890 671220
rect 131130 670980 131220 671220
rect 131460 670980 131570 671220
rect 131810 670980 131900 671220
rect 132140 670980 132230 671220
rect 132470 670980 132560 671220
rect 132800 670980 132910 671220
rect 133150 670980 133570 671220
rect 133810 670980 133900 671220
rect 134140 670980 134230 671220
rect 134470 670980 134560 671220
rect 134800 670980 134910 671220
rect 135150 670980 135240 671220
rect 135480 670980 135570 671220
rect 135810 670980 135900 671220
rect 136140 670980 136250 671220
rect 136490 670980 136580 671220
rect 136820 670980 136910 671220
rect 137150 670980 137240 671220
rect 137480 670980 137590 671220
rect 137830 670980 137920 671220
rect 138160 670980 138250 671220
rect 138490 670980 138580 671220
rect 138820 670980 138930 671220
rect 139170 670980 139260 671220
rect 139500 670980 139590 671220
rect 139830 670980 139920 671220
rect 140160 670980 140270 671220
rect 140510 670980 140600 671220
rect 140840 670980 140930 671220
rect 141170 670980 141260 671220
rect 141500 670980 141610 671220
rect 141850 670980 141940 671220
rect 142180 670980 142270 671220
rect 142510 670980 142600 671220
rect 142840 670980 142950 671220
rect 143190 670980 143280 671220
rect 143520 670980 143610 671220
rect 143850 670980 143940 671220
rect 144180 670980 144290 671220
rect 144530 670980 144950 671220
rect 145190 670980 145280 671220
rect 145520 670980 145610 671220
rect 145850 670980 145940 671220
rect 146180 670980 146290 671220
rect 146530 670980 146620 671220
rect 146860 670980 146950 671220
rect 147190 670980 147280 671220
rect 147520 670980 147630 671220
rect 147870 670980 147960 671220
rect 148200 670980 148290 671220
rect 148530 670980 148620 671220
rect 148860 670980 148970 671220
rect 149210 670980 149300 671220
rect 149540 670980 149630 671220
rect 149870 670980 149960 671220
rect 150200 670980 150310 671220
rect 150550 670980 150640 671220
rect 150880 670980 150970 671220
rect 151210 670980 151300 671220
rect 151540 670980 151650 671220
rect 151890 670980 151980 671220
rect 152220 670980 152310 671220
rect 152550 670980 152640 671220
rect 152880 670980 152990 671220
rect 153230 670980 153320 671220
rect 153560 670980 153650 671220
rect 153890 670980 153980 671220
rect 154220 670980 154330 671220
rect 154570 670980 154660 671220
rect 154900 670980 154990 671220
rect 155230 670980 155320 671220
rect 155560 670980 155670 671220
rect 155910 670980 155960 671220
rect 110760 670890 155960 670980
rect 110760 670650 110810 670890
rect 111050 670650 111140 670890
rect 111380 670650 111470 670890
rect 111710 670650 111800 670890
rect 112040 670650 112150 670890
rect 112390 670650 112480 670890
rect 112720 670650 112810 670890
rect 113050 670650 113140 670890
rect 113380 670650 113490 670890
rect 113730 670650 113820 670890
rect 114060 670650 114150 670890
rect 114390 670650 114480 670890
rect 114720 670650 114830 670890
rect 115070 670650 115160 670890
rect 115400 670650 115490 670890
rect 115730 670650 115820 670890
rect 116060 670650 116170 670890
rect 116410 670650 116500 670890
rect 116740 670650 116830 670890
rect 117070 670650 117160 670890
rect 117400 670650 117510 670890
rect 117750 670650 117840 670890
rect 118080 670650 118170 670890
rect 118410 670650 118500 670890
rect 118740 670650 118850 670890
rect 119090 670650 119180 670890
rect 119420 670650 119510 670890
rect 119750 670650 119840 670890
rect 120080 670650 120190 670890
rect 120430 670650 120520 670890
rect 120760 670650 120850 670890
rect 121090 670650 121180 670890
rect 121420 670650 121530 670890
rect 121770 670650 122190 670890
rect 122430 670650 122520 670890
rect 122760 670650 122850 670890
rect 123090 670650 123180 670890
rect 123420 670650 123530 670890
rect 123770 670650 123860 670890
rect 124100 670650 124190 670890
rect 124430 670650 124520 670890
rect 124760 670650 124870 670890
rect 125110 670650 125200 670890
rect 125440 670650 125530 670890
rect 125770 670650 125860 670890
rect 126100 670650 126210 670890
rect 126450 670650 126540 670890
rect 126780 670650 126870 670890
rect 127110 670650 127200 670890
rect 127440 670650 127550 670890
rect 127790 670650 127880 670890
rect 128120 670650 128210 670890
rect 128450 670650 128540 670890
rect 128780 670650 128890 670890
rect 129130 670650 129220 670890
rect 129460 670650 129550 670890
rect 129790 670650 129880 670890
rect 130120 670650 130230 670890
rect 130470 670650 130560 670890
rect 130800 670650 130890 670890
rect 131130 670650 131220 670890
rect 131460 670650 131570 670890
rect 131810 670650 131900 670890
rect 132140 670650 132230 670890
rect 132470 670650 132560 670890
rect 132800 670650 132910 670890
rect 133150 670650 133570 670890
rect 133810 670650 133900 670890
rect 134140 670650 134230 670890
rect 134470 670650 134560 670890
rect 134800 670650 134910 670890
rect 135150 670650 135240 670890
rect 135480 670650 135570 670890
rect 135810 670650 135900 670890
rect 136140 670650 136250 670890
rect 136490 670650 136580 670890
rect 136820 670650 136910 670890
rect 137150 670650 137240 670890
rect 137480 670650 137590 670890
rect 137830 670650 137920 670890
rect 138160 670650 138250 670890
rect 138490 670650 138580 670890
rect 138820 670650 138930 670890
rect 139170 670650 139260 670890
rect 139500 670650 139590 670890
rect 139830 670650 139920 670890
rect 140160 670650 140270 670890
rect 140510 670650 140600 670890
rect 140840 670650 140930 670890
rect 141170 670650 141260 670890
rect 141500 670650 141610 670890
rect 141850 670650 141940 670890
rect 142180 670650 142270 670890
rect 142510 670650 142600 670890
rect 142840 670650 142950 670890
rect 143190 670650 143280 670890
rect 143520 670650 143610 670890
rect 143850 670650 143940 670890
rect 144180 670650 144290 670890
rect 144530 670650 144950 670890
rect 145190 670650 145280 670890
rect 145520 670650 145610 670890
rect 145850 670650 145940 670890
rect 146180 670650 146290 670890
rect 146530 670650 146620 670890
rect 146860 670650 146950 670890
rect 147190 670650 147280 670890
rect 147520 670650 147630 670890
rect 147870 670650 147960 670890
rect 148200 670650 148290 670890
rect 148530 670650 148620 670890
rect 148860 670650 148970 670890
rect 149210 670650 149300 670890
rect 149540 670650 149630 670890
rect 149870 670650 149960 670890
rect 150200 670650 150310 670890
rect 150550 670650 150640 670890
rect 150880 670650 150970 670890
rect 151210 670650 151300 670890
rect 151540 670650 151650 670890
rect 151890 670650 151980 670890
rect 152220 670650 152310 670890
rect 152550 670650 152640 670890
rect 152880 670650 152990 670890
rect 153230 670650 153320 670890
rect 153560 670650 153650 670890
rect 153890 670650 153980 670890
rect 154220 670650 154330 670890
rect 154570 670650 154660 670890
rect 154900 670650 154990 670890
rect 155230 670650 155320 670890
rect 155560 670650 155670 670890
rect 155910 670650 155960 670890
rect 110760 670560 155960 670650
rect 110760 670320 110810 670560
rect 111050 670320 111140 670560
rect 111380 670320 111470 670560
rect 111710 670320 111800 670560
rect 112040 670320 112150 670560
rect 112390 670320 112480 670560
rect 112720 670320 112810 670560
rect 113050 670320 113140 670560
rect 113380 670320 113490 670560
rect 113730 670320 113820 670560
rect 114060 670320 114150 670560
rect 114390 670320 114480 670560
rect 114720 670320 114830 670560
rect 115070 670320 115160 670560
rect 115400 670320 115490 670560
rect 115730 670320 115820 670560
rect 116060 670320 116170 670560
rect 116410 670320 116500 670560
rect 116740 670320 116830 670560
rect 117070 670320 117160 670560
rect 117400 670320 117510 670560
rect 117750 670320 117840 670560
rect 118080 670320 118170 670560
rect 118410 670320 118500 670560
rect 118740 670320 118850 670560
rect 119090 670320 119180 670560
rect 119420 670320 119510 670560
rect 119750 670320 119840 670560
rect 120080 670320 120190 670560
rect 120430 670320 120520 670560
rect 120760 670320 120850 670560
rect 121090 670320 121180 670560
rect 121420 670320 121530 670560
rect 121770 670320 122190 670560
rect 122430 670320 122520 670560
rect 122760 670320 122850 670560
rect 123090 670320 123180 670560
rect 123420 670320 123530 670560
rect 123770 670320 123860 670560
rect 124100 670320 124190 670560
rect 124430 670320 124520 670560
rect 124760 670320 124870 670560
rect 125110 670320 125200 670560
rect 125440 670320 125530 670560
rect 125770 670320 125860 670560
rect 126100 670320 126210 670560
rect 126450 670320 126540 670560
rect 126780 670320 126870 670560
rect 127110 670320 127200 670560
rect 127440 670320 127550 670560
rect 127790 670320 127880 670560
rect 128120 670320 128210 670560
rect 128450 670320 128540 670560
rect 128780 670320 128890 670560
rect 129130 670320 129220 670560
rect 129460 670320 129550 670560
rect 129790 670320 129880 670560
rect 130120 670320 130230 670560
rect 130470 670320 130560 670560
rect 130800 670320 130890 670560
rect 131130 670320 131220 670560
rect 131460 670320 131570 670560
rect 131810 670320 131900 670560
rect 132140 670320 132230 670560
rect 132470 670320 132560 670560
rect 132800 670320 132910 670560
rect 133150 670320 133570 670560
rect 133810 670320 133900 670560
rect 134140 670320 134230 670560
rect 134470 670320 134560 670560
rect 134800 670320 134910 670560
rect 135150 670320 135240 670560
rect 135480 670320 135570 670560
rect 135810 670320 135900 670560
rect 136140 670320 136250 670560
rect 136490 670320 136580 670560
rect 136820 670320 136910 670560
rect 137150 670320 137240 670560
rect 137480 670320 137590 670560
rect 137830 670320 137920 670560
rect 138160 670320 138250 670560
rect 138490 670320 138580 670560
rect 138820 670320 138930 670560
rect 139170 670320 139260 670560
rect 139500 670320 139590 670560
rect 139830 670320 139920 670560
rect 140160 670320 140270 670560
rect 140510 670320 140600 670560
rect 140840 670320 140930 670560
rect 141170 670320 141260 670560
rect 141500 670320 141610 670560
rect 141850 670320 141940 670560
rect 142180 670320 142270 670560
rect 142510 670320 142600 670560
rect 142840 670320 142950 670560
rect 143190 670320 143280 670560
rect 143520 670320 143610 670560
rect 143850 670320 143940 670560
rect 144180 670320 144290 670560
rect 144530 670320 144950 670560
rect 145190 670320 145280 670560
rect 145520 670320 145610 670560
rect 145850 670320 145940 670560
rect 146180 670320 146290 670560
rect 146530 670320 146620 670560
rect 146860 670320 146950 670560
rect 147190 670320 147280 670560
rect 147520 670320 147630 670560
rect 147870 670320 147960 670560
rect 148200 670320 148290 670560
rect 148530 670320 148620 670560
rect 148860 670320 148970 670560
rect 149210 670320 149300 670560
rect 149540 670320 149630 670560
rect 149870 670320 149960 670560
rect 150200 670320 150310 670560
rect 150550 670320 150640 670560
rect 150880 670320 150970 670560
rect 151210 670320 151300 670560
rect 151540 670320 151650 670560
rect 151890 670320 151980 670560
rect 152220 670320 152310 670560
rect 152550 670320 152640 670560
rect 152880 670320 152990 670560
rect 153230 670320 153320 670560
rect 153560 670320 153650 670560
rect 153890 670320 153980 670560
rect 154220 670320 154330 670560
rect 154570 670320 154660 670560
rect 154900 670320 154990 670560
rect 155230 670320 155320 670560
rect 155560 670320 155670 670560
rect 155910 670320 155960 670560
rect 110760 670210 155960 670320
rect 110760 669970 110810 670210
rect 111050 669970 111140 670210
rect 111380 669970 111470 670210
rect 111710 669970 111800 670210
rect 112040 669970 112150 670210
rect 112390 669970 112480 670210
rect 112720 669970 112810 670210
rect 113050 669970 113140 670210
rect 113380 669970 113490 670210
rect 113730 669970 113820 670210
rect 114060 669970 114150 670210
rect 114390 669970 114480 670210
rect 114720 669970 114830 670210
rect 115070 669970 115160 670210
rect 115400 669970 115490 670210
rect 115730 669970 115820 670210
rect 116060 669970 116170 670210
rect 116410 669970 116500 670210
rect 116740 669970 116830 670210
rect 117070 669970 117160 670210
rect 117400 669970 117510 670210
rect 117750 669970 117840 670210
rect 118080 669970 118170 670210
rect 118410 669970 118500 670210
rect 118740 669970 118850 670210
rect 119090 669970 119180 670210
rect 119420 669970 119510 670210
rect 119750 669970 119840 670210
rect 120080 669970 120190 670210
rect 120430 669970 120520 670210
rect 120760 669970 120850 670210
rect 121090 669970 121180 670210
rect 121420 669970 121530 670210
rect 121770 669970 122190 670210
rect 122430 669970 122520 670210
rect 122760 669970 122850 670210
rect 123090 669970 123180 670210
rect 123420 669970 123530 670210
rect 123770 669970 123860 670210
rect 124100 669970 124190 670210
rect 124430 669970 124520 670210
rect 124760 669970 124870 670210
rect 125110 669970 125200 670210
rect 125440 669970 125530 670210
rect 125770 669970 125860 670210
rect 126100 669970 126210 670210
rect 126450 669970 126540 670210
rect 126780 669970 126870 670210
rect 127110 669970 127200 670210
rect 127440 669970 127550 670210
rect 127790 669970 127880 670210
rect 128120 669970 128210 670210
rect 128450 669970 128540 670210
rect 128780 669970 128890 670210
rect 129130 669970 129220 670210
rect 129460 669970 129550 670210
rect 129790 669970 129880 670210
rect 130120 669970 130230 670210
rect 130470 669970 130560 670210
rect 130800 669970 130890 670210
rect 131130 669970 131220 670210
rect 131460 669970 131570 670210
rect 131810 669970 131900 670210
rect 132140 669970 132230 670210
rect 132470 669970 132560 670210
rect 132800 669970 132910 670210
rect 133150 669970 133570 670210
rect 133810 669970 133900 670210
rect 134140 669970 134230 670210
rect 134470 669970 134560 670210
rect 134800 669970 134910 670210
rect 135150 669970 135240 670210
rect 135480 669970 135570 670210
rect 135810 669970 135900 670210
rect 136140 669970 136250 670210
rect 136490 669970 136580 670210
rect 136820 669970 136910 670210
rect 137150 669970 137240 670210
rect 137480 669970 137590 670210
rect 137830 669970 137920 670210
rect 138160 669970 138250 670210
rect 138490 669970 138580 670210
rect 138820 669970 138930 670210
rect 139170 669970 139260 670210
rect 139500 669970 139590 670210
rect 139830 669970 139920 670210
rect 140160 669970 140270 670210
rect 140510 669970 140600 670210
rect 140840 669970 140930 670210
rect 141170 669970 141260 670210
rect 141500 669970 141610 670210
rect 141850 669970 141940 670210
rect 142180 669970 142270 670210
rect 142510 669970 142600 670210
rect 142840 669970 142950 670210
rect 143190 669970 143280 670210
rect 143520 669970 143610 670210
rect 143850 669970 143940 670210
rect 144180 669970 144290 670210
rect 144530 669970 144950 670210
rect 145190 669970 145280 670210
rect 145520 669970 145610 670210
rect 145850 669970 145940 670210
rect 146180 669970 146290 670210
rect 146530 669970 146620 670210
rect 146860 669970 146950 670210
rect 147190 669970 147280 670210
rect 147520 669970 147630 670210
rect 147870 669970 147960 670210
rect 148200 669970 148290 670210
rect 148530 669970 148620 670210
rect 148860 669970 148970 670210
rect 149210 669970 149300 670210
rect 149540 669970 149630 670210
rect 149870 669970 149960 670210
rect 150200 669970 150310 670210
rect 150550 669970 150640 670210
rect 150880 669970 150970 670210
rect 151210 669970 151300 670210
rect 151540 669970 151650 670210
rect 151890 669970 151980 670210
rect 152220 669970 152310 670210
rect 152550 669970 152640 670210
rect 152880 669970 152990 670210
rect 153230 669970 153320 670210
rect 153560 669970 153650 670210
rect 153890 669970 153980 670210
rect 154220 669970 154330 670210
rect 154570 669970 154660 670210
rect 154900 669970 154990 670210
rect 155230 669970 155320 670210
rect 155560 669970 155670 670210
rect 155910 669970 155960 670210
rect 110760 669880 155960 669970
rect 110760 669640 110810 669880
rect 111050 669640 111140 669880
rect 111380 669640 111470 669880
rect 111710 669640 111800 669880
rect 112040 669640 112150 669880
rect 112390 669640 112480 669880
rect 112720 669640 112810 669880
rect 113050 669640 113140 669880
rect 113380 669640 113490 669880
rect 113730 669640 113820 669880
rect 114060 669640 114150 669880
rect 114390 669640 114480 669880
rect 114720 669640 114830 669880
rect 115070 669640 115160 669880
rect 115400 669640 115490 669880
rect 115730 669640 115820 669880
rect 116060 669640 116170 669880
rect 116410 669640 116500 669880
rect 116740 669640 116830 669880
rect 117070 669640 117160 669880
rect 117400 669640 117510 669880
rect 117750 669640 117840 669880
rect 118080 669640 118170 669880
rect 118410 669640 118500 669880
rect 118740 669640 118850 669880
rect 119090 669640 119180 669880
rect 119420 669640 119510 669880
rect 119750 669640 119840 669880
rect 120080 669640 120190 669880
rect 120430 669640 120520 669880
rect 120760 669640 120850 669880
rect 121090 669640 121180 669880
rect 121420 669640 121530 669880
rect 121770 669640 122190 669880
rect 122430 669640 122520 669880
rect 122760 669640 122850 669880
rect 123090 669640 123180 669880
rect 123420 669640 123530 669880
rect 123770 669640 123860 669880
rect 124100 669640 124190 669880
rect 124430 669640 124520 669880
rect 124760 669640 124870 669880
rect 125110 669640 125200 669880
rect 125440 669640 125530 669880
rect 125770 669640 125860 669880
rect 126100 669640 126210 669880
rect 126450 669640 126540 669880
rect 126780 669640 126870 669880
rect 127110 669640 127200 669880
rect 127440 669640 127550 669880
rect 127790 669640 127880 669880
rect 128120 669640 128210 669880
rect 128450 669640 128540 669880
rect 128780 669640 128890 669880
rect 129130 669640 129220 669880
rect 129460 669640 129550 669880
rect 129790 669640 129880 669880
rect 130120 669640 130230 669880
rect 130470 669640 130560 669880
rect 130800 669640 130890 669880
rect 131130 669640 131220 669880
rect 131460 669640 131570 669880
rect 131810 669640 131900 669880
rect 132140 669640 132230 669880
rect 132470 669640 132560 669880
rect 132800 669640 132910 669880
rect 133150 669640 133570 669880
rect 133810 669640 133900 669880
rect 134140 669640 134230 669880
rect 134470 669640 134560 669880
rect 134800 669640 134910 669880
rect 135150 669640 135240 669880
rect 135480 669640 135570 669880
rect 135810 669640 135900 669880
rect 136140 669640 136250 669880
rect 136490 669640 136580 669880
rect 136820 669640 136910 669880
rect 137150 669640 137240 669880
rect 137480 669640 137590 669880
rect 137830 669640 137920 669880
rect 138160 669640 138250 669880
rect 138490 669640 138580 669880
rect 138820 669640 138930 669880
rect 139170 669640 139260 669880
rect 139500 669640 139590 669880
rect 139830 669640 139920 669880
rect 140160 669640 140270 669880
rect 140510 669640 140600 669880
rect 140840 669640 140930 669880
rect 141170 669640 141260 669880
rect 141500 669640 141610 669880
rect 141850 669640 141940 669880
rect 142180 669640 142270 669880
rect 142510 669640 142600 669880
rect 142840 669640 142950 669880
rect 143190 669640 143280 669880
rect 143520 669640 143610 669880
rect 143850 669640 143940 669880
rect 144180 669640 144290 669880
rect 144530 669640 144950 669880
rect 145190 669640 145280 669880
rect 145520 669640 145610 669880
rect 145850 669640 145940 669880
rect 146180 669640 146290 669880
rect 146530 669640 146620 669880
rect 146860 669640 146950 669880
rect 147190 669640 147280 669880
rect 147520 669640 147630 669880
rect 147870 669640 147960 669880
rect 148200 669640 148290 669880
rect 148530 669640 148620 669880
rect 148860 669640 148970 669880
rect 149210 669640 149300 669880
rect 149540 669640 149630 669880
rect 149870 669640 149960 669880
rect 150200 669640 150310 669880
rect 150550 669640 150640 669880
rect 150880 669640 150970 669880
rect 151210 669640 151300 669880
rect 151540 669640 151650 669880
rect 151890 669640 151980 669880
rect 152220 669640 152310 669880
rect 152550 669640 152640 669880
rect 152880 669640 152990 669880
rect 153230 669640 153320 669880
rect 153560 669640 153650 669880
rect 153890 669640 153980 669880
rect 154220 669640 154330 669880
rect 154570 669640 154660 669880
rect 154900 669640 154990 669880
rect 155230 669640 155320 669880
rect 155560 669640 155670 669880
rect 155910 669640 155960 669880
rect 110760 669550 155960 669640
rect 110760 669310 110810 669550
rect 111050 669310 111140 669550
rect 111380 669310 111470 669550
rect 111710 669310 111800 669550
rect 112040 669310 112150 669550
rect 112390 669310 112480 669550
rect 112720 669310 112810 669550
rect 113050 669310 113140 669550
rect 113380 669310 113490 669550
rect 113730 669310 113820 669550
rect 114060 669310 114150 669550
rect 114390 669310 114480 669550
rect 114720 669310 114830 669550
rect 115070 669310 115160 669550
rect 115400 669310 115490 669550
rect 115730 669310 115820 669550
rect 116060 669310 116170 669550
rect 116410 669310 116500 669550
rect 116740 669310 116830 669550
rect 117070 669310 117160 669550
rect 117400 669310 117510 669550
rect 117750 669310 117840 669550
rect 118080 669310 118170 669550
rect 118410 669310 118500 669550
rect 118740 669310 118850 669550
rect 119090 669310 119180 669550
rect 119420 669310 119510 669550
rect 119750 669310 119840 669550
rect 120080 669310 120190 669550
rect 120430 669310 120520 669550
rect 120760 669310 120850 669550
rect 121090 669310 121180 669550
rect 121420 669310 121530 669550
rect 121770 669310 122190 669550
rect 122430 669310 122520 669550
rect 122760 669310 122850 669550
rect 123090 669310 123180 669550
rect 123420 669310 123530 669550
rect 123770 669310 123860 669550
rect 124100 669310 124190 669550
rect 124430 669310 124520 669550
rect 124760 669310 124870 669550
rect 125110 669310 125200 669550
rect 125440 669310 125530 669550
rect 125770 669310 125860 669550
rect 126100 669310 126210 669550
rect 126450 669310 126540 669550
rect 126780 669310 126870 669550
rect 127110 669310 127200 669550
rect 127440 669310 127550 669550
rect 127790 669310 127880 669550
rect 128120 669310 128210 669550
rect 128450 669310 128540 669550
rect 128780 669310 128890 669550
rect 129130 669310 129220 669550
rect 129460 669310 129550 669550
rect 129790 669310 129880 669550
rect 130120 669310 130230 669550
rect 130470 669310 130560 669550
rect 130800 669310 130890 669550
rect 131130 669310 131220 669550
rect 131460 669310 131570 669550
rect 131810 669310 131900 669550
rect 132140 669310 132230 669550
rect 132470 669310 132560 669550
rect 132800 669310 132910 669550
rect 133150 669310 133570 669550
rect 133810 669310 133900 669550
rect 134140 669310 134230 669550
rect 134470 669310 134560 669550
rect 134800 669310 134910 669550
rect 135150 669310 135240 669550
rect 135480 669310 135570 669550
rect 135810 669310 135900 669550
rect 136140 669310 136250 669550
rect 136490 669310 136580 669550
rect 136820 669310 136910 669550
rect 137150 669310 137240 669550
rect 137480 669310 137590 669550
rect 137830 669310 137920 669550
rect 138160 669310 138250 669550
rect 138490 669310 138580 669550
rect 138820 669310 138930 669550
rect 139170 669310 139260 669550
rect 139500 669310 139590 669550
rect 139830 669310 139920 669550
rect 140160 669310 140270 669550
rect 140510 669310 140600 669550
rect 140840 669310 140930 669550
rect 141170 669310 141260 669550
rect 141500 669310 141610 669550
rect 141850 669310 141940 669550
rect 142180 669310 142270 669550
rect 142510 669310 142600 669550
rect 142840 669310 142950 669550
rect 143190 669310 143280 669550
rect 143520 669310 143610 669550
rect 143850 669310 143940 669550
rect 144180 669310 144290 669550
rect 144530 669310 144950 669550
rect 145190 669310 145280 669550
rect 145520 669310 145610 669550
rect 145850 669310 145940 669550
rect 146180 669310 146290 669550
rect 146530 669310 146620 669550
rect 146860 669310 146950 669550
rect 147190 669310 147280 669550
rect 147520 669310 147630 669550
rect 147870 669310 147960 669550
rect 148200 669310 148290 669550
rect 148530 669310 148620 669550
rect 148860 669310 148970 669550
rect 149210 669310 149300 669550
rect 149540 669310 149630 669550
rect 149870 669310 149960 669550
rect 150200 669310 150310 669550
rect 150550 669310 150640 669550
rect 150880 669310 150970 669550
rect 151210 669310 151300 669550
rect 151540 669310 151650 669550
rect 151890 669310 151980 669550
rect 152220 669310 152310 669550
rect 152550 669310 152640 669550
rect 152880 669310 152990 669550
rect 153230 669310 153320 669550
rect 153560 669310 153650 669550
rect 153890 669310 153980 669550
rect 154220 669310 154330 669550
rect 154570 669310 154660 669550
rect 154900 669310 154990 669550
rect 155230 669310 155320 669550
rect 155560 669310 155670 669550
rect 155910 669310 155960 669550
rect 110760 669220 155960 669310
rect 110760 668980 110810 669220
rect 111050 668980 111140 669220
rect 111380 668980 111470 669220
rect 111710 668980 111800 669220
rect 112040 668980 112150 669220
rect 112390 668980 112480 669220
rect 112720 668980 112810 669220
rect 113050 668980 113140 669220
rect 113380 668980 113490 669220
rect 113730 668980 113820 669220
rect 114060 668980 114150 669220
rect 114390 668980 114480 669220
rect 114720 668980 114830 669220
rect 115070 668980 115160 669220
rect 115400 668980 115490 669220
rect 115730 668980 115820 669220
rect 116060 668980 116170 669220
rect 116410 668980 116500 669220
rect 116740 668980 116830 669220
rect 117070 668980 117160 669220
rect 117400 668980 117510 669220
rect 117750 668980 117840 669220
rect 118080 668980 118170 669220
rect 118410 668980 118500 669220
rect 118740 668980 118850 669220
rect 119090 668980 119180 669220
rect 119420 668980 119510 669220
rect 119750 668980 119840 669220
rect 120080 668980 120190 669220
rect 120430 668980 120520 669220
rect 120760 668980 120850 669220
rect 121090 668980 121180 669220
rect 121420 668980 121530 669220
rect 121770 668980 122190 669220
rect 122430 668980 122520 669220
rect 122760 668980 122850 669220
rect 123090 668980 123180 669220
rect 123420 668980 123530 669220
rect 123770 668980 123860 669220
rect 124100 668980 124190 669220
rect 124430 668980 124520 669220
rect 124760 668980 124870 669220
rect 125110 668980 125200 669220
rect 125440 668980 125530 669220
rect 125770 668980 125860 669220
rect 126100 668980 126210 669220
rect 126450 668980 126540 669220
rect 126780 668980 126870 669220
rect 127110 668980 127200 669220
rect 127440 668980 127550 669220
rect 127790 668980 127880 669220
rect 128120 668980 128210 669220
rect 128450 668980 128540 669220
rect 128780 668980 128890 669220
rect 129130 668980 129220 669220
rect 129460 668980 129550 669220
rect 129790 668980 129880 669220
rect 130120 668980 130230 669220
rect 130470 668980 130560 669220
rect 130800 668980 130890 669220
rect 131130 668980 131220 669220
rect 131460 668980 131570 669220
rect 131810 668980 131900 669220
rect 132140 668980 132230 669220
rect 132470 668980 132560 669220
rect 132800 668980 132910 669220
rect 133150 668980 133570 669220
rect 133810 668980 133900 669220
rect 134140 668980 134230 669220
rect 134470 668980 134560 669220
rect 134800 668980 134910 669220
rect 135150 668980 135240 669220
rect 135480 668980 135570 669220
rect 135810 668980 135900 669220
rect 136140 668980 136250 669220
rect 136490 668980 136580 669220
rect 136820 668980 136910 669220
rect 137150 668980 137240 669220
rect 137480 668980 137590 669220
rect 137830 668980 137920 669220
rect 138160 668980 138250 669220
rect 138490 668980 138580 669220
rect 138820 668980 138930 669220
rect 139170 668980 139260 669220
rect 139500 668980 139590 669220
rect 139830 668980 139920 669220
rect 140160 668980 140270 669220
rect 140510 668980 140600 669220
rect 140840 668980 140930 669220
rect 141170 668980 141260 669220
rect 141500 668980 141610 669220
rect 141850 668980 141940 669220
rect 142180 668980 142270 669220
rect 142510 668980 142600 669220
rect 142840 668980 142950 669220
rect 143190 668980 143280 669220
rect 143520 668980 143610 669220
rect 143850 668980 143940 669220
rect 144180 668980 144290 669220
rect 144530 668980 144950 669220
rect 145190 668980 145280 669220
rect 145520 668980 145610 669220
rect 145850 668980 145940 669220
rect 146180 668980 146290 669220
rect 146530 668980 146620 669220
rect 146860 668980 146950 669220
rect 147190 668980 147280 669220
rect 147520 668980 147630 669220
rect 147870 668980 147960 669220
rect 148200 668980 148290 669220
rect 148530 668980 148620 669220
rect 148860 668980 148970 669220
rect 149210 668980 149300 669220
rect 149540 668980 149630 669220
rect 149870 668980 149960 669220
rect 150200 668980 150310 669220
rect 150550 668980 150640 669220
rect 150880 668980 150970 669220
rect 151210 668980 151300 669220
rect 151540 668980 151650 669220
rect 151890 668980 151980 669220
rect 152220 668980 152310 669220
rect 152550 668980 152640 669220
rect 152880 668980 152990 669220
rect 153230 668980 153320 669220
rect 153560 668980 153650 669220
rect 153890 668980 153980 669220
rect 154220 668980 154330 669220
rect 154570 668980 154660 669220
rect 154900 668980 154990 669220
rect 155230 668980 155320 669220
rect 155560 668980 155670 669220
rect 155910 668980 155960 669220
rect 110760 668870 155960 668980
rect 110760 668630 110810 668870
rect 111050 668630 111140 668870
rect 111380 668630 111470 668870
rect 111710 668630 111800 668870
rect 112040 668630 112150 668870
rect 112390 668630 112480 668870
rect 112720 668630 112810 668870
rect 113050 668630 113140 668870
rect 113380 668630 113490 668870
rect 113730 668630 113820 668870
rect 114060 668630 114150 668870
rect 114390 668630 114480 668870
rect 114720 668630 114830 668870
rect 115070 668630 115160 668870
rect 115400 668630 115490 668870
rect 115730 668630 115820 668870
rect 116060 668630 116170 668870
rect 116410 668630 116500 668870
rect 116740 668630 116830 668870
rect 117070 668630 117160 668870
rect 117400 668630 117510 668870
rect 117750 668630 117840 668870
rect 118080 668630 118170 668870
rect 118410 668630 118500 668870
rect 118740 668630 118850 668870
rect 119090 668630 119180 668870
rect 119420 668630 119510 668870
rect 119750 668630 119840 668870
rect 120080 668630 120190 668870
rect 120430 668630 120520 668870
rect 120760 668630 120850 668870
rect 121090 668630 121180 668870
rect 121420 668630 121530 668870
rect 121770 668630 122190 668870
rect 122430 668630 122520 668870
rect 122760 668630 122850 668870
rect 123090 668630 123180 668870
rect 123420 668630 123530 668870
rect 123770 668630 123860 668870
rect 124100 668630 124190 668870
rect 124430 668630 124520 668870
rect 124760 668630 124870 668870
rect 125110 668630 125200 668870
rect 125440 668630 125530 668870
rect 125770 668630 125860 668870
rect 126100 668630 126210 668870
rect 126450 668630 126540 668870
rect 126780 668630 126870 668870
rect 127110 668630 127200 668870
rect 127440 668630 127550 668870
rect 127790 668630 127880 668870
rect 128120 668630 128210 668870
rect 128450 668630 128540 668870
rect 128780 668630 128890 668870
rect 129130 668630 129220 668870
rect 129460 668630 129550 668870
rect 129790 668630 129880 668870
rect 130120 668630 130230 668870
rect 130470 668630 130560 668870
rect 130800 668630 130890 668870
rect 131130 668630 131220 668870
rect 131460 668630 131570 668870
rect 131810 668630 131900 668870
rect 132140 668630 132230 668870
rect 132470 668630 132560 668870
rect 132800 668630 132910 668870
rect 133150 668630 133570 668870
rect 133810 668630 133900 668870
rect 134140 668630 134230 668870
rect 134470 668630 134560 668870
rect 134800 668630 134910 668870
rect 135150 668630 135240 668870
rect 135480 668630 135570 668870
rect 135810 668630 135900 668870
rect 136140 668630 136250 668870
rect 136490 668630 136580 668870
rect 136820 668630 136910 668870
rect 137150 668630 137240 668870
rect 137480 668630 137590 668870
rect 137830 668630 137920 668870
rect 138160 668630 138250 668870
rect 138490 668630 138580 668870
rect 138820 668630 138930 668870
rect 139170 668630 139260 668870
rect 139500 668630 139590 668870
rect 139830 668630 139920 668870
rect 140160 668630 140270 668870
rect 140510 668630 140600 668870
rect 140840 668630 140930 668870
rect 141170 668630 141260 668870
rect 141500 668630 141610 668870
rect 141850 668630 141940 668870
rect 142180 668630 142270 668870
rect 142510 668630 142600 668870
rect 142840 668630 142950 668870
rect 143190 668630 143280 668870
rect 143520 668630 143610 668870
rect 143850 668630 143940 668870
rect 144180 668630 144290 668870
rect 144530 668630 144950 668870
rect 145190 668630 145280 668870
rect 145520 668630 145610 668870
rect 145850 668630 145940 668870
rect 146180 668630 146290 668870
rect 146530 668630 146620 668870
rect 146860 668630 146950 668870
rect 147190 668630 147280 668870
rect 147520 668630 147630 668870
rect 147870 668630 147960 668870
rect 148200 668630 148290 668870
rect 148530 668630 148620 668870
rect 148860 668630 148970 668870
rect 149210 668630 149300 668870
rect 149540 668630 149630 668870
rect 149870 668630 149960 668870
rect 150200 668630 150310 668870
rect 150550 668630 150640 668870
rect 150880 668630 150970 668870
rect 151210 668630 151300 668870
rect 151540 668630 151650 668870
rect 151890 668630 151980 668870
rect 152220 668630 152310 668870
rect 152550 668630 152640 668870
rect 152880 668630 152990 668870
rect 153230 668630 153320 668870
rect 153560 668630 153650 668870
rect 153890 668630 153980 668870
rect 154220 668630 154330 668870
rect 154570 668630 154660 668870
rect 154900 668630 154990 668870
rect 155230 668630 155320 668870
rect 155560 668630 155670 668870
rect 155910 668630 155960 668870
rect 110760 668540 155960 668630
rect 110760 668300 110810 668540
rect 111050 668300 111140 668540
rect 111380 668300 111470 668540
rect 111710 668300 111800 668540
rect 112040 668300 112150 668540
rect 112390 668300 112480 668540
rect 112720 668300 112810 668540
rect 113050 668300 113140 668540
rect 113380 668300 113490 668540
rect 113730 668300 113820 668540
rect 114060 668300 114150 668540
rect 114390 668300 114480 668540
rect 114720 668300 114830 668540
rect 115070 668300 115160 668540
rect 115400 668300 115490 668540
rect 115730 668300 115820 668540
rect 116060 668300 116170 668540
rect 116410 668300 116500 668540
rect 116740 668300 116830 668540
rect 117070 668300 117160 668540
rect 117400 668300 117510 668540
rect 117750 668300 117840 668540
rect 118080 668300 118170 668540
rect 118410 668300 118500 668540
rect 118740 668300 118850 668540
rect 119090 668300 119180 668540
rect 119420 668300 119510 668540
rect 119750 668300 119840 668540
rect 120080 668300 120190 668540
rect 120430 668300 120520 668540
rect 120760 668300 120850 668540
rect 121090 668300 121180 668540
rect 121420 668300 121530 668540
rect 121770 668300 122190 668540
rect 122430 668300 122520 668540
rect 122760 668300 122850 668540
rect 123090 668300 123180 668540
rect 123420 668300 123530 668540
rect 123770 668300 123860 668540
rect 124100 668300 124190 668540
rect 124430 668300 124520 668540
rect 124760 668300 124870 668540
rect 125110 668300 125200 668540
rect 125440 668300 125530 668540
rect 125770 668300 125860 668540
rect 126100 668300 126210 668540
rect 126450 668300 126540 668540
rect 126780 668300 126870 668540
rect 127110 668300 127200 668540
rect 127440 668300 127550 668540
rect 127790 668300 127880 668540
rect 128120 668300 128210 668540
rect 128450 668300 128540 668540
rect 128780 668300 128890 668540
rect 129130 668300 129220 668540
rect 129460 668300 129550 668540
rect 129790 668300 129880 668540
rect 130120 668300 130230 668540
rect 130470 668300 130560 668540
rect 130800 668300 130890 668540
rect 131130 668300 131220 668540
rect 131460 668300 131570 668540
rect 131810 668300 131900 668540
rect 132140 668300 132230 668540
rect 132470 668300 132560 668540
rect 132800 668300 132910 668540
rect 133150 668300 133570 668540
rect 133810 668300 133900 668540
rect 134140 668300 134230 668540
rect 134470 668300 134560 668540
rect 134800 668300 134910 668540
rect 135150 668300 135240 668540
rect 135480 668300 135570 668540
rect 135810 668300 135900 668540
rect 136140 668300 136250 668540
rect 136490 668300 136580 668540
rect 136820 668300 136910 668540
rect 137150 668300 137240 668540
rect 137480 668300 137590 668540
rect 137830 668300 137920 668540
rect 138160 668300 138250 668540
rect 138490 668300 138580 668540
rect 138820 668300 138930 668540
rect 139170 668300 139260 668540
rect 139500 668300 139590 668540
rect 139830 668300 139920 668540
rect 140160 668300 140270 668540
rect 140510 668300 140600 668540
rect 140840 668300 140930 668540
rect 141170 668300 141260 668540
rect 141500 668300 141610 668540
rect 141850 668300 141940 668540
rect 142180 668300 142270 668540
rect 142510 668300 142600 668540
rect 142840 668300 142950 668540
rect 143190 668300 143280 668540
rect 143520 668300 143610 668540
rect 143850 668300 143940 668540
rect 144180 668300 144290 668540
rect 144530 668300 144950 668540
rect 145190 668300 145280 668540
rect 145520 668300 145610 668540
rect 145850 668300 145940 668540
rect 146180 668300 146290 668540
rect 146530 668300 146620 668540
rect 146860 668300 146950 668540
rect 147190 668300 147280 668540
rect 147520 668300 147630 668540
rect 147870 668300 147960 668540
rect 148200 668300 148290 668540
rect 148530 668300 148620 668540
rect 148860 668300 148970 668540
rect 149210 668300 149300 668540
rect 149540 668300 149630 668540
rect 149870 668300 149960 668540
rect 150200 668300 150310 668540
rect 150550 668300 150640 668540
rect 150880 668300 150970 668540
rect 151210 668300 151300 668540
rect 151540 668300 151650 668540
rect 151890 668300 151980 668540
rect 152220 668300 152310 668540
rect 152550 668300 152640 668540
rect 152880 668300 152990 668540
rect 153230 668300 153320 668540
rect 153560 668300 153650 668540
rect 153890 668300 153980 668540
rect 154220 668300 154330 668540
rect 154570 668300 154660 668540
rect 154900 668300 154990 668540
rect 155230 668300 155320 668540
rect 155560 668300 155670 668540
rect 155910 668300 155960 668540
rect 110760 668210 155960 668300
rect 110760 667970 110810 668210
rect 111050 667970 111140 668210
rect 111380 667970 111470 668210
rect 111710 667970 111800 668210
rect 112040 667970 112150 668210
rect 112390 667970 112480 668210
rect 112720 667970 112810 668210
rect 113050 667970 113140 668210
rect 113380 667970 113490 668210
rect 113730 667970 113820 668210
rect 114060 667970 114150 668210
rect 114390 667970 114480 668210
rect 114720 667970 114830 668210
rect 115070 667970 115160 668210
rect 115400 667970 115490 668210
rect 115730 667970 115820 668210
rect 116060 667970 116170 668210
rect 116410 667970 116500 668210
rect 116740 667970 116830 668210
rect 117070 667970 117160 668210
rect 117400 667970 117510 668210
rect 117750 667970 117840 668210
rect 118080 667970 118170 668210
rect 118410 667970 118500 668210
rect 118740 667970 118850 668210
rect 119090 667970 119180 668210
rect 119420 667970 119510 668210
rect 119750 667970 119840 668210
rect 120080 667970 120190 668210
rect 120430 667970 120520 668210
rect 120760 667970 120850 668210
rect 121090 667970 121180 668210
rect 121420 667970 121530 668210
rect 121770 667970 122190 668210
rect 122430 667970 122520 668210
rect 122760 667970 122850 668210
rect 123090 667970 123180 668210
rect 123420 667970 123530 668210
rect 123770 667970 123860 668210
rect 124100 667970 124190 668210
rect 124430 667970 124520 668210
rect 124760 667970 124870 668210
rect 125110 667970 125200 668210
rect 125440 667970 125530 668210
rect 125770 667970 125860 668210
rect 126100 667970 126210 668210
rect 126450 667970 126540 668210
rect 126780 667970 126870 668210
rect 127110 667970 127200 668210
rect 127440 667970 127550 668210
rect 127790 667970 127880 668210
rect 128120 667970 128210 668210
rect 128450 667970 128540 668210
rect 128780 667970 128890 668210
rect 129130 667970 129220 668210
rect 129460 667970 129550 668210
rect 129790 667970 129880 668210
rect 130120 667970 130230 668210
rect 130470 667970 130560 668210
rect 130800 667970 130890 668210
rect 131130 667970 131220 668210
rect 131460 667970 131570 668210
rect 131810 667970 131900 668210
rect 132140 667970 132230 668210
rect 132470 667970 132560 668210
rect 132800 667970 132910 668210
rect 133150 667970 133570 668210
rect 133810 667970 133900 668210
rect 134140 667970 134230 668210
rect 134470 667970 134560 668210
rect 134800 667970 134910 668210
rect 135150 667970 135240 668210
rect 135480 667970 135570 668210
rect 135810 667970 135900 668210
rect 136140 667970 136250 668210
rect 136490 667970 136580 668210
rect 136820 667970 136910 668210
rect 137150 667970 137240 668210
rect 137480 667970 137590 668210
rect 137830 667970 137920 668210
rect 138160 667970 138250 668210
rect 138490 667970 138580 668210
rect 138820 667970 138930 668210
rect 139170 667970 139260 668210
rect 139500 667970 139590 668210
rect 139830 667970 139920 668210
rect 140160 667970 140270 668210
rect 140510 667970 140600 668210
rect 140840 667970 140930 668210
rect 141170 667970 141260 668210
rect 141500 667970 141610 668210
rect 141850 667970 141940 668210
rect 142180 667970 142270 668210
rect 142510 667970 142600 668210
rect 142840 667970 142950 668210
rect 143190 667970 143280 668210
rect 143520 667970 143610 668210
rect 143850 667970 143940 668210
rect 144180 667970 144290 668210
rect 144530 667970 144950 668210
rect 145190 667970 145280 668210
rect 145520 667970 145610 668210
rect 145850 667970 145940 668210
rect 146180 667970 146290 668210
rect 146530 667970 146620 668210
rect 146860 667970 146950 668210
rect 147190 667970 147280 668210
rect 147520 667970 147630 668210
rect 147870 667970 147960 668210
rect 148200 667970 148290 668210
rect 148530 667970 148620 668210
rect 148860 667970 148970 668210
rect 149210 667970 149300 668210
rect 149540 667970 149630 668210
rect 149870 667970 149960 668210
rect 150200 667970 150310 668210
rect 150550 667970 150640 668210
rect 150880 667970 150970 668210
rect 151210 667970 151300 668210
rect 151540 667970 151650 668210
rect 151890 667970 151980 668210
rect 152220 667970 152310 668210
rect 152550 667970 152640 668210
rect 152880 667970 152990 668210
rect 153230 667970 153320 668210
rect 153560 667970 153650 668210
rect 153890 667970 153980 668210
rect 154220 667970 154330 668210
rect 154570 667970 154660 668210
rect 154900 667970 154990 668210
rect 155230 667970 155320 668210
rect 155560 667970 155670 668210
rect 155910 667970 155960 668210
rect 110760 667880 155960 667970
rect 110760 667640 110810 667880
rect 111050 667640 111140 667880
rect 111380 667640 111470 667880
rect 111710 667640 111800 667880
rect 112040 667640 112150 667880
rect 112390 667640 112480 667880
rect 112720 667640 112810 667880
rect 113050 667640 113140 667880
rect 113380 667640 113490 667880
rect 113730 667640 113820 667880
rect 114060 667640 114150 667880
rect 114390 667640 114480 667880
rect 114720 667640 114830 667880
rect 115070 667640 115160 667880
rect 115400 667640 115490 667880
rect 115730 667640 115820 667880
rect 116060 667640 116170 667880
rect 116410 667640 116500 667880
rect 116740 667640 116830 667880
rect 117070 667640 117160 667880
rect 117400 667640 117510 667880
rect 117750 667640 117840 667880
rect 118080 667640 118170 667880
rect 118410 667640 118500 667880
rect 118740 667640 118850 667880
rect 119090 667640 119180 667880
rect 119420 667640 119510 667880
rect 119750 667640 119840 667880
rect 120080 667640 120190 667880
rect 120430 667640 120520 667880
rect 120760 667640 120850 667880
rect 121090 667640 121180 667880
rect 121420 667640 121530 667880
rect 121770 667640 122190 667880
rect 122430 667640 122520 667880
rect 122760 667640 122850 667880
rect 123090 667640 123180 667880
rect 123420 667640 123530 667880
rect 123770 667640 123860 667880
rect 124100 667640 124190 667880
rect 124430 667640 124520 667880
rect 124760 667640 124870 667880
rect 125110 667640 125200 667880
rect 125440 667640 125530 667880
rect 125770 667640 125860 667880
rect 126100 667640 126210 667880
rect 126450 667640 126540 667880
rect 126780 667640 126870 667880
rect 127110 667640 127200 667880
rect 127440 667640 127550 667880
rect 127790 667640 127880 667880
rect 128120 667640 128210 667880
rect 128450 667640 128540 667880
rect 128780 667640 128890 667880
rect 129130 667640 129220 667880
rect 129460 667640 129550 667880
rect 129790 667640 129880 667880
rect 130120 667640 130230 667880
rect 130470 667640 130560 667880
rect 130800 667640 130890 667880
rect 131130 667640 131220 667880
rect 131460 667640 131570 667880
rect 131810 667640 131900 667880
rect 132140 667640 132230 667880
rect 132470 667640 132560 667880
rect 132800 667640 132910 667880
rect 133150 667640 133570 667880
rect 133810 667640 133900 667880
rect 134140 667640 134230 667880
rect 134470 667640 134560 667880
rect 134800 667640 134910 667880
rect 135150 667640 135240 667880
rect 135480 667640 135570 667880
rect 135810 667640 135900 667880
rect 136140 667640 136250 667880
rect 136490 667640 136580 667880
rect 136820 667640 136910 667880
rect 137150 667640 137240 667880
rect 137480 667640 137590 667880
rect 137830 667640 137920 667880
rect 138160 667640 138250 667880
rect 138490 667640 138580 667880
rect 138820 667640 138930 667880
rect 139170 667640 139260 667880
rect 139500 667640 139590 667880
rect 139830 667640 139920 667880
rect 140160 667640 140270 667880
rect 140510 667640 140600 667880
rect 140840 667640 140930 667880
rect 141170 667640 141260 667880
rect 141500 667640 141610 667880
rect 141850 667640 141940 667880
rect 142180 667640 142270 667880
rect 142510 667640 142600 667880
rect 142840 667640 142950 667880
rect 143190 667640 143280 667880
rect 143520 667640 143610 667880
rect 143850 667640 143940 667880
rect 144180 667640 144290 667880
rect 144530 667640 144950 667880
rect 145190 667640 145280 667880
rect 145520 667640 145610 667880
rect 145850 667640 145940 667880
rect 146180 667640 146290 667880
rect 146530 667640 146620 667880
rect 146860 667640 146950 667880
rect 147190 667640 147280 667880
rect 147520 667640 147630 667880
rect 147870 667640 147960 667880
rect 148200 667640 148290 667880
rect 148530 667640 148620 667880
rect 148860 667640 148970 667880
rect 149210 667640 149300 667880
rect 149540 667640 149630 667880
rect 149870 667640 149960 667880
rect 150200 667640 150310 667880
rect 150550 667640 150640 667880
rect 150880 667640 150970 667880
rect 151210 667640 151300 667880
rect 151540 667640 151650 667880
rect 151890 667640 151980 667880
rect 152220 667640 152310 667880
rect 152550 667640 152640 667880
rect 152880 667640 152990 667880
rect 153230 667640 153320 667880
rect 153560 667640 153650 667880
rect 153890 667640 153980 667880
rect 154220 667640 154330 667880
rect 154570 667640 154660 667880
rect 154900 667640 154990 667880
rect 155230 667640 155320 667880
rect 155560 667640 155670 667880
rect 155910 667640 155960 667880
rect 110760 667530 155960 667640
rect 110760 667290 110810 667530
rect 111050 667290 111140 667530
rect 111380 667290 111470 667530
rect 111710 667290 111800 667530
rect 112040 667290 112150 667530
rect 112390 667290 112480 667530
rect 112720 667290 112810 667530
rect 113050 667290 113140 667530
rect 113380 667290 113490 667530
rect 113730 667290 113820 667530
rect 114060 667290 114150 667530
rect 114390 667290 114480 667530
rect 114720 667290 114830 667530
rect 115070 667290 115160 667530
rect 115400 667290 115490 667530
rect 115730 667290 115820 667530
rect 116060 667290 116170 667530
rect 116410 667290 116500 667530
rect 116740 667290 116830 667530
rect 117070 667290 117160 667530
rect 117400 667290 117510 667530
rect 117750 667290 117840 667530
rect 118080 667290 118170 667530
rect 118410 667290 118500 667530
rect 118740 667290 118850 667530
rect 119090 667290 119180 667530
rect 119420 667290 119510 667530
rect 119750 667290 119840 667530
rect 120080 667290 120190 667530
rect 120430 667290 120520 667530
rect 120760 667290 120850 667530
rect 121090 667290 121180 667530
rect 121420 667290 121530 667530
rect 121770 667290 122190 667530
rect 122430 667290 122520 667530
rect 122760 667290 122850 667530
rect 123090 667290 123180 667530
rect 123420 667290 123530 667530
rect 123770 667290 123860 667530
rect 124100 667290 124190 667530
rect 124430 667290 124520 667530
rect 124760 667290 124870 667530
rect 125110 667290 125200 667530
rect 125440 667290 125530 667530
rect 125770 667290 125860 667530
rect 126100 667290 126210 667530
rect 126450 667290 126540 667530
rect 126780 667290 126870 667530
rect 127110 667290 127200 667530
rect 127440 667290 127550 667530
rect 127790 667290 127880 667530
rect 128120 667290 128210 667530
rect 128450 667290 128540 667530
rect 128780 667290 128890 667530
rect 129130 667290 129220 667530
rect 129460 667290 129550 667530
rect 129790 667290 129880 667530
rect 130120 667290 130230 667530
rect 130470 667290 130560 667530
rect 130800 667290 130890 667530
rect 131130 667290 131220 667530
rect 131460 667290 131570 667530
rect 131810 667290 131900 667530
rect 132140 667290 132230 667530
rect 132470 667290 132560 667530
rect 132800 667290 132910 667530
rect 133150 667290 133570 667530
rect 133810 667290 133900 667530
rect 134140 667290 134230 667530
rect 134470 667290 134560 667530
rect 134800 667290 134910 667530
rect 135150 667290 135240 667530
rect 135480 667290 135570 667530
rect 135810 667290 135900 667530
rect 136140 667290 136250 667530
rect 136490 667290 136580 667530
rect 136820 667290 136910 667530
rect 137150 667290 137240 667530
rect 137480 667290 137590 667530
rect 137830 667290 137920 667530
rect 138160 667290 138250 667530
rect 138490 667290 138580 667530
rect 138820 667290 138930 667530
rect 139170 667290 139260 667530
rect 139500 667290 139590 667530
rect 139830 667290 139920 667530
rect 140160 667290 140270 667530
rect 140510 667290 140600 667530
rect 140840 667290 140930 667530
rect 141170 667290 141260 667530
rect 141500 667290 141610 667530
rect 141850 667290 141940 667530
rect 142180 667290 142270 667530
rect 142510 667290 142600 667530
rect 142840 667290 142950 667530
rect 143190 667290 143280 667530
rect 143520 667290 143610 667530
rect 143850 667290 143940 667530
rect 144180 667290 144290 667530
rect 144530 667290 144950 667530
rect 145190 667290 145280 667530
rect 145520 667290 145610 667530
rect 145850 667290 145940 667530
rect 146180 667290 146290 667530
rect 146530 667290 146620 667530
rect 146860 667290 146950 667530
rect 147190 667290 147280 667530
rect 147520 667290 147630 667530
rect 147870 667290 147960 667530
rect 148200 667290 148290 667530
rect 148530 667290 148620 667530
rect 148860 667290 148970 667530
rect 149210 667290 149300 667530
rect 149540 667290 149630 667530
rect 149870 667290 149960 667530
rect 150200 667290 150310 667530
rect 150550 667290 150640 667530
rect 150880 667290 150970 667530
rect 151210 667290 151300 667530
rect 151540 667290 151650 667530
rect 151890 667290 151980 667530
rect 152220 667290 152310 667530
rect 152550 667290 152640 667530
rect 152880 667290 152990 667530
rect 153230 667290 153320 667530
rect 153560 667290 153650 667530
rect 153890 667290 153980 667530
rect 154220 667290 154330 667530
rect 154570 667290 154660 667530
rect 154900 667290 154990 667530
rect 155230 667290 155320 667530
rect 155560 667290 155670 667530
rect 155910 667290 155960 667530
rect 110760 667200 155960 667290
rect 110760 666960 110810 667200
rect 111050 666960 111140 667200
rect 111380 666960 111470 667200
rect 111710 666960 111800 667200
rect 112040 666960 112150 667200
rect 112390 666960 112480 667200
rect 112720 666960 112810 667200
rect 113050 666960 113140 667200
rect 113380 666960 113490 667200
rect 113730 666960 113820 667200
rect 114060 666960 114150 667200
rect 114390 666960 114480 667200
rect 114720 666960 114830 667200
rect 115070 666960 115160 667200
rect 115400 666960 115490 667200
rect 115730 666960 115820 667200
rect 116060 666960 116170 667200
rect 116410 666960 116500 667200
rect 116740 666960 116830 667200
rect 117070 666960 117160 667200
rect 117400 666960 117510 667200
rect 117750 666960 117840 667200
rect 118080 666960 118170 667200
rect 118410 666960 118500 667200
rect 118740 666960 118850 667200
rect 119090 666960 119180 667200
rect 119420 666960 119510 667200
rect 119750 666960 119840 667200
rect 120080 666960 120190 667200
rect 120430 666960 120520 667200
rect 120760 666960 120850 667200
rect 121090 666960 121180 667200
rect 121420 666960 121530 667200
rect 121770 666960 122190 667200
rect 122430 666960 122520 667200
rect 122760 666960 122850 667200
rect 123090 666960 123180 667200
rect 123420 666960 123530 667200
rect 123770 666960 123860 667200
rect 124100 666960 124190 667200
rect 124430 666960 124520 667200
rect 124760 666960 124870 667200
rect 125110 666960 125200 667200
rect 125440 666960 125530 667200
rect 125770 666960 125860 667200
rect 126100 666960 126210 667200
rect 126450 666960 126540 667200
rect 126780 666960 126870 667200
rect 127110 666960 127200 667200
rect 127440 666960 127550 667200
rect 127790 666960 127880 667200
rect 128120 666960 128210 667200
rect 128450 666960 128540 667200
rect 128780 666960 128890 667200
rect 129130 666960 129220 667200
rect 129460 666960 129550 667200
rect 129790 666960 129880 667200
rect 130120 666960 130230 667200
rect 130470 666960 130560 667200
rect 130800 666960 130890 667200
rect 131130 666960 131220 667200
rect 131460 666960 131570 667200
rect 131810 666960 131900 667200
rect 132140 666960 132230 667200
rect 132470 666960 132560 667200
rect 132800 666960 132910 667200
rect 133150 666960 133570 667200
rect 133810 666960 133900 667200
rect 134140 666960 134230 667200
rect 134470 666960 134560 667200
rect 134800 666960 134910 667200
rect 135150 666960 135240 667200
rect 135480 666960 135570 667200
rect 135810 666960 135900 667200
rect 136140 666960 136250 667200
rect 136490 666960 136580 667200
rect 136820 666960 136910 667200
rect 137150 666960 137240 667200
rect 137480 666960 137590 667200
rect 137830 666960 137920 667200
rect 138160 666960 138250 667200
rect 138490 666960 138580 667200
rect 138820 666960 138930 667200
rect 139170 666960 139260 667200
rect 139500 666960 139590 667200
rect 139830 666960 139920 667200
rect 140160 666960 140270 667200
rect 140510 666960 140600 667200
rect 140840 666960 140930 667200
rect 141170 666960 141260 667200
rect 141500 666960 141610 667200
rect 141850 666960 141940 667200
rect 142180 666960 142270 667200
rect 142510 666960 142600 667200
rect 142840 666960 142950 667200
rect 143190 666960 143280 667200
rect 143520 666960 143610 667200
rect 143850 666960 143940 667200
rect 144180 666960 144290 667200
rect 144530 666960 144950 667200
rect 145190 666960 145280 667200
rect 145520 666960 145610 667200
rect 145850 666960 145940 667200
rect 146180 666960 146290 667200
rect 146530 666960 146620 667200
rect 146860 666960 146950 667200
rect 147190 666960 147280 667200
rect 147520 666960 147630 667200
rect 147870 666960 147960 667200
rect 148200 666960 148290 667200
rect 148530 666960 148620 667200
rect 148860 666960 148970 667200
rect 149210 666960 149300 667200
rect 149540 666960 149630 667200
rect 149870 666960 149960 667200
rect 150200 666960 150310 667200
rect 150550 666960 150640 667200
rect 150880 666960 150970 667200
rect 151210 666960 151300 667200
rect 151540 666960 151650 667200
rect 151890 666960 151980 667200
rect 152220 666960 152310 667200
rect 152550 666960 152640 667200
rect 152880 666960 152990 667200
rect 153230 666960 153320 667200
rect 153560 666960 153650 667200
rect 153890 666960 153980 667200
rect 154220 666960 154330 667200
rect 154570 666960 154660 667200
rect 154900 666960 154990 667200
rect 155230 666960 155320 667200
rect 155560 666960 155670 667200
rect 155910 666960 155960 667200
rect 110760 666870 155960 666960
rect 110760 666630 110810 666870
rect 111050 666630 111140 666870
rect 111380 666630 111470 666870
rect 111710 666630 111800 666870
rect 112040 666630 112150 666870
rect 112390 666630 112480 666870
rect 112720 666630 112810 666870
rect 113050 666630 113140 666870
rect 113380 666630 113490 666870
rect 113730 666630 113820 666870
rect 114060 666630 114150 666870
rect 114390 666630 114480 666870
rect 114720 666630 114830 666870
rect 115070 666630 115160 666870
rect 115400 666630 115490 666870
rect 115730 666630 115820 666870
rect 116060 666630 116170 666870
rect 116410 666630 116500 666870
rect 116740 666630 116830 666870
rect 117070 666630 117160 666870
rect 117400 666630 117510 666870
rect 117750 666630 117840 666870
rect 118080 666630 118170 666870
rect 118410 666630 118500 666870
rect 118740 666630 118850 666870
rect 119090 666630 119180 666870
rect 119420 666630 119510 666870
rect 119750 666630 119840 666870
rect 120080 666630 120190 666870
rect 120430 666630 120520 666870
rect 120760 666630 120850 666870
rect 121090 666630 121180 666870
rect 121420 666630 121530 666870
rect 121770 666630 122190 666870
rect 122430 666630 122520 666870
rect 122760 666630 122850 666870
rect 123090 666630 123180 666870
rect 123420 666630 123530 666870
rect 123770 666630 123860 666870
rect 124100 666630 124190 666870
rect 124430 666630 124520 666870
rect 124760 666630 124870 666870
rect 125110 666630 125200 666870
rect 125440 666630 125530 666870
rect 125770 666630 125860 666870
rect 126100 666630 126210 666870
rect 126450 666630 126540 666870
rect 126780 666630 126870 666870
rect 127110 666630 127200 666870
rect 127440 666630 127550 666870
rect 127790 666630 127880 666870
rect 128120 666630 128210 666870
rect 128450 666630 128540 666870
rect 128780 666630 128890 666870
rect 129130 666630 129220 666870
rect 129460 666630 129550 666870
rect 129790 666630 129880 666870
rect 130120 666630 130230 666870
rect 130470 666630 130560 666870
rect 130800 666630 130890 666870
rect 131130 666630 131220 666870
rect 131460 666630 131570 666870
rect 131810 666630 131900 666870
rect 132140 666630 132230 666870
rect 132470 666630 132560 666870
rect 132800 666630 132910 666870
rect 133150 666630 133570 666870
rect 133810 666630 133900 666870
rect 134140 666630 134230 666870
rect 134470 666630 134560 666870
rect 134800 666630 134910 666870
rect 135150 666630 135240 666870
rect 135480 666630 135570 666870
rect 135810 666630 135900 666870
rect 136140 666630 136250 666870
rect 136490 666630 136580 666870
rect 136820 666630 136910 666870
rect 137150 666630 137240 666870
rect 137480 666630 137590 666870
rect 137830 666630 137920 666870
rect 138160 666630 138250 666870
rect 138490 666630 138580 666870
rect 138820 666630 138930 666870
rect 139170 666630 139260 666870
rect 139500 666630 139590 666870
rect 139830 666630 139920 666870
rect 140160 666630 140270 666870
rect 140510 666630 140600 666870
rect 140840 666630 140930 666870
rect 141170 666630 141260 666870
rect 141500 666630 141610 666870
rect 141850 666630 141940 666870
rect 142180 666630 142270 666870
rect 142510 666630 142600 666870
rect 142840 666630 142950 666870
rect 143190 666630 143280 666870
rect 143520 666630 143610 666870
rect 143850 666630 143940 666870
rect 144180 666630 144290 666870
rect 144530 666630 144950 666870
rect 145190 666630 145280 666870
rect 145520 666630 145610 666870
rect 145850 666630 145940 666870
rect 146180 666630 146290 666870
rect 146530 666630 146620 666870
rect 146860 666630 146950 666870
rect 147190 666630 147280 666870
rect 147520 666630 147630 666870
rect 147870 666630 147960 666870
rect 148200 666630 148290 666870
rect 148530 666630 148620 666870
rect 148860 666630 148970 666870
rect 149210 666630 149300 666870
rect 149540 666630 149630 666870
rect 149870 666630 149960 666870
rect 150200 666630 150310 666870
rect 150550 666630 150640 666870
rect 150880 666630 150970 666870
rect 151210 666630 151300 666870
rect 151540 666630 151650 666870
rect 151890 666630 151980 666870
rect 152220 666630 152310 666870
rect 152550 666630 152640 666870
rect 152880 666630 152990 666870
rect 153230 666630 153320 666870
rect 153560 666630 153650 666870
rect 153890 666630 153980 666870
rect 154220 666630 154330 666870
rect 154570 666630 154660 666870
rect 154900 666630 154990 666870
rect 155230 666630 155320 666870
rect 155560 666630 155670 666870
rect 155910 666630 155960 666870
rect 110760 666540 155960 666630
rect 110760 666300 110810 666540
rect 111050 666300 111140 666540
rect 111380 666300 111470 666540
rect 111710 666300 111800 666540
rect 112040 666300 112150 666540
rect 112390 666300 112480 666540
rect 112720 666300 112810 666540
rect 113050 666300 113140 666540
rect 113380 666300 113490 666540
rect 113730 666300 113820 666540
rect 114060 666300 114150 666540
rect 114390 666300 114480 666540
rect 114720 666300 114830 666540
rect 115070 666300 115160 666540
rect 115400 666300 115490 666540
rect 115730 666300 115820 666540
rect 116060 666300 116170 666540
rect 116410 666300 116500 666540
rect 116740 666300 116830 666540
rect 117070 666300 117160 666540
rect 117400 666300 117510 666540
rect 117750 666300 117840 666540
rect 118080 666300 118170 666540
rect 118410 666300 118500 666540
rect 118740 666300 118850 666540
rect 119090 666300 119180 666540
rect 119420 666300 119510 666540
rect 119750 666300 119840 666540
rect 120080 666300 120190 666540
rect 120430 666300 120520 666540
rect 120760 666300 120850 666540
rect 121090 666300 121180 666540
rect 121420 666300 121530 666540
rect 121770 666300 122190 666540
rect 122430 666300 122520 666540
rect 122760 666300 122850 666540
rect 123090 666300 123180 666540
rect 123420 666300 123530 666540
rect 123770 666300 123860 666540
rect 124100 666300 124190 666540
rect 124430 666300 124520 666540
rect 124760 666300 124870 666540
rect 125110 666300 125200 666540
rect 125440 666300 125530 666540
rect 125770 666300 125860 666540
rect 126100 666300 126210 666540
rect 126450 666300 126540 666540
rect 126780 666300 126870 666540
rect 127110 666300 127200 666540
rect 127440 666300 127550 666540
rect 127790 666300 127880 666540
rect 128120 666300 128210 666540
rect 128450 666300 128540 666540
rect 128780 666300 128890 666540
rect 129130 666300 129220 666540
rect 129460 666300 129550 666540
rect 129790 666300 129880 666540
rect 130120 666300 130230 666540
rect 130470 666300 130560 666540
rect 130800 666300 130890 666540
rect 131130 666300 131220 666540
rect 131460 666300 131570 666540
rect 131810 666300 131900 666540
rect 132140 666300 132230 666540
rect 132470 666300 132560 666540
rect 132800 666300 132910 666540
rect 133150 666300 133570 666540
rect 133810 666300 133900 666540
rect 134140 666300 134230 666540
rect 134470 666300 134560 666540
rect 134800 666300 134910 666540
rect 135150 666300 135240 666540
rect 135480 666300 135570 666540
rect 135810 666300 135900 666540
rect 136140 666300 136250 666540
rect 136490 666300 136580 666540
rect 136820 666300 136910 666540
rect 137150 666300 137240 666540
rect 137480 666300 137590 666540
rect 137830 666300 137920 666540
rect 138160 666300 138250 666540
rect 138490 666300 138580 666540
rect 138820 666300 138930 666540
rect 139170 666300 139260 666540
rect 139500 666300 139590 666540
rect 139830 666300 139920 666540
rect 140160 666300 140270 666540
rect 140510 666300 140600 666540
rect 140840 666300 140930 666540
rect 141170 666300 141260 666540
rect 141500 666300 141610 666540
rect 141850 666300 141940 666540
rect 142180 666300 142270 666540
rect 142510 666300 142600 666540
rect 142840 666300 142950 666540
rect 143190 666300 143280 666540
rect 143520 666300 143610 666540
rect 143850 666300 143940 666540
rect 144180 666300 144290 666540
rect 144530 666300 144950 666540
rect 145190 666300 145280 666540
rect 145520 666300 145610 666540
rect 145850 666300 145940 666540
rect 146180 666300 146290 666540
rect 146530 666300 146620 666540
rect 146860 666300 146950 666540
rect 147190 666300 147280 666540
rect 147520 666300 147630 666540
rect 147870 666300 147960 666540
rect 148200 666300 148290 666540
rect 148530 666300 148620 666540
rect 148860 666300 148970 666540
rect 149210 666300 149300 666540
rect 149540 666300 149630 666540
rect 149870 666300 149960 666540
rect 150200 666300 150310 666540
rect 150550 666300 150640 666540
rect 150880 666300 150970 666540
rect 151210 666300 151300 666540
rect 151540 666300 151650 666540
rect 151890 666300 151980 666540
rect 152220 666300 152310 666540
rect 152550 666300 152640 666540
rect 152880 666300 152990 666540
rect 153230 666300 153320 666540
rect 153560 666300 153650 666540
rect 153890 666300 153980 666540
rect 154220 666300 154330 666540
rect 154570 666300 154660 666540
rect 154900 666300 154990 666540
rect 155230 666300 155320 666540
rect 155560 666300 155670 666540
rect 155910 666300 155960 666540
rect 110760 666190 155960 666300
rect 110760 665950 110810 666190
rect 111050 665950 111140 666190
rect 111380 665950 111470 666190
rect 111710 665950 111800 666190
rect 112040 665950 112150 666190
rect 112390 665950 112480 666190
rect 112720 665950 112810 666190
rect 113050 665950 113140 666190
rect 113380 665950 113490 666190
rect 113730 665950 113820 666190
rect 114060 665950 114150 666190
rect 114390 665950 114480 666190
rect 114720 665950 114830 666190
rect 115070 665950 115160 666190
rect 115400 665950 115490 666190
rect 115730 665950 115820 666190
rect 116060 665950 116170 666190
rect 116410 665950 116500 666190
rect 116740 665950 116830 666190
rect 117070 665950 117160 666190
rect 117400 665950 117510 666190
rect 117750 665950 117840 666190
rect 118080 665950 118170 666190
rect 118410 665950 118500 666190
rect 118740 665950 118850 666190
rect 119090 665950 119180 666190
rect 119420 665950 119510 666190
rect 119750 665950 119840 666190
rect 120080 665950 120190 666190
rect 120430 665950 120520 666190
rect 120760 665950 120850 666190
rect 121090 665950 121180 666190
rect 121420 665950 121530 666190
rect 121770 665950 122190 666190
rect 122430 665950 122520 666190
rect 122760 665950 122850 666190
rect 123090 665950 123180 666190
rect 123420 665950 123530 666190
rect 123770 665950 123860 666190
rect 124100 665950 124190 666190
rect 124430 665950 124520 666190
rect 124760 665950 124870 666190
rect 125110 665950 125200 666190
rect 125440 665950 125530 666190
rect 125770 665950 125860 666190
rect 126100 665950 126210 666190
rect 126450 665950 126540 666190
rect 126780 665950 126870 666190
rect 127110 665950 127200 666190
rect 127440 665950 127550 666190
rect 127790 665950 127880 666190
rect 128120 665950 128210 666190
rect 128450 665950 128540 666190
rect 128780 665950 128890 666190
rect 129130 665950 129220 666190
rect 129460 665950 129550 666190
rect 129790 665950 129880 666190
rect 130120 665950 130230 666190
rect 130470 665950 130560 666190
rect 130800 665950 130890 666190
rect 131130 665950 131220 666190
rect 131460 665950 131570 666190
rect 131810 665950 131900 666190
rect 132140 665950 132230 666190
rect 132470 665950 132560 666190
rect 132800 665950 132910 666190
rect 133150 665950 133570 666190
rect 133810 665950 133900 666190
rect 134140 665950 134230 666190
rect 134470 665950 134560 666190
rect 134800 665950 134910 666190
rect 135150 665950 135240 666190
rect 135480 665950 135570 666190
rect 135810 665950 135900 666190
rect 136140 665950 136250 666190
rect 136490 665950 136580 666190
rect 136820 665950 136910 666190
rect 137150 665950 137240 666190
rect 137480 665950 137590 666190
rect 137830 665950 137920 666190
rect 138160 665950 138250 666190
rect 138490 665950 138580 666190
rect 138820 665950 138930 666190
rect 139170 665950 139260 666190
rect 139500 665950 139590 666190
rect 139830 665950 139920 666190
rect 140160 665950 140270 666190
rect 140510 665950 140600 666190
rect 140840 665950 140930 666190
rect 141170 665950 141260 666190
rect 141500 665950 141610 666190
rect 141850 665950 141940 666190
rect 142180 665950 142270 666190
rect 142510 665950 142600 666190
rect 142840 665950 142950 666190
rect 143190 665950 143280 666190
rect 143520 665950 143610 666190
rect 143850 665950 143940 666190
rect 144180 665950 144290 666190
rect 144530 665950 144950 666190
rect 145190 665950 145280 666190
rect 145520 665950 145610 666190
rect 145850 665950 145940 666190
rect 146180 665950 146290 666190
rect 146530 665950 146620 666190
rect 146860 665950 146950 666190
rect 147190 665950 147280 666190
rect 147520 665950 147630 666190
rect 147870 665950 147960 666190
rect 148200 665950 148290 666190
rect 148530 665950 148620 666190
rect 148860 665950 148970 666190
rect 149210 665950 149300 666190
rect 149540 665950 149630 666190
rect 149870 665950 149960 666190
rect 150200 665950 150310 666190
rect 150550 665950 150640 666190
rect 150880 665950 150970 666190
rect 151210 665950 151300 666190
rect 151540 665950 151650 666190
rect 151890 665950 151980 666190
rect 152220 665950 152310 666190
rect 152550 665950 152640 666190
rect 152880 665950 152990 666190
rect 153230 665950 153320 666190
rect 153560 665950 153650 666190
rect 153890 665950 153980 666190
rect 154220 665950 154330 666190
rect 154570 665950 154660 666190
rect 154900 665950 154990 666190
rect 155230 665950 155320 666190
rect 155560 665950 155670 666190
rect 155910 665950 155960 666190
rect 110760 665860 155960 665950
rect 110760 665620 110810 665860
rect 111050 665620 111140 665860
rect 111380 665620 111470 665860
rect 111710 665620 111800 665860
rect 112040 665620 112150 665860
rect 112390 665620 112480 665860
rect 112720 665620 112810 665860
rect 113050 665620 113140 665860
rect 113380 665620 113490 665860
rect 113730 665620 113820 665860
rect 114060 665620 114150 665860
rect 114390 665620 114480 665860
rect 114720 665620 114830 665860
rect 115070 665620 115160 665860
rect 115400 665620 115490 665860
rect 115730 665620 115820 665860
rect 116060 665620 116170 665860
rect 116410 665620 116500 665860
rect 116740 665620 116830 665860
rect 117070 665620 117160 665860
rect 117400 665620 117510 665860
rect 117750 665620 117840 665860
rect 118080 665620 118170 665860
rect 118410 665620 118500 665860
rect 118740 665620 118850 665860
rect 119090 665620 119180 665860
rect 119420 665620 119510 665860
rect 119750 665620 119840 665860
rect 120080 665620 120190 665860
rect 120430 665620 120520 665860
rect 120760 665620 120850 665860
rect 121090 665620 121180 665860
rect 121420 665620 121530 665860
rect 121770 665620 122190 665860
rect 122430 665620 122520 665860
rect 122760 665620 122850 665860
rect 123090 665620 123180 665860
rect 123420 665620 123530 665860
rect 123770 665620 123860 665860
rect 124100 665620 124190 665860
rect 124430 665620 124520 665860
rect 124760 665620 124870 665860
rect 125110 665620 125200 665860
rect 125440 665620 125530 665860
rect 125770 665620 125860 665860
rect 126100 665620 126210 665860
rect 126450 665620 126540 665860
rect 126780 665620 126870 665860
rect 127110 665620 127200 665860
rect 127440 665620 127550 665860
rect 127790 665620 127880 665860
rect 128120 665620 128210 665860
rect 128450 665620 128540 665860
rect 128780 665620 128890 665860
rect 129130 665620 129220 665860
rect 129460 665620 129550 665860
rect 129790 665620 129880 665860
rect 130120 665620 130230 665860
rect 130470 665620 130560 665860
rect 130800 665620 130890 665860
rect 131130 665620 131220 665860
rect 131460 665620 131570 665860
rect 131810 665620 131900 665860
rect 132140 665620 132230 665860
rect 132470 665620 132560 665860
rect 132800 665620 132910 665860
rect 133150 665620 133570 665860
rect 133810 665620 133900 665860
rect 134140 665620 134230 665860
rect 134470 665620 134560 665860
rect 134800 665620 134910 665860
rect 135150 665620 135240 665860
rect 135480 665620 135570 665860
rect 135810 665620 135900 665860
rect 136140 665620 136250 665860
rect 136490 665620 136580 665860
rect 136820 665620 136910 665860
rect 137150 665620 137240 665860
rect 137480 665620 137590 665860
rect 137830 665620 137920 665860
rect 138160 665620 138250 665860
rect 138490 665620 138580 665860
rect 138820 665620 138930 665860
rect 139170 665620 139260 665860
rect 139500 665620 139590 665860
rect 139830 665620 139920 665860
rect 140160 665620 140270 665860
rect 140510 665620 140600 665860
rect 140840 665620 140930 665860
rect 141170 665620 141260 665860
rect 141500 665620 141610 665860
rect 141850 665620 141940 665860
rect 142180 665620 142270 665860
rect 142510 665620 142600 665860
rect 142840 665620 142950 665860
rect 143190 665620 143280 665860
rect 143520 665620 143610 665860
rect 143850 665620 143940 665860
rect 144180 665620 144290 665860
rect 144530 665620 144950 665860
rect 145190 665620 145280 665860
rect 145520 665620 145610 665860
rect 145850 665620 145940 665860
rect 146180 665620 146290 665860
rect 146530 665620 146620 665860
rect 146860 665620 146950 665860
rect 147190 665620 147280 665860
rect 147520 665620 147630 665860
rect 147870 665620 147960 665860
rect 148200 665620 148290 665860
rect 148530 665620 148620 665860
rect 148860 665620 148970 665860
rect 149210 665620 149300 665860
rect 149540 665620 149630 665860
rect 149870 665620 149960 665860
rect 150200 665620 150310 665860
rect 150550 665620 150640 665860
rect 150880 665620 150970 665860
rect 151210 665620 151300 665860
rect 151540 665620 151650 665860
rect 151890 665620 151980 665860
rect 152220 665620 152310 665860
rect 152550 665620 152640 665860
rect 152880 665620 152990 665860
rect 153230 665620 153320 665860
rect 153560 665620 153650 665860
rect 153890 665620 153980 665860
rect 154220 665620 154330 665860
rect 154570 665620 154660 665860
rect 154900 665620 154990 665860
rect 155230 665620 155320 665860
rect 155560 665620 155670 665860
rect 155910 665620 155960 665860
rect 110760 665530 155960 665620
rect 110760 665290 110810 665530
rect 111050 665290 111140 665530
rect 111380 665290 111470 665530
rect 111710 665290 111800 665530
rect 112040 665290 112150 665530
rect 112390 665290 112480 665530
rect 112720 665290 112810 665530
rect 113050 665290 113140 665530
rect 113380 665290 113490 665530
rect 113730 665290 113820 665530
rect 114060 665290 114150 665530
rect 114390 665290 114480 665530
rect 114720 665290 114830 665530
rect 115070 665290 115160 665530
rect 115400 665290 115490 665530
rect 115730 665290 115820 665530
rect 116060 665290 116170 665530
rect 116410 665290 116500 665530
rect 116740 665290 116830 665530
rect 117070 665290 117160 665530
rect 117400 665290 117510 665530
rect 117750 665290 117840 665530
rect 118080 665290 118170 665530
rect 118410 665290 118500 665530
rect 118740 665290 118850 665530
rect 119090 665290 119180 665530
rect 119420 665290 119510 665530
rect 119750 665290 119840 665530
rect 120080 665290 120190 665530
rect 120430 665290 120520 665530
rect 120760 665290 120850 665530
rect 121090 665290 121180 665530
rect 121420 665290 121530 665530
rect 121770 665290 122190 665530
rect 122430 665290 122520 665530
rect 122760 665290 122850 665530
rect 123090 665290 123180 665530
rect 123420 665290 123530 665530
rect 123770 665290 123860 665530
rect 124100 665290 124190 665530
rect 124430 665290 124520 665530
rect 124760 665290 124870 665530
rect 125110 665290 125200 665530
rect 125440 665290 125530 665530
rect 125770 665290 125860 665530
rect 126100 665290 126210 665530
rect 126450 665290 126540 665530
rect 126780 665290 126870 665530
rect 127110 665290 127200 665530
rect 127440 665290 127550 665530
rect 127790 665290 127880 665530
rect 128120 665290 128210 665530
rect 128450 665290 128540 665530
rect 128780 665290 128890 665530
rect 129130 665290 129220 665530
rect 129460 665290 129550 665530
rect 129790 665290 129880 665530
rect 130120 665290 130230 665530
rect 130470 665290 130560 665530
rect 130800 665290 130890 665530
rect 131130 665290 131220 665530
rect 131460 665290 131570 665530
rect 131810 665290 131900 665530
rect 132140 665290 132230 665530
rect 132470 665290 132560 665530
rect 132800 665290 132910 665530
rect 133150 665290 133570 665530
rect 133810 665290 133900 665530
rect 134140 665290 134230 665530
rect 134470 665290 134560 665530
rect 134800 665290 134910 665530
rect 135150 665290 135240 665530
rect 135480 665290 135570 665530
rect 135810 665290 135900 665530
rect 136140 665290 136250 665530
rect 136490 665290 136580 665530
rect 136820 665290 136910 665530
rect 137150 665290 137240 665530
rect 137480 665290 137590 665530
rect 137830 665290 137920 665530
rect 138160 665290 138250 665530
rect 138490 665290 138580 665530
rect 138820 665290 138930 665530
rect 139170 665290 139260 665530
rect 139500 665290 139590 665530
rect 139830 665290 139920 665530
rect 140160 665290 140270 665530
rect 140510 665290 140600 665530
rect 140840 665290 140930 665530
rect 141170 665290 141260 665530
rect 141500 665290 141610 665530
rect 141850 665290 141940 665530
rect 142180 665290 142270 665530
rect 142510 665290 142600 665530
rect 142840 665290 142950 665530
rect 143190 665290 143280 665530
rect 143520 665290 143610 665530
rect 143850 665290 143940 665530
rect 144180 665290 144290 665530
rect 144530 665290 144950 665530
rect 145190 665290 145280 665530
rect 145520 665290 145610 665530
rect 145850 665290 145940 665530
rect 146180 665290 146290 665530
rect 146530 665290 146620 665530
rect 146860 665290 146950 665530
rect 147190 665290 147280 665530
rect 147520 665290 147630 665530
rect 147870 665290 147960 665530
rect 148200 665290 148290 665530
rect 148530 665290 148620 665530
rect 148860 665290 148970 665530
rect 149210 665290 149300 665530
rect 149540 665290 149630 665530
rect 149870 665290 149960 665530
rect 150200 665290 150310 665530
rect 150550 665290 150640 665530
rect 150880 665290 150970 665530
rect 151210 665290 151300 665530
rect 151540 665290 151650 665530
rect 151890 665290 151980 665530
rect 152220 665290 152310 665530
rect 152550 665290 152640 665530
rect 152880 665290 152990 665530
rect 153230 665290 153320 665530
rect 153560 665290 153650 665530
rect 153890 665290 153980 665530
rect 154220 665290 154330 665530
rect 154570 665290 154660 665530
rect 154900 665290 154990 665530
rect 155230 665290 155320 665530
rect 155560 665290 155670 665530
rect 155910 665290 155960 665530
rect 110760 665200 155960 665290
rect 110760 664960 110810 665200
rect 111050 664960 111140 665200
rect 111380 664960 111470 665200
rect 111710 664960 111800 665200
rect 112040 664960 112150 665200
rect 112390 664960 112480 665200
rect 112720 664960 112810 665200
rect 113050 664960 113140 665200
rect 113380 664960 113490 665200
rect 113730 664960 113820 665200
rect 114060 664960 114150 665200
rect 114390 664960 114480 665200
rect 114720 664960 114830 665200
rect 115070 664960 115160 665200
rect 115400 664960 115490 665200
rect 115730 664960 115820 665200
rect 116060 664960 116170 665200
rect 116410 664960 116500 665200
rect 116740 664960 116830 665200
rect 117070 664960 117160 665200
rect 117400 664960 117510 665200
rect 117750 664960 117840 665200
rect 118080 664960 118170 665200
rect 118410 664960 118500 665200
rect 118740 664960 118850 665200
rect 119090 664960 119180 665200
rect 119420 664960 119510 665200
rect 119750 664960 119840 665200
rect 120080 664960 120190 665200
rect 120430 664960 120520 665200
rect 120760 664960 120850 665200
rect 121090 664960 121180 665200
rect 121420 664960 121530 665200
rect 121770 664960 122190 665200
rect 122430 664960 122520 665200
rect 122760 664960 122850 665200
rect 123090 664960 123180 665200
rect 123420 664960 123530 665200
rect 123770 664960 123860 665200
rect 124100 664960 124190 665200
rect 124430 664960 124520 665200
rect 124760 664960 124870 665200
rect 125110 664960 125200 665200
rect 125440 664960 125530 665200
rect 125770 664960 125860 665200
rect 126100 664960 126210 665200
rect 126450 664960 126540 665200
rect 126780 664960 126870 665200
rect 127110 664960 127200 665200
rect 127440 664960 127550 665200
rect 127790 664960 127880 665200
rect 128120 664960 128210 665200
rect 128450 664960 128540 665200
rect 128780 664960 128890 665200
rect 129130 664960 129220 665200
rect 129460 664960 129550 665200
rect 129790 664960 129880 665200
rect 130120 664960 130230 665200
rect 130470 664960 130560 665200
rect 130800 664960 130890 665200
rect 131130 664960 131220 665200
rect 131460 664960 131570 665200
rect 131810 664960 131900 665200
rect 132140 664960 132230 665200
rect 132470 664960 132560 665200
rect 132800 664960 132910 665200
rect 133150 664960 133570 665200
rect 133810 664960 133900 665200
rect 134140 664960 134230 665200
rect 134470 664960 134560 665200
rect 134800 664960 134910 665200
rect 135150 664960 135240 665200
rect 135480 664960 135570 665200
rect 135810 664960 135900 665200
rect 136140 664960 136250 665200
rect 136490 664960 136580 665200
rect 136820 664960 136910 665200
rect 137150 664960 137240 665200
rect 137480 664960 137590 665200
rect 137830 664960 137920 665200
rect 138160 664960 138250 665200
rect 138490 664960 138580 665200
rect 138820 664960 138930 665200
rect 139170 664960 139260 665200
rect 139500 664960 139590 665200
rect 139830 664960 139920 665200
rect 140160 664960 140270 665200
rect 140510 664960 140600 665200
rect 140840 664960 140930 665200
rect 141170 664960 141260 665200
rect 141500 664960 141610 665200
rect 141850 664960 141940 665200
rect 142180 664960 142270 665200
rect 142510 664960 142600 665200
rect 142840 664960 142950 665200
rect 143190 664960 143280 665200
rect 143520 664960 143610 665200
rect 143850 664960 143940 665200
rect 144180 664960 144290 665200
rect 144530 664960 144950 665200
rect 145190 664960 145280 665200
rect 145520 664960 145610 665200
rect 145850 664960 145940 665200
rect 146180 664960 146290 665200
rect 146530 664960 146620 665200
rect 146860 664960 146950 665200
rect 147190 664960 147280 665200
rect 147520 664960 147630 665200
rect 147870 664960 147960 665200
rect 148200 664960 148290 665200
rect 148530 664960 148620 665200
rect 148860 664960 148970 665200
rect 149210 664960 149300 665200
rect 149540 664960 149630 665200
rect 149870 664960 149960 665200
rect 150200 664960 150310 665200
rect 150550 664960 150640 665200
rect 150880 664960 150970 665200
rect 151210 664960 151300 665200
rect 151540 664960 151650 665200
rect 151890 664960 151980 665200
rect 152220 664960 152310 665200
rect 152550 664960 152640 665200
rect 152880 664960 152990 665200
rect 153230 664960 153320 665200
rect 153560 664960 153650 665200
rect 153890 664960 153980 665200
rect 154220 664960 154330 665200
rect 154570 664960 154660 665200
rect 154900 664960 154990 665200
rect 155230 664960 155320 665200
rect 155560 664960 155670 665200
rect 155910 664960 155960 665200
rect 110760 664850 155960 664960
rect 110760 664610 110810 664850
rect 111050 664610 111140 664850
rect 111380 664610 111470 664850
rect 111710 664610 111800 664850
rect 112040 664610 112150 664850
rect 112390 664610 112480 664850
rect 112720 664610 112810 664850
rect 113050 664610 113140 664850
rect 113380 664610 113490 664850
rect 113730 664610 113820 664850
rect 114060 664610 114150 664850
rect 114390 664610 114480 664850
rect 114720 664610 114830 664850
rect 115070 664610 115160 664850
rect 115400 664610 115490 664850
rect 115730 664610 115820 664850
rect 116060 664610 116170 664850
rect 116410 664610 116500 664850
rect 116740 664610 116830 664850
rect 117070 664610 117160 664850
rect 117400 664610 117510 664850
rect 117750 664610 117840 664850
rect 118080 664610 118170 664850
rect 118410 664610 118500 664850
rect 118740 664610 118850 664850
rect 119090 664610 119180 664850
rect 119420 664610 119510 664850
rect 119750 664610 119840 664850
rect 120080 664610 120190 664850
rect 120430 664610 120520 664850
rect 120760 664610 120850 664850
rect 121090 664610 121180 664850
rect 121420 664610 121530 664850
rect 121770 664610 122190 664850
rect 122430 664610 122520 664850
rect 122760 664610 122850 664850
rect 123090 664610 123180 664850
rect 123420 664610 123530 664850
rect 123770 664610 123860 664850
rect 124100 664610 124190 664850
rect 124430 664610 124520 664850
rect 124760 664610 124870 664850
rect 125110 664610 125200 664850
rect 125440 664610 125530 664850
rect 125770 664610 125860 664850
rect 126100 664610 126210 664850
rect 126450 664610 126540 664850
rect 126780 664610 126870 664850
rect 127110 664610 127200 664850
rect 127440 664610 127550 664850
rect 127790 664610 127880 664850
rect 128120 664610 128210 664850
rect 128450 664610 128540 664850
rect 128780 664610 128890 664850
rect 129130 664610 129220 664850
rect 129460 664610 129550 664850
rect 129790 664610 129880 664850
rect 130120 664610 130230 664850
rect 130470 664610 130560 664850
rect 130800 664610 130890 664850
rect 131130 664610 131220 664850
rect 131460 664610 131570 664850
rect 131810 664610 131900 664850
rect 132140 664610 132230 664850
rect 132470 664610 132560 664850
rect 132800 664610 132910 664850
rect 133150 664610 133570 664850
rect 133810 664610 133900 664850
rect 134140 664610 134230 664850
rect 134470 664610 134560 664850
rect 134800 664610 134910 664850
rect 135150 664610 135240 664850
rect 135480 664610 135570 664850
rect 135810 664610 135900 664850
rect 136140 664610 136250 664850
rect 136490 664610 136580 664850
rect 136820 664610 136910 664850
rect 137150 664610 137240 664850
rect 137480 664610 137590 664850
rect 137830 664610 137920 664850
rect 138160 664610 138250 664850
rect 138490 664610 138580 664850
rect 138820 664610 138930 664850
rect 139170 664610 139260 664850
rect 139500 664610 139590 664850
rect 139830 664610 139920 664850
rect 140160 664610 140270 664850
rect 140510 664610 140600 664850
rect 140840 664610 140930 664850
rect 141170 664610 141260 664850
rect 141500 664610 141610 664850
rect 141850 664610 141940 664850
rect 142180 664610 142270 664850
rect 142510 664610 142600 664850
rect 142840 664610 142950 664850
rect 143190 664610 143280 664850
rect 143520 664610 143610 664850
rect 143850 664610 143940 664850
rect 144180 664610 144290 664850
rect 144530 664610 144950 664850
rect 145190 664610 145280 664850
rect 145520 664610 145610 664850
rect 145850 664610 145940 664850
rect 146180 664610 146290 664850
rect 146530 664610 146620 664850
rect 146860 664610 146950 664850
rect 147190 664610 147280 664850
rect 147520 664610 147630 664850
rect 147870 664610 147960 664850
rect 148200 664610 148290 664850
rect 148530 664610 148620 664850
rect 148860 664610 148970 664850
rect 149210 664610 149300 664850
rect 149540 664610 149630 664850
rect 149870 664610 149960 664850
rect 150200 664610 150310 664850
rect 150550 664610 150640 664850
rect 150880 664610 150970 664850
rect 151210 664610 151300 664850
rect 151540 664610 151650 664850
rect 151890 664610 151980 664850
rect 152220 664610 152310 664850
rect 152550 664610 152640 664850
rect 152880 664610 152990 664850
rect 153230 664610 153320 664850
rect 153560 664610 153650 664850
rect 153890 664610 153980 664850
rect 154220 664610 154330 664850
rect 154570 664610 154660 664850
rect 154900 664610 154990 664850
rect 155230 664610 155320 664850
rect 155560 664610 155670 664850
rect 155910 664610 155960 664850
rect 110760 664520 155960 664610
rect 110760 664280 110810 664520
rect 111050 664280 111140 664520
rect 111380 664280 111470 664520
rect 111710 664280 111800 664520
rect 112040 664280 112150 664520
rect 112390 664280 112480 664520
rect 112720 664280 112810 664520
rect 113050 664280 113140 664520
rect 113380 664280 113490 664520
rect 113730 664280 113820 664520
rect 114060 664280 114150 664520
rect 114390 664280 114480 664520
rect 114720 664280 114830 664520
rect 115070 664280 115160 664520
rect 115400 664280 115490 664520
rect 115730 664280 115820 664520
rect 116060 664280 116170 664520
rect 116410 664280 116500 664520
rect 116740 664280 116830 664520
rect 117070 664280 117160 664520
rect 117400 664280 117510 664520
rect 117750 664280 117840 664520
rect 118080 664280 118170 664520
rect 118410 664280 118500 664520
rect 118740 664280 118850 664520
rect 119090 664280 119180 664520
rect 119420 664280 119510 664520
rect 119750 664280 119840 664520
rect 120080 664280 120190 664520
rect 120430 664280 120520 664520
rect 120760 664280 120850 664520
rect 121090 664280 121180 664520
rect 121420 664280 121530 664520
rect 121770 664280 122190 664520
rect 122430 664280 122520 664520
rect 122760 664280 122850 664520
rect 123090 664280 123180 664520
rect 123420 664280 123530 664520
rect 123770 664280 123860 664520
rect 124100 664280 124190 664520
rect 124430 664280 124520 664520
rect 124760 664280 124870 664520
rect 125110 664280 125200 664520
rect 125440 664280 125530 664520
rect 125770 664280 125860 664520
rect 126100 664280 126210 664520
rect 126450 664280 126540 664520
rect 126780 664280 126870 664520
rect 127110 664280 127200 664520
rect 127440 664280 127550 664520
rect 127790 664280 127880 664520
rect 128120 664280 128210 664520
rect 128450 664280 128540 664520
rect 128780 664280 128890 664520
rect 129130 664280 129220 664520
rect 129460 664280 129550 664520
rect 129790 664280 129880 664520
rect 130120 664280 130230 664520
rect 130470 664280 130560 664520
rect 130800 664280 130890 664520
rect 131130 664280 131220 664520
rect 131460 664280 131570 664520
rect 131810 664280 131900 664520
rect 132140 664280 132230 664520
rect 132470 664280 132560 664520
rect 132800 664280 132910 664520
rect 133150 664280 133570 664520
rect 133810 664280 133900 664520
rect 134140 664280 134230 664520
rect 134470 664280 134560 664520
rect 134800 664280 134910 664520
rect 135150 664280 135240 664520
rect 135480 664280 135570 664520
rect 135810 664280 135900 664520
rect 136140 664280 136250 664520
rect 136490 664280 136580 664520
rect 136820 664280 136910 664520
rect 137150 664280 137240 664520
rect 137480 664280 137590 664520
rect 137830 664280 137920 664520
rect 138160 664280 138250 664520
rect 138490 664280 138580 664520
rect 138820 664280 138930 664520
rect 139170 664280 139260 664520
rect 139500 664280 139590 664520
rect 139830 664280 139920 664520
rect 140160 664280 140270 664520
rect 140510 664280 140600 664520
rect 140840 664280 140930 664520
rect 141170 664280 141260 664520
rect 141500 664280 141610 664520
rect 141850 664280 141940 664520
rect 142180 664280 142270 664520
rect 142510 664280 142600 664520
rect 142840 664280 142950 664520
rect 143190 664280 143280 664520
rect 143520 664280 143610 664520
rect 143850 664280 143940 664520
rect 144180 664280 144290 664520
rect 144530 664280 144950 664520
rect 145190 664280 145280 664520
rect 145520 664280 145610 664520
rect 145850 664280 145940 664520
rect 146180 664280 146290 664520
rect 146530 664280 146620 664520
rect 146860 664280 146950 664520
rect 147190 664280 147280 664520
rect 147520 664280 147630 664520
rect 147870 664280 147960 664520
rect 148200 664280 148290 664520
rect 148530 664280 148620 664520
rect 148860 664280 148970 664520
rect 149210 664280 149300 664520
rect 149540 664280 149630 664520
rect 149870 664280 149960 664520
rect 150200 664280 150310 664520
rect 150550 664280 150640 664520
rect 150880 664280 150970 664520
rect 151210 664280 151300 664520
rect 151540 664280 151650 664520
rect 151890 664280 151980 664520
rect 152220 664280 152310 664520
rect 152550 664280 152640 664520
rect 152880 664280 152990 664520
rect 153230 664280 153320 664520
rect 153560 664280 153650 664520
rect 153890 664280 153980 664520
rect 154220 664280 154330 664520
rect 154570 664280 154660 664520
rect 154900 664280 154990 664520
rect 155230 664280 155320 664520
rect 155560 664280 155670 664520
rect 155910 664280 155960 664520
rect 110760 664190 155960 664280
rect 110760 663950 110810 664190
rect 111050 663950 111140 664190
rect 111380 663950 111470 664190
rect 111710 663950 111800 664190
rect 112040 663950 112150 664190
rect 112390 663950 112480 664190
rect 112720 663950 112810 664190
rect 113050 663950 113140 664190
rect 113380 663950 113490 664190
rect 113730 663950 113820 664190
rect 114060 663950 114150 664190
rect 114390 663950 114480 664190
rect 114720 663950 114830 664190
rect 115070 663950 115160 664190
rect 115400 663950 115490 664190
rect 115730 663950 115820 664190
rect 116060 663950 116170 664190
rect 116410 663950 116500 664190
rect 116740 663950 116830 664190
rect 117070 663950 117160 664190
rect 117400 663950 117510 664190
rect 117750 663950 117840 664190
rect 118080 663950 118170 664190
rect 118410 663950 118500 664190
rect 118740 663950 118850 664190
rect 119090 663950 119180 664190
rect 119420 663950 119510 664190
rect 119750 663950 119840 664190
rect 120080 663950 120190 664190
rect 120430 663950 120520 664190
rect 120760 663950 120850 664190
rect 121090 663950 121180 664190
rect 121420 663950 121530 664190
rect 121770 663950 122190 664190
rect 122430 663950 122520 664190
rect 122760 663950 122850 664190
rect 123090 663950 123180 664190
rect 123420 663950 123530 664190
rect 123770 663950 123860 664190
rect 124100 663950 124190 664190
rect 124430 663950 124520 664190
rect 124760 663950 124870 664190
rect 125110 663950 125200 664190
rect 125440 663950 125530 664190
rect 125770 663950 125860 664190
rect 126100 663950 126210 664190
rect 126450 663950 126540 664190
rect 126780 663950 126870 664190
rect 127110 663950 127200 664190
rect 127440 663950 127550 664190
rect 127790 663950 127880 664190
rect 128120 663950 128210 664190
rect 128450 663950 128540 664190
rect 128780 663950 128890 664190
rect 129130 663950 129220 664190
rect 129460 663950 129550 664190
rect 129790 663950 129880 664190
rect 130120 663950 130230 664190
rect 130470 663950 130560 664190
rect 130800 663950 130890 664190
rect 131130 663950 131220 664190
rect 131460 663950 131570 664190
rect 131810 663950 131900 664190
rect 132140 663950 132230 664190
rect 132470 663950 132560 664190
rect 132800 663950 132910 664190
rect 133150 663950 133570 664190
rect 133810 663950 133900 664190
rect 134140 663950 134230 664190
rect 134470 663950 134560 664190
rect 134800 663950 134910 664190
rect 135150 663950 135240 664190
rect 135480 663950 135570 664190
rect 135810 663950 135900 664190
rect 136140 663950 136250 664190
rect 136490 663950 136580 664190
rect 136820 663950 136910 664190
rect 137150 663950 137240 664190
rect 137480 663950 137590 664190
rect 137830 663950 137920 664190
rect 138160 663950 138250 664190
rect 138490 663950 138580 664190
rect 138820 663950 138930 664190
rect 139170 663950 139260 664190
rect 139500 663950 139590 664190
rect 139830 663950 139920 664190
rect 140160 663950 140270 664190
rect 140510 663950 140600 664190
rect 140840 663950 140930 664190
rect 141170 663950 141260 664190
rect 141500 663950 141610 664190
rect 141850 663950 141940 664190
rect 142180 663950 142270 664190
rect 142510 663950 142600 664190
rect 142840 663950 142950 664190
rect 143190 663950 143280 664190
rect 143520 663950 143610 664190
rect 143850 663950 143940 664190
rect 144180 663950 144290 664190
rect 144530 663950 144950 664190
rect 145190 663950 145280 664190
rect 145520 663950 145610 664190
rect 145850 663950 145940 664190
rect 146180 663950 146290 664190
rect 146530 663950 146620 664190
rect 146860 663950 146950 664190
rect 147190 663950 147280 664190
rect 147520 663950 147630 664190
rect 147870 663950 147960 664190
rect 148200 663950 148290 664190
rect 148530 663950 148620 664190
rect 148860 663950 148970 664190
rect 149210 663950 149300 664190
rect 149540 663950 149630 664190
rect 149870 663950 149960 664190
rect 150200 663950 150310 664190
rect 150550 663950 150640 664190
rect 150880 663950 150970 664190
rect 151210 663950 151300 664190
rect 151540 663950 151650 664190
rect 151890 663950 151980 664190
rect 152220 663950 152310 664190
rect 152550 663950 152640 664190
rect 152880 663950 152990 664190
rect 153230 663950 153320 664190
rect 153560 663950 153650 664190
rect 153890 663950 153980 664190
rect 154220 663950 154330 664190
rect 154570 663950 154660 664190
rect 154900 663950 154990 664190
rect 155230 663950 155320 664190
rect 155560 663950 155670 664190
rect 155910 663950 155960 664190
rect 110760 663860 155960 663950
rect 110760 663620 110810 663860
rect 111050 663620 111140 663860
rect 111380 663620 111470 663860
rect 111710 663620 111800 663860
rect 112040 663620 112150 663860
rect 112390 663620 112480 663860
rect 112720 663620 112810 663860
rect 113050 663620 113140 663860
rect 113380 663620 113490 663860
rect 113730 663620 113820 663860
rect 114060 663620 114150 663860
rect 114390 663620 114480 663860
rect 114720 663620 114830 663860
rect 115070 663620 115160 663860
rect 115400 663620 115490 663860
rect 115730 663620 115820 663860
rect 116060 663620 116170 663860
rect 116410 663620 116500 663860
rect 116740 663620 116830 663860
rect 117070 663620 117160 663860
rect 117400 663620 117510 663860
rect 117750 663620 117840 663860
rect 118080 663620 118170 663860
rect 118410 663620 118500 663860
rect 118740 663620 118850 663860
rect 119090 663620 119180 663860
rect 119420 663620 119510 663860
rect 119750 663620 119840 663860
rect 120080 663620 120190 663860
rect 120430 663620 120520 663860
rect 120760 663620 120850 663860
rect 121090 663620 121180 663860
rect 121420 663620 121530 663860
rect 121770 663620 122190 663860
rect 122430 663620 122520 663860
rect 122760 663620 122850 663860
rect 123090 663620 123180 663860
rect 123420 663620 123530 663860
rect 123770 663620 123860 663860
rect 124100 663620 124190 663860
rect 124430 663620 124520 663860
rect 124760 663620 124870 663860
rect 125110 663620 125200 663860
rect 125440 663620 125530 663860
rect 125770 663620 125860 663860
rect 126100 663620 126210 663860
rect 126450 663620 126540 663860
rect 126780 663620 126870 663860
rect 127110 663620 127200 663860
rect 127440 663620 127550 663860
rect 127790 663620 127880 663860
rect 128120 663620 128210 663860
rect 128450 663620 128540 663860
rect 128780 663620 128890 663860
rect 129130 663620 129220 663860
rect 129460 663620 129550 663860
rect 129790 663620 129880 663860
rect 130120 663620 130230 663860
rect 130470 663620 130560 663860
rect 130800 663620 130890 663860
rect 131130 663620 131220 663860
rect 131460 663620 131570 663860
rect 131810 663620 131900 663860
rect 132140 663620 132230 663860
rect 132470 663620 132560 663860
rect 132800 663620 132910 663860
rect 133150 663620 133570 663860
rect 133810 663620 133900 663860
rect 134140 663620 134230 663860
rect 134470 663620 134560 663860
rect 134800 663620 134910 663860
rect 135150 663620 135240 663860
rect 135480 663620 135570 663860
rect 135810 663620 135900 663860
rect 136140 663620 136250 663860
rect 136490 663620 136580 663860
rect 136820 663620 136910 663860
rect 137150 663620 137240 663860
rect 137480 663620 137590 663860
rect 137830 663620 137920 663860
rect 138160 663620 138250 663860
rect 138490 663620 138580 663860
rect 138820 663620 138930 663860
rect 139170 663620 139260 663860
rect 139500 663620 139590 663860
rect 139830 663620 139920 663860
rect 140160 663620 140270 663860
rect 140510 663620 140600 663860
rect 140840 663620 140930 663860
rect 141170 663620 141260 663860
rect 141500 663620 141610 663860
rect 141850 663620 141940 663860
rect 142180 663620 142270 663860
rect 142510 663620 142600 663860
rect 142840 663620 142950 663860
rect 143190 663620 143280 663860
rect 143520 663620 143610 663860
rect 143850 663620 143940 663860
rect 144180 663620 144290 663860
rect 144530 663620 144950 663860
rect 145190 663620 145280 663860
rect 145520 663620 145610 663860
rect 145850 663620 145940 663860
rect 146180 663620 146290 663860
rect 146530 663620 146620 663860
rect 146860 663620 146950 663860
rect 147190 663620 147280 663860
rect 147520 663620 147630 663860
rect 147870 663620 147960 663860
rect 148200 663620 148290 663860
rect 148530 663620 148620 663860
rect 148860 663620 148970 663860
rect 149210 663620 149300 663860
rect 149540 663620 149630 663860
rect 149870 663620 149960 663860
rect 150200 663620 150310 663860
rect 150550 663620 150640 663860
rect 150880 663620 150970 663860
rect 151210 663620 151300 663860
rect 151540 663620 151650 663860
rect 151890 663620 151980 663860
rect 152220 663620 152310 663860
rect 152550 663620 152640 663860
rect 152880 663620 152990 663860
rect 153230 663620 153320 663860
rect 153560 663620 153650 663860
rect 153890 663620 153980 663860
rect 154220 663620 154330 663860
rect 154570 663620 154660 663860
rect 154900 663620 154990 663860
rect 155230 663620 155320 663860
rect 155560 663620 155670 663860
rect 155910 663620 155960 663860
rect 110760 663510 155960 663620
rect 110760 663270 110810 663510
rect 111050 663270 111140 663510
rect 111380 663270 111470 663510
rect 111710 663270 111800 663510
rect 112040 663270 112150 663510
rect 112390 663270 112480 663510
rect 112720 663270 112810 663510
rect 113050 663270 113140 663510
rect 113380 663270 113490 663510
rect 113730 663270 113820 663510
rect 114060 663270 114150 663510
rect 114390 663270 114480 663510
rect 114720 663270 114830 663510
rect 115070 663270 115160 663510
rect 115400 663270 115490 663510
rect 115730 663270 115820 663510
rect 116060 663270 116170 663510
rect 116410 663270 116500 663510
rect 116740 663270 116830 663510
rect 117070 663270 117160 663510
rect 117400 663270 117510 663510
rect 117750 663270 117840 663510
rect 118080 663270 118170 663510
rect 118410 663270 118500 663510
rect 118740 663270 118850 663510
rect 119090 663270 119180 663510
rect 119420 663270 119510 663510
rect 119750 663270 119840 663510
rect 120080 663270 120190 663510
rect 120430 663270 120520 663510
rect 120760 663270 120850 663510
rect 121090 663270 121180 663510
rect 121420 663270 121530 663510
rect 121770 663270 122190 663510
rect 122430 663270 122520 663510
rect 122760 663270 122850 663510
rect 123090 663270 123180 663510
rect 123420 663270 123530 663510
rect 123770 663270 123860 663510
rect 124100 663270 124190 663510
rect 124430 663270 124520 663510
rect 124760 663270 124870 663510
rect 125110 663270 125200 663510
rect 125440 663270 125530 663510
rect 125770 663270 125860 663510
rect 126100 663270 126210 663510
rect 126450 663270 126540 663510
rect 126780 663270 126870 663510
rect 127110 663270 127200 663510
rect 127440 663270 127550 663510
rect 127790 663270 127880 663510
rect 128120 663270 128210 663510
rect 128450 663270 128540 663510
rect 128780 663270 128890 663510
rect 129130 663270 129220 663510
rect 129460 663270 129550 663510
rect 129790 663270 129880 663510
rect 130120 663270 130230 663510
rect 130470 663270 130560 663510
rect 130800 663270 130890 663510
rect 131130 663270 131220 663510
rect 131460 663270 131570 663510
rect 131810 663270 131900 663510
rect 132140 663270 132230 663510
rect 132470 663270 132560 663510
rect 132800 663270 132910 663510
rect 133150 663270 133570 663510
rect 133810 663270 133900 663510
rect 134140 663270 134230 663510
rect 134470 663270 134560 663510
rect 134800 663270 134910 663510
rect 135150 663270 135240 663510
rect 135480 663270 135570 663510
rect 135810 663270 135900 663510
rect 136140 663270 136250 663510
rect 136490 663270 136580 663510
rect 136820 663270 136910 663510
rect 137150 663270 137240 663510
rect 137480 663270 137590 663510
rect 137830 663270 137920 663510
rect 138160 663270 138250 663510
rect 138490 663270 138580 663510
rect 138820 663270 138930 663510
rect 139170 663270 139260 663510
rect 139500 663270 139590 663510
rect 139830 663270 139920 663510
rect 140160 663270 140270 663510
rect 140510 663270 140600 663510
rect 140840 663270 140930 663510
rect 141170 663270 141260 663510
rect 141500 663270 141610 663510
rect 141850 663270 141940 663510
rect 142180 663270 142270 663510
rect 142510 663270 142600 663510
rect 142840 663270 142950 663510
rect 143190 663270 143280 663510
rect 143520 663270 143610 663510
rect 143850 663270 143940 663510
rect 144180 663270 144290 663510
rect 144530 663270 144950 663510
rect 145190 663270 145280 663510
rect 145520 663270 145610 663510
rect 145850 663270 145940 663510
rect 146180 663270 146290 663510
rect 146530 663270 146620 663510
rect 146860 663270 146950 663510
rect 147190 663270 147280 663510
rect 147520 663270 147630 663510
rect 147870 663270 147960 663510
rect 148200 663270 148290 663510
rect 148530 663270 148620 663510
rect 148860 663270 148970 663510
rect 149210 663270 149300 663510
rect 149540 663270 149630 663510
rect 149870 663270 149960 663510
rect 150200 663270 150310 663510
rect 150550 663270 150640 663510
rect 150880 663270 150970 663510
rect 151210 663270 151300 663510
rect 151540 663270 151650 663510
rect 151890 663270 151980 663510
rect 152220 663270 152310 663510
rect 152550 663270 152640 663510
rect 152880 663270 152990 663510
rect 153230 663270 153320 663510
rect 153560 663270 153650 663510
rect 153890 663270 153980 663510
rect 154220 663270 154330 663510
rect 154570 663270 154660 663510
rect 154900 663270 154990 663510
rect 155230 663270 155320 663510
rect 155560 663270 155670 663510
rect 155910 663270 155960 663510
rect 110760 663180 155960 663270
rect 110760 662940 110810 663180
rect 111050 662940 111140 663180
rect 111380 662940 111470 663180
rect 111710 662940 111800 663180
rect 112040 662940 112150 663180
rect 112390 662940 112480 663180
rect 112720 662940 112810 663180
rect 113050 662940 113140 663180
rect 113380 662940 113490 663180
rect 113730 662940 113820 663180
rect 114060 662940 114150 663180
rect 114390 662940 114480 663180
rect 114720 662940 114830 663180
rect 115070 662940 115160 663180
rect 115400 662940 115490 663180
rect 115730 662940 115820 663180
rect 116060 662940 116170 663180
rect 116410 662940 116500 663180
rect 116740 662940 116830 663180
rect 117070 662940 117160 663180
rect 117400 662940 117510 663180
rect 117750 662940 117840 663180
rect 118080 662940 118170 663180
rect 118410 662940 118500 663180
rect 118740 662940 118850 663180
rect 119090 662940 119180 663180
rect 119420 662940 119510 663180
rect 119750 662940 119840 663180
rect 120080 662940 120190 663180
rect 120430 662940 120520 663180
rect 120760 662940 120850 663180
rect 121090 662940 121180 663180
rect 121420 662940 121530 663180
rect 121770 662940 122190 663180
rect 122430 662940 122520 663180
rect 122760 662940 122850 663180
rect 123090 662940 123180 663180
rect 123420 662940 123530 663180
rect 123770 662940 123860 663180
rect 124100 662940 124190 663180
rect 124430 662940 124520 663180
rect 124760 662940 124870 663180
rect 125110 662940 125200 663180
rect 125440 662940 125530 663180
rect 125770 662940 125860 663180
rect 126100 662940 126210 663180
rect 126450 662940 126540 663180
rect 126780 662940 126870 663180
rect 127110 662940 127200 663180
rect 127440 662940 127550 663180
rect 127790 662940 127880 663180
rect 128120 662940 128210 663180
rect 128450 662940 128540 663180
rect 128780 662940 128890 663180
rect 129130 662940 129220 663180
rect 129460 662940 129550 663180
rect 129790 662940 129880 663180
rect 130120 662940 130230 663180
rect 130470 662940 130560 663180
rect 130800 662940 130890 663180
rect 131130 662940 131220 663180
rect 131460 662940 131570 663180
rect 131810 662940 131900 663180
rect 132140 662940 132230 663180
rect 132470 662940 132560 663180
rect 132800 662940 132910 663180
rect 133150 662940 133570 663180
rect 133810 662940 133900 663180
rect 134140 662940 134230 663180
rect 134470 662940 134560 663180
rect 134800 662940 134910 663180
rect 135150 662940 135240 663180
rect 135480 662940 135570 663180
rect 135810 662940 135900 663180
rect 136140 662940 136250 663180
rect 136490 662940 136580 663180
rect 136820 662940 136910 663180
rect 137150 662940 137240 663180
rect 137480 662940 137590 663180
rect 137830 662940 137920 663180
rect 138160 662940 138250 663180
rect 138490 662940 138580 663180
rect 138820 662940 138930 663180
rect 139170 662940 139260 663180
rect 139500 662940 139590 663180
rect 139830 662940 139920 663180
rect 140160 662940 140270 663180
rect 140510 662940 140600 663180
rect 140840 662940 140930 663180
rect 141170 662940 141260 663180
rect 141500 662940 141610 663180
rect 141850 662940 141940 663180
rect 142180 662940 142270 663180
rect 142510 662940 142600 663180
rect 142840 662940 142950 663180
rect 143190 662940 143280 663180
rect 143520 662940 143610 663180
rect 143850 662940 143940 663180
rect 144180 662940 144290 663180
rect 144530 662940 144950 663180
rect 145190 662940 145280 663180
rect 145520 662940 145610 663180
rect 145850 662940 145940 663180
rect 146180 662940 146290 663180
rect 146530 662940 146620 663180
rect 146860 662940 146950 663180
rect 147190 662940 147280 663180
rect 147520 662940 147630 663180
rect 147870 662940 147960 663180
rect 148200 662940 148290 663180
rect 148530 662940 148620 663180
rect 148860 662940 148970 663180
rect 149210 662940 149300 663180
rect 149540 662940 149630 663180
rect 149870 662940 149960 663180
rect 150200 662940 150310 663180
rect 150550 662940 150640 663180
rect 150880 662940 150970 663180
rect 151210 662940 151300 663180
rect 151540 662940 151650 663180
rect 151890 662940 151980 663180
rect 152220 662940 152310 663180
rect 152550 662940 152640 663180
rect 152880 662940 152990 663180
rect 153230 662940 153320 663180
rect 153560 662940 153650 663180
rect 153890 662940 153980 663180
rect 154220 662940 154330 663180
rect 154570 662940 154660 663180
rect 154900 662940 154990 663180
rect 155230 662940 155320 663180
rect 155560 662940 155670 663180
rect 155910 662940 155960 663180
rect 110760 662850 155960 662940
rect 110760 662610 110810 662850
rect 111050 662610 111140 662850
rect 111380 662610 111470 662850
rect 111710 662610 111800 662850
rect 112040 662610 112150 662850
rect 112390 662610 112480 662850
rect 112720 662610 112810 662850
rect 113050 662610 113140 662850
rect 113380 662610 113490 662850
rect 113730 662610 113820 662850
rect 114060 662610 114150 662850
rect 114390 662610 114480 662850
rect 114720 662610 114830 662850
rect 115070 662610 115160 662850
rect 115400 662610 115490 662850
rect 115730 662610 115820 662850
rect 116060 662610 116170 662850
rect 116410 662610 116500 662850
rect 116740 662610 116830 662850
rect 117070 662610 117160 662850
rect 117400 662610 117510 662850
rect 117750 662610 117840 662850
rect 118080 662610 118170 662850
rect 118410 662610 118500 662850
rect 118740 662610 118850 662850
rect 119090 662610 119180 662850
rect 119420 662610 119510 662850
rect 119750 662610 119840 662850
rect 120080 662610 120190 662850
rect 120430 662610 120520 662850
rect 120760 662610 120850 662850
rect 121090 662610 121180 662850
rect 121420 662610 121530 662850
rect 121770 662610 122190 662850
rect 122430 662610 122520 662850
rect 122760 662610 122850 662850
rect 123090 662610 123180 662850
rect 123420 662610 123530 662850
rect 123770 662610 123860 662850
rect 124100 662610 124190 662850
rect 124430 662610 124520 662850
rect 124760 662610 124870 662850
rect 125110 662610 125200 662850
rect 125440 662610 125530 662850
rect 125770 662610 125860 662850
rect 126100 662610 126210 662850
rect 126450 662610 126540 662850
rect 126780 662610 126870 662850
rect 127110 662610 127200 662850
rect 127440 662610 127550 662850
rect 127790 662610 127880 662850
rect 128120 662610 128210 662850
rect 128450 662610 128540 662850
rect 128780 662610 128890 662850
rect 129130 662610 129220 662850
rect 129460 662610 129550 662850
rect 129790 662610 129880 662850
rect 130120 662610 130230 662850
rect 130470 662610 130560 662850
rect 130800 662610 130890 662850
rect 131130 662610 131220 662850
rect 131460 662610 131570 662850
rect 131810 662610 131900 662850
rect 132140 662610 132230 662850
rect 132470 662610 132560 662850
rect 132800 662610 132910 662850
rect 133150 662610 133570 662850
rect 133810 662610 133900 662850
rect 134140 662610 134230 662850
rect 134470 662610 134560 662850
rect 134800 662610 134910 662850
rect 135150 662610 135240 662850
rect 135480 662610 135570 662850
rect 135810 662610 135900 662850
rect 136140 662610 136250 662850
rect 136490 662610 136580 662850
rect 136820 662610 136910 662850
rect 137150 662610 137240 662850
rect 137480 662610 137590 662850
rect 137830 662610 137920 662850
rect 138160 662610 138250 662850
rect 138490 662610 138580 662850
rect 138820 662610 138930 662850
rect 139170 662610 139260 662850
rect 139500 662610 139590 662850
rect 139830 662610 139920 662850
rect 140160 662610 140270 662850
rect 140510 662610 140600 662850
rect 140840 662610 140930 662850
rect 141170 662610 141260 662850
rect 141500 662610 141610 662850
rect 141850 662610 141940 662850
rect 142180 662610 142270 662850
rect 142510 662610 142600 662850
rect 142840 662610 142950 662850
rect 143190 662610 143280 662850
rect 143520 662610 143610 662850
rect 143850 662610 143940 662850
rect 144180 662610 144290 662850
rect 144530 662610 144950 662850
rect 145190 662610 145280 662850
rect 145520 662610 145610 662850
rect 145850 662610 145940 662850
rect 146180 662610 146290 662850
rect 146530 662610 146620 662850
rect 146860 662610 146950 662850
rect 147190 662610 147280 662850
rect 147520 662610 147630 662850
rect 147870 662610 147960 662850
rect 148200 662610 148290 662850
rect 148530 662610 148620 662850
rect 148860 662610 148970 662850
rect 149210 662610 149300 662850
rect 149540 662610 149630 662850
rect 149870 662610 149960 662850
rect 150200 662610 150310 662850
rect 150550 662610 150640 662850
rect 150880 662610 150970 662850
rect 151210 662610 151300 662850
rect 151540 662610 151650 662850
rect 151890 662610 151980 662850
rect 152220 662610 152310 662850
rect 152550 662610 152640 662850
rect 152880 662610 152990 662850
rect 153230 662610 153320 662850
rect 153560 662610 153650 662850
rect 153890 662610 153980 662850
rect 154220 662610 154330 662850
rect 154570 662610 154660 662850
rect 154900 662610 154990 662850
rect 155230 662610 155320 662850
rect 155560 662610 155670 662850
rect 155910 662610 155960 662850
rect 110760 662520 155960 662610
rect 110760 662280 110810 662520
rect 111050 662280 111140 662520
rect 111380 662280 111470 662520
rect 111710 662280 111800 662520
rect 112040 662280 112150 662520
rect 112390 662280 112480 662520
rect 112720 662280 112810 662520
rect 113050 662280 113140 662520
rect 113380 662280 113490 662520
rect 113730 662280 113820 662520
rect 114060 662280 114150 662520
rect 114390 662280 114480 662520
rect 114720 662280 114830 662520
rect 115070 662280 115160 662520
rect 115400 662280 115490 662520
rect 115730 662280 115820 662520
rect 116060 662280 116170 662520
rect 116410 662280 116500 662520
rect 116740 662280 116830 662520
rect 117070 662280 117160 662520
rect 117400 662280 117510 662520
rect 117750 662280 117840 662520
rect 118080 662280 118170 662520
rect 118410 662280 118500 662520
rect 118740 662280 118850 662520
rect 119090 662280 119180 662520
rect 119420 662280 119510 662520
rect 119750 662280 119840 662520
rect 120080 662280 120190 662520
rect 120430 662280 120520 662520
rect 120760 662280 120850 662520
rect 121090 662280 121180 662520
rect 121420 662280 121530 662520
rect 121770 662280 122190 662520
rect 122430 662280 122520 662520
rect 122760 662280 122850 662520
rect 123090 662280 123180 662520
rect 123420 662280 123530 662520
rect 123770 662280 123860 662520
rect 124100 662280 124190 662520
rect 124430 662280 124520 662520
rect 124760 662280 124870 662520
rect 125110 662280 125200 662520
rect 125440 662280 125530 662520
rect 125770 662280 125860 662520
rect 126100 662280 126210 662520
rect 126450 662280 126540 662520
rect 126780 662280 126870 662520
rect 127110 662280 127200 662520
rect 127440 662280 127550 662520
rect 127790 662280 127880 662520
rect 128120 662280 128210 662520
rect 128450 662280 128540 662520
rect 128780 662280 128890 662520
rect 129130 662280 129220 662520
rect 129460 662280 129550 662520
rect 129790 662280 129880 662520
rect 130120 662280 130230 662520
rect 130470 662280 130560 662520
rect 130800 662280 130890 662520
rect 131130 662280 131220 662520
rect 131460 662280 131570 662520
rect 131810 662280 131900 662520
rect 132140 662280 132230 662520
rect 132470 662280 132560 662520
rect 132800 662280 132910 662520
rect 133150 662280 133570 662520
rect 133810 662280 133900 662520
rect 134140 662280 134230 662520
rect 134470 662280 134560 662520
rect 134800 662280 134910 662520
rect 135150 662280 135240 662520
rect 135480 662280 135570 662520
rect 135810 662280 135900 662520
rect 136140 662280 136250 662520
rect 136490 662280 136580 662520
rect 136820 662280 136910 662520
rect 137150 662280 137240 662520
rect 137480 662280 137590 662520
rect 137830 662280 137920 662520
rect 138160 662280 138250 662520
rect 138490 662280 138580 662520
rect 138820 662280 138930 662520
rect 139170 662280 139260 662520
rect 139500 662280 139590 662520
rect 139830 662280 139920 662520
rect 140160 662280 140270 662520
rect 140510 662280 140600 662520
rect 140840 662280 140930 662520
rect 141170 662280 141260 662520
rect 141500 662280 141610 662520
rect 141850 662280 141940 662520
rect 142180 662280 142270 662520
rect 142510 662280 142600 662520
rect 142840 662280 142950 662520
rect 143190 662280 143280 662520
rect 143520 662280 143610 662520
rect 143850 662280 143940 662520
rect 144180 662280 144290 662520
rect 144530 662280 144950 662520
rect 145190 662280 145280 662520
rect 145520 662280 145610 662520
rect 145850 662280 145940 662520
rect 146180 662280 146290 662520
rect 146530 662280 146620 662520
rect 146860 662280 146950 662520
rect 147190 662280 147280 662520
rect 147520 662280 147630 662520
rect 147870 662280 147960 662520
rect 148200 662280 148290 662520
rect 148530 662280 148620 662520
rect 148860 662280 148970 662520
rect 149210 662280 149300 662520
rect 149540 662280 149630 662520
rect 149870 662280 149960 662520
rect 150200 662280 150310 662520
rect 150550 662280 150640 662520
rect 150880 662280 150970 662520
rect 151210 662280 151300 662520
rect 151540 662280 151650 662520
rect 151890 662280 151980 662520
rect 152220 662280 152310 662520
rect 152550 662280 152640 662520
rect 152880 662280 152990 662520
rect 153230 662280 153320 662520
rect 153560 662280 153650 662520
rect 153890 662280 153980 662520
rect 154220 662280 154330 662520
rect 154570 662280 154660 662520
rect 154900 662280 154990 662520
rect 155230 662280 155320 662520
rect 155560 662280 155670 662520
rect 155910 662280 155960 662520
rect 110760 662170 155960 662280
rect 110760 661930 110810 662170
rect 111050 661930 111140 662170
rect 111380 661930 111470 662170
rect 111710 661930 111800 662170
rect 112040 661930 112150 662170
rect 112390 661930 112480 662170
rect 112720 661930 112810 662170
rect 113050 661930 113140 662170
rect 113380 661930 113490 662170
rect 113730 661930 113820 662170
rect 114060 661930 114150 662170
rect 114390 661930 114480 662170
rect 114720 661930 114830 662170
rect 115070 661930 115160 662170
rect 115400 661930 115490 662170
rect 115730 661930 115820 662170
rect 116060 661930 116170 662170
rect 116410 661930 116500 662170
rect 116740 661930 116830 662170
rect 117070 661930 117160 662170
rect 117400 661930 117510 662170
rect 117750 661930 117840 662170
rect 118080 661930 118170 662170
rect 118410 661930 118500 662170
rect 118740 661930 118850 662170
rect 119090 661930 119180 662170
rect 119420 661930 119510 662170
rect 119750 661930 119840 662170
rect 120080 661930 120190 662170
rect 120430 661930 120520 662170
rect 120760 661930 120850 662170
rect 121090 661930 121180 662170
rect 121420 661930 121530 662170
rect 121770 661930 122190 662170
rect 122430 661930 122520 662170
rect 122760 661930 122850 662170
rect 123090 661930 123180 662170
rect 123420 661930 123530 662170
rect 123770 661930 123860 662170
rect 124100 661930 124190 662170
rect 124430 661930 124520 662170
rect 124760 661930 124870 662170
rect 125110 661930 125200 662170
rect 125440 661930 125530 662170
rect 125770 661930 125860 662170
rect 126100 661930 126210 662170
rect 126450 661930 126540 662170
rect 126780 661930 126870 662170
rect 127110 661930 127200 662170
rect 127440 661930 127550 662170
rect 127790 661930 127880 662170
rect 128120 661930 128210 662170
rect 128450 661930 128540 662170
rect 128780 661930 128890 662170
rect 129130 661930 129220 662170
rect 129460 661930 129550 662170
rect 129790 661930 129880 662170
rect 130120 661930 130230 662170
rect 130470 661930 130560 662170
rect 130800 661930 130890 662170
rect 131130 661930 131220 662170
rect 131460 661930 131570 662170
rect 131810 661930 131900 662170
rect 132140 661930 132230 662170
rect 132470 661930 132560 662170
rect 132800 661930 132910 662170
rect 133150 661930 133570 662170
rect 133810 661930 133900 662170
rect 134140 661930 134230 662170
rect 134470 661930 134560 662170
rect 134800 661930 134910 662170
rect 135150 661930 135240 662170
rect 135480 661930 135570 662170
rect 135810 661930 135900 662170
rect 136140 661930 136250 662170
rect 136490 661930 136580 662170
rect 136820 661930 136910 662170
rect 137150 661930 137240 662170
rect 137480 661930 137590 662170
rect 137830 661930 137920 662170
rect 138160 661930 138250 662170
rect 138490 661930 138580 662170
rect 138820 661930 138930 662170
rect 139170 661930 139260 662170
rect 139500 661930 139590 662170
rect 139830 661930 139920 662170
rect 140160 661930 140270 662170
rect 140510 661930 140600 662170
rect 140840 661930 140930 662170
rect 141170 661930 141260 662170
rect 141500 661930 141610 662170
rect 141850 661930 141940 662170
rect 142180 661930 142270 662170
rect 142510 661930 142600 662170
rect 142840 661930 142950 662170
rect 143190 661930 143280 662170
rect 143520 661930 143610 662170
rect 143850 661930 143940 662170
rect 144180 661930 144290 662170
rect 144530 661930 144950 662170
rect 145190 661930 145280 662170
rect 145520 661930 145610 662170
rect 145850 661930 145940 662170
rect 146180 661930 146290 662170
rect 146530 661930 146620 662170
rect 146860 661930 146950 662170
rect 147190 661930 147280 662170
rect 147520 661930 147630 662170
rect 147870 661930 147960 662170
rect 148200 661930 148290 662170
rect 148530 661930 148620 662170
rect 148860 661930 148970 662170
rect 149210 661930 149300 662170
rect 149540 661930 149630 662170
rect 149870 661930 149960 662170
rect 150200 661930 150310 662170
rect 150550 661930 150640 662170
rect 150880 661930 150970 662170
rect 151210 661930 151300 662170
rect 151540 661930 151650 662170
rect 151890 661930 151980 662170
rect 152220 661930 152310 662170
rect 152550 661930 152640 662170
rect 152880 661930 152990 662170
rect 153230 661930 153320 662170
rect 153560 661930 153650 662170
rect 153890 661930 153980 662170
rect 154220 661930 154330 662170
rect 154570 661930 154660 662170
rect 154900 661930 154990 662170
rect 155230 661930 155320 662170
rect 155560 661930 155670 662170
rect 155910 661930 155960 662170
rect 110760 661840 155960 661930
rect 110760 661600 110810 661840
rect 111050 661600 111140 661840
rect 111380 661600 111470 661840
rect 111710 661600 111800 661840
rect 112040 661600 112150 661840
rect 112390 661600 112480 661840
rect 112720 661600 112810 661840
rect 113050 661600 113140 661840
rect 113380 661600 113490 661840
rect 113730 661600 113820 661840
rect 114060 661600 114150 661840
rect 114390 661600 114480 661840
rect 114720 661600 114830 661840
rect 115070 661600 115160 661840
rect 115400 661600 115490 661840
rect 115730 661600 115820 661840
rect 116060 661600 116170 661840
rect 116410 661600 116500 661840
rect 116740 661600 116830 661840
rect 117070 661600 117160 661840
rect 117400 661600 117510 661840
rect 117750 661600 117840 661840
rect 118080 661600 118170 661840
rect 118410 661600 118500 661840
rect 118740 661600 118850 661840
rect 119090 661600 119180 661840
rect 119420 661600 119510 661840
rect 119750 661600 119840 661840
rect 120080 661600 120190 661840
rect 120430 661600 120520 661840
rect 120760 661600 120850 661840
rect 121090 661600 121180 661840
rect 121420 661600 121530 661840
rect 121770 661600 122190 661840
rect 122430 661600 122520 661840
rect 122760 661600 122850 661840
rect 123090 661600 123180 661840
rect 123420 661600 123530 661840
rect 123770 661600 123860 661840
rect 124100 661600 124190 661840
rect 124430 661600 124520 661840
rect 124760 661600 124870 661840
rect 125110 661600 125200 661840
rect 125440 661600 125530 661840
rect 125770 661600 125860 661840
rect 126100 661600 126210 661840
rect 126450 661600 126540 661840
rect 126780 661600 126870 661840
rect 127110 661600 127200 661840
rect 127440 661600 127550 661840
rect 127790 661600 127880 661840
rect 128120 661600 128210 661840
rect 128450 661600 128540 661840
rect 128780 661600 128890 661840
rect 129130 661600 129220 661840
rect 129460 661600 129550 661840
rect 129790 661600 129880 661840
rect 130120 661600 130230 661840
rect 130470 661600 130560 661840
rect 130800 661600 130890 661840
rect 131130 661600 131220 661840
rect 131460 661600 131570 661840
rect 131810 661600 131900 661840
rect 132140 661600 132230 661840
rect 132470 661600 132560 661840
rect 132800 661600 132910 661840
rect 133150 661600 133570 661840
rect 133810 661600 133900 661840
rect 134140 661600 134230 661840
rect 134470 661600 134560 661840
rect 134800 661600 134910 661840
rect 135150 661600 135240 661840
rect 135480 661600 135570 661840
rect 135810 661600 135900 661840
rect 136140 661600 136250 661840
rect 136490 661600 136580 661840
rect 136820 661600 136910 661840
rect 137150 661600 137240 661840
rect 137480 661600 137590 661840
rect 137830 661600 137920 661840
rect 138160 661600 138250 661840
rect 138490 661600 138580 661840
rect 138820 661600 138930 661840
rect 139170 661600 139260 661840
rect 139500 661600 139590 661840
rect 139830 661600 139920 661840
rect 140160 661600 140270 661840
rect 140510 661600 140600 661840
rect 140840 661600 140930 661840
rect 141170 661600 141260 661840
rect 141500 661600 141610 661840
rect 141850 661600 141940 661840
rect 142180 661600 142270 661840
rect 142510 661600 142600 661840
rect 142840 661600 142950 661840
rect 143190 661600 143280 661840
rect 143520 661600 143610 661840
rect 143850 661600 143940 661840
rect 144180 661600 144290 661840
rect 144530 661600 144950 661840
rect 145190 661600 145280 661840
rect 145520 661600 145610 661840
rect 145850 661600 145940 661840
rect 146180 661600 146290 661840
rect 146530 661600 146620 661840
rect 146860 661600 146950 661840
rect 147190 661600 147280 661840
rect 147520 661600 147630 661840
rect 147870 661600 147960 661840
rect 148200 661600 148290 661840
rect 148530 661600 148620 661840
rect 148860 661600 148970 661840
rect 149210 661600 149300 661840
rect 149540 661600 149630 661840
rect 149870 661600 149960 661840
rect 150200 661600 150310 661840
rect 150550 661600 150640 661840
rect 150880 661600 150970 661840
rect 151210 661600 151300 661840
rect 151540 661600 151650 661840
rect 151890 661600 151980 661840
rect 152220 661600 152310 661840
rect 152550 661600 152640 661840
rect 152880 661600 152990 661840
rect 153230 661600 153320 661840
rect 153560 661600 153650 661840
rect 153890 661600 153980 661840
rect 154220 661600 154330 661840
rect 154570 661600 154660 661840
rect 154900 661600 154990 661840
rect 155230 661600 155320 661840
rect 155560 661600 155670 661840
rect 155910 661600 155960 661840
rect 110760 661510 155960 661600
rect 110760 661270 110810 661510
rect 111050 661270 111140 661510
rect 111380 661270 111470 661510
rect 111710 661270 111800 661510
rect 112040 661270 112150 661510
rect 112390 661270 112480 661510
rect 112720 661270 112810 661510
rect 113050 661270 113140 661510
rect 113380 661270 113490 661510
rect 113730 661270 113820 661510
rect 114060 661270 114150 661510
rect 114390 661270 114480 661510
rect 114720 661270 114830 661510
rect 115070 661270 115160 661510
rect 115400 661270 115490 661510
rect 115730 661270 115820 661510
rect 116060 661270 116170 661510
rect 116410 661270 116500 661510
rect 116740 661270 116830 661510
rect 117070 661270 117160 661510
rect 117400 661270 117510 661510
rect 117750 661270 117840 661510
rect 118080 661270 118170 661510
rect 118410 661270 118500 661510
rect 118740 661270 118850 661510
rect 119090 661270 119180 661510
rect 119420 661270 119510 661510
rect 119750 661270 119840 661510
rect 120080 661270 120190 661510
rect 120430 661270 120520 661510
rect 120760 661270 120850 661510
rect 121090 661270 121180 661510
rect 121420 661270 121530 661510
rect 121770 661270 122190 661510
rect 122430 661270 122520 661510
rect 122760 661270 122850 661510
rect 123090 661270 123180 661510
rect 123420 661270 123530 661510
rect 123770 661270 123860 661510
rect 124100 661270 124190 661510
rect 124430 661270 124520 661510
rect 124760 661270 124870 661510
rect 125110 661270 125200 661510
rect 125440 661270 125530 661510
rect 125770 661270 125860 661510
rect 126100 661270 126210 661510
rect 126450 661270 126540 661510
rect 126780 661270 126870 661510
rect 127110 661270 127200 661510
rect 127440 661270 127550 661510
rect 127790 661270 127880 661510
rect 128120 661270 128210 661510
rect 128450 661270 128540 661510
rect 128780 661270 128890 661510
rect 129130 661270 129220 661510
rect 129460 661270 129550 661510
rect 129790 661270 129880 661510
rect 130120 661270 130230 661510
rect 130470 661270 130560 661510
rect 130800 661270 130890 661510
rect 131130 661270 131220 661510
rect 131460 661270 131570 661510
rect 131810 661270 131900 661510
rect 132140 661270 132230 661510
rect 132470 661270 132560 661510
rect 132800 661270 132910 661510
rect 133150 661270 133570 661510
rect 133810 661270 133900 661510
rect 134140 661270 134230 661510
rect 134470 661270 134560 661510
rect 134800 661270 134910 661510
rect 135150 661270 135240 661510
rect 135480 661270 135570 661510
rect 135810 661270 135900 661510
rect 136140 661270 136250 661510
rect 136490 661270 136580 661510
rect 136820 661270 136910 661510
rect 137150 661270 137240 661510
rect 137480 661270 137590 661510
rect 137830 661270 137920 661510
rect 138160 661270 138250 661510
rect 138490 661270 138580 661510
rect 138820 661270 138930 661510
rect 139170 661270 139260 661510
rect 139500 661270 139590 661510
rect 139830 661270 139920 661510
rect 140160 661270 140270 661510
rect 140510 661270 140600 661510
rect 140840 661270 140930 661510
rect 141170 661270 141260 661510
rect 141500 661270 141610 661510
rect 141850 661270 141940 661510
rect 142180 661270 142270 661510
rect 142510 661270 142600 661510
rect 142840 661270 142950 661510
rect 143190 661270 143280 661510
rect 143520 661270 143610 661510
rect 143850 661270 143940 661510
rect 144180 661270 144290 661510
rect 144530 661270 144950 661510
rect 145190 661270 145280 661510
rect 145520 661270 145610 661510
rect 145850 661270 145940 661510
rect 146180 661270 146290 661510
rect 146530 661270 146620 661510
rect 146860 661270 146950 661510
rect 147190 661270 147280 661510
rect 147520 661270 147630 661510
rect 147870 661270 147960 661510
rect 148200 661270 148290 661510
rect 148530 661270 148620 661510
rect 148860 661270 148970 661510
rect 149210 661270 149300 661510
rect 149540 661270 149630 661510
rect 149870 661270 149960 661510
rect 150200 661270 150310 661510
rect 150550 661270 150640 661510
rect 150880 661270 150970 661510
rect 151210 661270 151300 661510
rect 151540 661270 151650 661510
rect 151890 661270 151980 661510
rect 152220 661270 152310 661510
rect 152550 661270 152640 661510
rect 152880 661270 152990 661510
rect 153230 661270 153320 661510
rect 153560 661270 153650 661510
rect 153890 661270 153980 661510
rect 154220 661270 154330 661510
rect 154570 661270 154660 661510
rect 154900 661270 154990 661510
rect 155230 661270 155320 661510
rect 155560 661270 155670 661510
rect 155910 661270 155960 661510
rect 110760 661180 155960 661270
rect 110760 660940 110810 661180
rect 111050 660940 111140 661180
rect 111380 660940 111470 661180
rect 111710 660940 111800 661180
rect 112040 660940 112150 661180
rect 112390 660940 112480 661180
rect 112720 660940 112810 661180
rect 113050 660940 113140 661180
rect 113380 660940 113490 661180
rect 113730 660940 113820 661180
rect 114060 660940 114150 661180
rect 114390 660940 114480 661180
rect 114720 660940 114830 661180
rect 115070 660940 115160 661180
rect 115400 660940 115490 661180
rect 115730 660940 115820 661180
rect 116060 660940 116170 661180
rect 116410 660940 116500 661180
rect 116740 660940 116830 661180
rect 117070 660940 117160 661180
rect 117400 660940 117510 661180
rect 117750 660940 117840 661180
rect 118080 660940 118170 661180
rect 118410 660940 118500 661180
rect 118740 660940 118850 661180
rect 119090 660940 119180 661180
rect 119420 660940 119510 661180
rect 119750 660940 119840 661180
rect 120080 660940 120190 661180
rect 120430 660940 120520 661180
rect 120760 660940 120850 661180
rect 121090 660940 121180 661180
rect 121420 660940 121530 661180
rect 121770 660940 122190 661180
rect 122430 660940 122520 661180
rect 122760 660940 122850 661180
rect 123090 660940 123180 661180
rect 123420 660940 123530 661180
rect 123770 660940 123860 661180
rect 124100 660940 124190 661180
rect 124430 660940 124520 661180
rect 124760 660940 124870 661180
rect 125110 660940 125200 661180
rect 125440 660940 125530 661180
rect 125770 660940 125860 661180
rect 126100 660940 126210 661180
rect 126450 660940 126540 661180
rect 126780 660940 126870 661180
rect 127110 660940 127200 661180
rect 127440 660940 127550 661180
rect 127790 660940 127880 661180
rect 128120 660940 128210 661180
rect 128450 660940 128540 661180
rect 128780 660940 128890 661180
rect 129130 660940 129220 661180
rect 129460 660940 129550 661180
rect 129790 660940 129880 661180
rect 130120 660940 130230 661180
rect 130470 660940 130560 661180
rect 130800 660940 130890 661180
rect 131130 660940 131220 661180
rect 131460 660940 131570 661180
rect 131810 660940 131900 661180
rect 132140 660940 132230 661180
rect 132470 660940 132560 661180
rect 132800 660940 132910 661180
rect 133150 660940 133570 661180
rect 133810 660940 133900 661180
rect 134140 660940 134230 661180
rect 134470 660940 134560 661180
rect 134800 660940 134910 661180
rect 135150 660940 135240 661180
rect 135480 660940 135570 661180
rect 135810 660940 135900 661180
rect 136140 660940 136250 661180
rect 136490 660940 136580 661180
rect 136820 660940 136910 661180
rect 137150 660940 137240 661180
rect 137480 660940 137590 661180
rect 137830 660940 137920 661180
rect 138160 660940 138250 661180
rect 138490 660940 138580 661180
rect 138820 660940 138930 661180
rect 139170 660940 139260 661180
rect 139500 660940 139590 661180
rect 139830 660940 139920 661180
rect 140160 660940 140270 661180
rect 140510 660940 140600 661180
rect 140840 660940 140930 661180
rect 141170 660940 141260 661180
rect 141500 660940 141610 661180
rect 141850 660940 141940 661180
rect 142180 660940 142270 661180
rect 142510 660940 142600 661180
rect 142840 660940 142950 661180
rect 143190 660940 143280 661180
rect 143520 660940 143610 661180
rect 143850 660940 143940 661180
rect 144180 660940 144290 661180
rect 144530 660940 144950 661180
rect 145190 660940 145280 661180
rect 145520 660940 145610 661180
rect 145850 660940 145940 661180
rect 146180 660940 146290 661180
rect 146530 660940 146620 661180
rect 146860 660940 146950 661180
rect 147190 660940 147280 661180
rect 147520 660940 147630 661180
rect 147870 660940 147960 661180
rect 148200 660940 148290 661180
rect 148530 660940 148620 661180
rect 148860 660940 148970 661180
rect 149210 660940 149300 661180
rect 149540 660940 149630 661180
rect 149870 660940 149960 661180
rect 150200 660940 150310 661180
rect 150550 660940 150640 661180
rect 150880 660940 150970 661180
rect 151210 660940 151300 661180
rect 151540 660940 151650 661180
rect 151890 660940 151980 661180
rect 152220 660940 152310 661180
rect 152550 660940 152640 661180
rect 152880 660940 152990 661180
rect 153230 660940 153320 661180
rect 153560 660940 153650 661180
rect 153890 660940 153980 661180
rect 154220 660940 154330 661180
rect 154570 660940 154660 661180
rect 154900 660940 154990 661180
rect 155230 660940 155320 661180
rect 155560 660940 155670 661180
rect 155910 660940 155960 661180
rect 110760 660890 155960 660940
rect 121820 660790 122140 660800
rect 133200 660790 133520 660800
rect 144580 660790 144900 660800
rect 110760 660760 155960 660790
rect 110760 660520 110890 660760
rect 111130 660520 111220 660760
rect 111460 660520 111550 660760
rect 111790 660520 111880 660760
rect 112120 660520 112210 660760
rect 112450 660520 112540 660760
rect 112780 660520 112870 660760
rect 113110 660520 113200 660760
rect 113440 660520 113530 660760
rect 113770 660520 113860 660760
rect 114100 660520 114190 660760
rect 114430 660520 114520 660760
rect 114760 660520 114850 660760
rect 115090 660520 115180 660760
rect 115420 660520 115510 660760
rect 115750 660520 115840 660760
rect 116080 660520 116170 660760
rect 116410 660520 116500 660760
rect 116740 660520 116830 660760
rect 117070 660520 117160 660760
rect 117400 660520 117490 660760
rect 117730 660520 117820 660760
rect 118060 660520 118150 660760
rect 118390 660520 118480 660760
rect 118720 660520 118810 660760
rect 119050 660520 119140 660760
rect 119380 660520 119470 660760
rect 119710 660520 119800 660760
rect 120040 660520 120130 660760
rect 120370 660520 120460 660760
rect 120700 660520 120790 660760
rect 121030 660520 121120 660760
rect 121360 660520 121450 660760
rect 121690 660520 122270 660760
rect 122510 660520 122600 660760
rect 122840 660520 122930 660760
rect 123170 660520 123260 660760
rect 123500 660520 123590 660760
rect 123830 660520 123920 660760
rect 124160 660520 124250 660760
rect 124490 660520 124580 660760
rect 124820 660520 124910 660760
rect 125150 660520 125240 660760
rect 125480 660520 125570 660760
rect 125810 660520 125900 660760
rect 126140 660520 126230 660760
rect 126470 660520 126560 660760
rect 126800 660520 126890 660760
rect 127130 660520 127220 660760
rect 127460 660520 127550 660760
rect 127790 660520 127880 660760
rect 128120 660520 128210 660760
rect 128450 660520 128540 660760
rect 128780 660520 128870 660760
rect 129110 660520 129200 660760
rect 129440 660520 129530 660760
rect 129770 660520 129860 660760
rect 130100 660520 130190 660760
rect 130430 660520 130520 660760
rect 130760 660520 130850 660760
rect 131090 660520 131180 660760
rect 131420 660520 131510 660760
rect 131750 660520 131840 660760
rect 132080 660520 132170 660760
rect 132410 660520 132500 660760
rect 132740 660520 132830 660760
rect 133070 660520 133650 660760
rect 133890 660520 133980 660760
rect 134220 660520 134310 660760
rect 134550 660520 134640 660760
rect 134880 660520 134970 660760
rect 135210 660520 135300 660760
rect 135540 660520 135630 660760
rect 135870 660520 135960 660760
rect 136200 660520 136290 660760
rect 136530 660520 136620 660760
rect 136860 660520 136950 660760
rect 137190 660520 137280 660760
rect 137520 660520 137610 660760
rect 137850 660520 137940 660760
rect 138180 660520 138270 660760
rect 138510 660520 138600 660760
rect 138840 660520 138930 660760
rect 139170 660520 139260 660760
rect 139500 660520 139590 660760
rect 139830 660520 139920 660760
rect 140160 660520 140250 660760
rect 140490 660520 140580 660760
rect 140820 660520 140910 660760
rect 141150 660520 141240 660760
rect 141480 660520 141570 660760
rect 141810 660520 141900 660760
rect 142140 660520 142230 660760
rect 142470 660520 142560 660760
rect 142800 660520 142890 660760
rect 143130 660520 143220 660760
rect 143460 660520 143550 660760
rect 143790 660520 143880 660760
rect 144120 660520 144210 660760
rect 144450 660520 145030 660760
rect 145270 660520 145360 660760
rect 145600 660520 145690 660760
rect 145930 660520 146020 660760
rect 146260 660520 146350 660760
rect 146590 660520 146680 660760
rect 146920 660520 147010 660760
rect 147250 660520 147340 660760
rect 147580 660520 147670 660760
rect 147910 660520 148000 660760
rect 148240 660520 148330 660760
rect 148570 660520 148660 660760
rect 148900 660520 148990 660760
rect 149230 660520 149320 660760
rect 149560 660520 149650 660760
rect 149890 660520 149980 660760
rect 150220 660520 150310 660760
rect 150550 660520 150640 660760
rect 150880 660520 150970 660760
rect 151210 660520 151300 660760
rect 151540 660520 151630 660760
rect 151870 660520 151960 660760
rect 152200 660520 152290 660760
rect 152530 660520 152620 660760
rect 152860 660520 152950 660760
rect 153190 660520 153280 660760
rect 153520 660520 153610 660760
rect 153850 660520 153940 660760
rect 154180 660520 154270 660760
rect 154510 660520 154600 660760
rect 154840 660520 154930 660760
rect 155170 660520 155260 660760
rect 155500 660520 155590 660760
rect 155830 660520 155960 660760
rect 110760 660490 155960 660520
rect 121820 660480 122140 660490
rect 133200 660480 133520 660490
rect 144580 660480 144900 660490
rect 110760 660340 155960 660390
rect 110760 660100 110810 660340
rect 111050 660100 111160 660340
rect 111400 660100 111490 660340
rect 111730 660100 111820 660340
rect 112060 660100 112150 660340
rect 112390 660100 112500 660340
rect 112740 660100 112830 660340
rect 113070 660100 113160 660340
rect 113400 660100 113490 660340
rect 113730 660100 113840 660340
rect 114080 660100 114170 660340
rect 114410 660100 114500 660340
rect 114740 660100 114830 660340
rect 115070 660100 115180 660340
rect 115420 660100 115510 660340
rect 115750 660100 115840 660340
rect 116080 660100 116170 660340
rect 116410 660100 116520 660340
rect 116760 660100 116850 660340
rect 117090 660100 117180 660340
rect 117420 660100 117510 660340
rect 117750 660100 117860 660340
rect 118100 660100 118190 660340
rect 118430 660100 118520 660340
rect 118760 660100 118850 660340
rect 119090 660100 119200 660340
rect 119440 660100 119530 660340
rect 119770 660100 119860 660340
rect 120100 660100 120190 660340
rect 120430 660100 120540 660340
rect 120780 660100 120870 660340
rect 121110 660100 121200 660340
rect 121440 660100 121530 660340
rect 121770 660100 122190 660340
rect 122430 660100 122540 660340
rect 122780 660100 122870 660340
rect 123110 660100 123200 660340
rect 123440 660100 123530 660340
rect 123770 660100 123880 660340
rect 124120 660100 124210 660340
rect 124450 660100 124540 660340
rect 124780 660100 124870 660340
rect 125110 660100 125220 660340
rect 125460 660100 125550 660340
rect 125790 660100 125880 660340
rect 126120 660100 126210 660340
rect 126450 660100 126560 660340
rect 126800 660100 126890 660340
rect 127130 660100 127220 660340
rect 127460 660100 127550 660340
rect 127790 660100 127900 660340
rect 128140 660100 128230 660340
rect 128470 660100 128560 660340
rect 128800 660100 128890 660340
rect 129130 660100 129240 660340
rect 129480 660100 129570 660340
rect 129810 660100 129900 660340
rect 130140 660100 130230 660340
rect 130470 660100 130580 660340
rect 130820 660100 130910 660340
rect 131150 660100 131240 660340
rect 131480 660100 131570 660340
rect 131810 660100 131920 660340
rect 132160 660100 132250 660340
rect 132490 660100 132580 660340
rect 132820 660100 132910 660340
rect 133150 660100 133570 660340
rect 133810 660100 133920 660340
rect 134160 660100 134250 660340
rect 134490 660100 134580 660340
rect 134820 660100 134910 660340
rect 135150 660100 135260 660340
rect 135500 660100 135590 660340
rect 135830 660100 135920 660340
rect 136160 660100 136250 660340
rect 136490 660100 136600 660340
rect 136840 660100 136930 660340
rect 137170 660100 137260 660340
rect 137500 660100 137590 660340
rect 137830 660100 137940 660340
rect 138180 660100 138270 660340
rect 138510 660100 138600 660340
rect 138840 660100 138930 660340
rect 139170 660100 139280 660340
rect 139520 660100 139610 660340
rect 139850 660100 139940 660340
rect 140180 660100 140270 660340
rect 140510 660100 140620 660340
rect 140860 660100 140950 660340
rect 141190 660100 141280 660340
rect 141520 660100 141610 660340
rect 141850 660100 141960 660340
rect 142200 660100 142290 660340
rect 142530 660100 142620 660340
rect 142860 660100 142950 660340
rect 143190 660100 143300 660340
rect 143540 660100 143630 660340
rect 143870 660100 143960 660340
rect 144200 660100 144290 660340
rect 144530 660100 144950 660340
rect 145190 660100 145300 660340
rect 145540 660100 145630 660340
rect 145870 660100 145960 660340
rect 146200 660100 146290 660340
rect 146530 660100 146640 660340
rect 146880 660100 146970 660340
rect 147210 660100 147300 660340
rect 147540 660100 147630 660340
rect 147870 660100 147980 660340
rect 148220 660100 148310 660340
rect 148550 660100 148640 660340
rect 148880 660100 148970 660340
rect 149210 660100 149320 660340
rect 149560 660100 149650 660340
rect 149890 660100 149980 660340
rect 150220 660100 150310 660340
rect 150550 660100 150660 660340
rect 150900 660100 150990 660340
rect 151230 660100 151320 660340
rect 151560 660100 151650 660340
rect 151890 660100 152000 660340
rect 152240 660100 152330 660340
rect 152570 660100 152660 660340
rect 152900 660100 152990 660340
rect 153230 660100 153340 660340
rect 153580 660100 153670 660340
rect 153910 660100 154000 660340
rect 154240 660100 154330 660340
rect 154570 660100 154680 660340
rect 154920 660100 155010 660340
rect 155250 660100 155340 660340
rect 155580 660100 155670 660340
rect 155910 660100 155960 660340
rect 110760 660010 155960 660100
rect 110760 659770 110810 660010
rect 111050 659770 111160 660010
rect 111400 659770 111490 660010
rect 111730 659770 111820 660010
rect 112060 659770 112150 660010
rect 112390 659770 112500 660010
rect 112740 659770 112830 660010
rect 113070 659770 113160 660010
rect 113400 659770 113490 660010
rect 113730 659770 113840 660010
rect 114080 659770 114170 660010
rect 114410 659770 114500 660010
rect 114740 659770 114830 660010
rect 115070 659770 115180 660010
rect 115420 659770 115510 660010
rect 115750 659770 115840 660010
rect 116080 659770 116170 660010
rect 116410 659770 116520 660010
rect 116760 659770 116850 660010
rect 117090 659770 117180 660010
rect 117420 659770 117510 660010
rect 117750 659770 117860 660010
rect 118100 659770 118190 660010
rect 118430 659770 118520 660010
rect 118760 659770 118850 660010
rect 119090 659770 119200 660010
rect 119440 659770 119530 660010
rect 119770 659770 119860 660010
rect 120100 659770 120190 660010
rect 120430 659770 120540 660010
rect 120780 659770 120870 660010
rect 121110 659770 121200 660010
rect 121440 659770 121530 660010
rect 121770 659770 122190 660010
rect 122430 659770 122540 660010
rect 122780 659770 122870 660010
rect 123110 659770 123200 660010
rect 123440 659770 123530 660010
rect 123770 659770 123880 660010
rect 124120 659770 124210 660010
rect 124450 659770 124540 660010
rect 124780 659770 124870 660010
rect 125110 659770 125220 660010
rect 125460 659770 125550 660010
rect 125790 659770 125880 660010
rect 126120 659770 126210 660010
rect 126450 659770 126560 660010
rect 126800 659770 126890 660010
rect 127130 659770 127220 660010
rect 127460 659770 127550 660010
rect 127790 659770 127900 660010
rect 128140 659770 128230 660010
rect 128470 659770 128560 660010
rect 128800 659770 128890 660010
rect 129130 659770 129240 660010
rect 129480 659770 129570 660010
rect 129810 659770 129900 660010
rect 130140 659770 130230 660010
rect 130470 659770 130580 660010
rect 130820 659770 130910 660010
rect 131150 659770 131240 660010
rect 131480 659770 131570 660010
rect 131810 659770 131920 660010
rect 132160 659770 132250 660010
rect 132490 659770 132580 660010
rect 132820 659770 132910 660010
rect 133150 659770 133570 660010
rect 133810 659770 133920 660010
rect 134160 659770 134250 660010
rect 134490 659770 134580 660010
rect 134820 659770 134910 660010
rect 135150 659770 135260 660010
rect 135500 659770 135590 660010
rect 135830 659770 135920 660010
rect 136160 659770 136250 660010
rect 136490 659770 136600 660010
rect 136840 659770 136930 660010
rect 137170 659770 137260 660010
rect 137500 659770 137590 660010
rect 137830 659770 137940 660010
rect 138180 659770 138270 660010
rect 138510 659770 138600 660010
rect 138840 659770 138930 660010
rect 139170 659770 139280 660010
rect 139520 659770 139610 660010
rect 139850 659770 139940 660010
rect 140180 659770 140270 660010
rect 140510 659770 140620 660010
rect 140860 659770 140950 660010
rect 141190 659770 141280 660010
rect 141520 659770 141610 660010
rect 141850 659770 141960 660010
rect 142200 659770 142290 660010
rect 142530 659770 142620 660010
rect 142860 659770 142950 660010
rect 143190 659770 143300 660010
rect 143540 659770 143630 660010
rect 143870 659770 143960 660010
rect 144200 659770 144290 660010
rect 144530 659770 144950 660010
rect 145190 659770 145300 660010
rect 145540 659770 145630 660010
rect 145870 659770 145960 660010
rect 146200 659770 146290 660010
rect 146530 659770 146640 660010
rect 146880 659770 146970 660010
rect 147210 659770 147300 660010
rect 147540 659770 147630 660010
rect 147870 659770 147980 660010
rect 148220 659770 148310 660010
rect 148550 659770 148640 660010
rect 148880 659770 148970 660010
rect 149210 659770 149320 660010
rect 149560 659770 149650 660010
rect 149890 659770 149980 660010
rect 150220 659770 150310 660010
rect 150550 659770 150660 660010
rect 150900 659770 150990 660010
rect 151230 659770 151320 660010
rect 151560 659770 151650 660010
rect 151890 659770 152000 660010
rect 152240 659770 152330 660010
rect 152570 659770 152660 660010
rect 152900 659770 152990 660010
rect 153230 659770 153340 660010
rect 153580 659770 153670 660010
rect 153910 659770 154000 660010
rect 154240 659770 154330 660010
rect 154570 659770 154680 660010
rect 154920 659770 155010 660010
rect 155250 659770 155340 660010
rect 155580 659770 155670 660010
rect 155910 659770 155960 660010
rect 110760 659680 155960 659770
rect 110760 659440 110810 659680
rect 111050 659440 111160 659680
rect 111400 659440 111490 659680
rect 111730 659440 111820 659680
rect 112060 659440 112150 659680
rect 112390 659440 112500 659680
rect 112740 659440 112830 659680
rect 113070 659440 113160 659680
rect 113400 659440 113490 659680
rect 113730 659440 113840 659680
rect 114080 659440 114170 659680
rect 114410 659440 114500 659680
rect 114740 659440 114830 659680
rect 115070 659440 115180 659680
rect 115420 659440 115510 659680
rect 115750 659440 115840 659680
rect 116080 659440 116170 659680
rect 116410 659440 116520 659680
rect 116760 659440 116850 659680
rect 117090 659440 117180 659680
rect 117420 659440 117510 659680
rect 117750 659440 117860 659680
rect 118100 659440 118190 659680
rect 118430 659440 118520 659680
rect 118760 659440 118850 659680
rect 119090 659440 119200 659680
rect 119440 659440 119530 659680
rect 119770 659440 119860 659680
rect 120100 659440 120190 659680
rect 120430 659440 120540 659680
rect 120780 659440 120870 659680
rect 121110 659440 121200 659680
rect 121440 659440 121530 659680
rect 121770 659440 122190 659680
rect 122430 659440 122540 659680
rect 122780 659440 122870 659680
rect 123110 659440 123200 659680
rect 123440 659440 123530 659680
rect 123770 659440 123880 659680
rect 124120 659440 124210 659680
rect 124450 659440 124540 659680
rect 124780 659440 124870 659680
rect 125110 659440 125220 659680
rect 125460 659440 125550 659680
rect 125790 659440 125880 659680
rect 126120 659440 126210 659680
rect 126450 659440 126560 659680
rect 126800 659440 126890 659680
rect 127130 659440 127220 659680
rect 127460 659440 127550 659680
rect 127790 659440 127900 659680
rect 128140 659440 128230 659680
rect 128470 659440 128560 659680
rect 128800 659440 128890 659680
rect 129130 659440 129240 659680
rect 129480 659440 129570 659680
rect 129810 659440 129900 659680
rect 130140 659440 130230 659680
rect 130470 659440 130580 659680
rect 130820 659440 130910 659680
rect 131150 659440 131240 659680
rect 131480 659440 131570 659680
rect 131810 659440 131920 659680
rect 132160 659440 132250 659680
rect 132490 659440 132580 659680
rect 132820 659440 132910 659680
rect 133150 659440 133570 659680
rect 133810 659440 133920 659680
rect 134160 659440 134250 659680
rect 134490 659440 134580 659680
rect 134820 659440 134910 659680
rect 135150 659440 135260 659680
rect 135500 659440 135590 659680
rect 135830 659440 135920 659680
rect 136160 659440 136250 659680
rect 136490 659440 136600 659680
rect 136840 659440 136930 659680
rect 137170 659440 137260 659680
rect 137500 659440 137590 659680
rect 137830 659440 137940 659680
rect 138180 659440 138270 659680
rect 138510 659440 138600 659680
rect 138840 659440 138930 659680
rect 139170 659440 139280 659680
rect 139520 659440 139610 659680
rect 139850 659440 139940 659680
rect 140180 659440 140270 659680
rect 140510 659440 140620 659680
rect 140860 659440 140950 659680
rect 141190 659440 141280 659680
rect 141520 659440 141610 659680
rect 141850 659440 141960 659680
rect 142200 659440 142290 659680
rect 142530 659440 142620 659680
rect 142860 659440 142950 659680
rect 143190 659440 143300 659680
rect 143540 659440 143630 659680
rect 143870 659440 143960 659680
rect 144200 659440 144290 659680
rect 144530 659440 144950 659680
rect 145190 659440 145300 659680
rect 145540 659440 145630 659680
rect 145870 659440 145960 659680
rect 146200 659440 146290 659680
rect 146530 659440 146640 659680
rect 146880 659440 146970 659680
rect 147210 659440 147300 659680
rect 147540 659440 147630 659680
rect 147870 659440 147980 659680
rect 148220 659440 148310 659680
rect 148550 659440 148640 659680
rect 148880 659440 148970 659680
rect 149210 659440 149320 659680
rect 149560 659440 149650 659680
rect 149890 659440 149980 659680
rect 150220 659440 150310 659680
rect 150550 659440 150660 659680
rect 150900 659440 150990 659680
rect 151230 659440 151320 659680
rect 151560 659440 151650 659680
rect 151890 659440 152000 659680
rect 152240 659440 152330 659680
rect 152570 659440 152660 659680
rect 152900 659440 152990 659680
rect 153230 659440 153340 659680
rect 153580 659440 153670 659680
rect 153910 659440 154000 659680
rect 154240 659440 154330 659680
rect 154570 659440 154680 659680
rect 154920 659440 155010 659680
rect 155250 659440 155340 659680
rect 155580 659440 155670 659680
rect 155910 659440 155960 659680
rect 110760 659350 155960 659440
rect 110760 659110 110810 659350
rect 111050 659110 111160 659350
rect 111400 659110 111490 659350
rect 111730 659110 111820 659350
rect 112060 659110 112150 659350
rect 112390 659110 112500 659350
rect 112740 659110 112830 659350
rect 113070 659110 113160 659350
rect 113400 659110 113490 659350
rect 113730 659110 113840 659350
rect 114080 659110 114170 659350
rect 114410 659110 114500 659350
rect 114740 659110 114830 659350
rect 115070 659110 115180 659350
rect 115420 659110 115510 659350
rect 115750 659110 115840 659350
rect 116080 659110 116170 659350
rect 116410 659110 116520 659350
rect 116760 659110 116850 659350
rect 117090 659110 117180 659350
rect 117420 659110 117510 659350
rect 117750 659110 117860 659350
rect 118100 659110 118190 659350
rect 118430 659110 118520 659350
rect 118760 659110 118850 659350
rect 119090 659110 119200 659350
rect 119440 659110 119530 659350
rect 119770 659110 119860 659350
rect 120100 659110 120190 659350
rect 120430 659110 120540 659350
rect 120780 659110 120870 659350
rect 121110 659110 121200 659350
rect 121440 659110 121530 659350
rect 121770 659110 122190 659350
rect 122430 659110 122540 659350
rect 122780 659110 122870 659350
rect 123110 659110 123200 659350
rect 123440 659110 123530 659350
rect 123770 659110 123880 659350
rect 124120 659110 124210 659350
rect 124450 659110 124540 659350
rect 124780 659110 124870 659350
rect 125110 659110 125220 659350
rect 125460 659110 125550 659350
rect 125790 659110 125880 659350
rect 126120 659110 126210 659350
rect 126450 659110 126560 659350
rect 126800 659110 126890 659350
rect 127130 659110 127220 659350
rect 127460 659110 127550 659350
rect 127790 659110 127900 659350
rect 128140 659110 128230 659350
rect 128470 659110 128560 659350
rect 128800 659110 128890 659350
rect 129130 659110 129240 659350
rect 129480 659110 129570 659350
rect 129810 659110 129900 659350
rect 130140 659110 130230 659350
rect 130470 659110 130580 659350
rect 130820 659110 130910 659350
rect 131150 659110 131240 659350
rect 131480 659110 131570 659350
rect 131810 659110 131920 659350
rect 132160 659110 132250 659350
rect 132490 659110 132580 659350
rect 132820 659110 132910 659350
rect 133150 659110 133570 659350
rect 133810 659110 133920 659350
rect 134160 659110 134250 659350
rect 134490 659110 134580 659350
rect 134820 659110 134910 659350
rect 135150 659110 135260 659350
rect 135500 659110 135590 659350
rect 135830 659110 135920 659350
rect 136160 659110 136250 659350
rect 136490 659110 136600 659350
rect 136840 659110 136930 659350
rect 137170 659110 137260 659350
rect 137500 659110 137590 659350
rect 137830 659110 137940 659350
rect 138180 659110 138270 659350
rect 138510 659110 138600 659350
rect 138840 659110 138930 659350
rect 139170 659110 139280 659350
rect 139520 659110 139610 659350
rect 139850 659110 139940 659350
rect 140180 659110 140270 659350
rect 140510 659110 140620 659350
rect 140860 659110 140950 659350
rect 141190 659110 141280 659350
rect 141520 659110 141610 659350
rect 141850 659110 141960 659350
rect 142200 659110 142290 659350
rect 142530 659110 142620 659350
rect 142860 659110 142950 659350
rect 143190 659110 143300 659350
rect 143540 659110 143630 659350
rect 143870 659110 143960 659350
rect 144200 659110 144290 659350
rect 144530 659110 144950 659350
rect 145190 659110 145300 659350
rect 145540 659110 145630 659350
rect 145870 659110 145960 659350
rect 146200 659110 146290 659350
rect 146530 659110 146640 659350
rect 146880 659110 146970 659350
rect 147210 659110 147300 659350
rect 147540 659110 147630 659350
rect 147870 659110 147980 659350
rect 148220 659110 148310 659350
rect 148550 659110 148640 659350
rect 148880 659110 148970 659350
rect 149210 659110 149320 659350
rect 149560 659110 149650 659350
rect 149890 659110 149980 659350
rect 150220 659110 150310 659350
rect 150550 659110 150660 659350
rect 150900 659110 150990 659350
rect 151230 659110 151320 659350
rect 151560 659110 151650 659350
rect 151890 659110 152000 659350
rect 152240 659110 152330 659350
rect 152570 659110 152660 659350
rect 152900 659110 152990 659350
rect 153230 659110 153340 659350
rect 153580 659110 153670 659350
rect 153910 659110 154000 659350
rect 154240 659110 154330 659350
rect 154570 659110 154680 659350
rect 154920 659110 155010 659350
rect 155250 659110 155340 659350
rect 155580 659110 155670 659350
rect 155910 659110 155960 659350
rect 110760 659000 155960 659110
rect 110760 658760 110810 659000
rect 111050 658760 111160 659000
rect 111400 658760 111490 659000
rect 111730 658760 111820 659000
rect 112060 658760 112150 659000
rect 112390 658760 112500 659000
rect 112740 658760 112830 659000
rect 113070 658760 113160 659000
rect 113400 658760 113490 659000
rect 113730 658760 113840 659000
rect 114080 658760 114170 659000
rect 114410 658760 114500 659000
rect 114740 658760 114830 659000
rect 115070 658760 115180 659000
rect 115420 658760 115510 659000
rect 115750 658760 115840 659000
rect 116080 658760 116170 659000
rect 116410 658760 116520 659000
rect 116760 658760 116850 659000
rect 117090 658760 117180 659000
rect 117420 658760 117510 659000
rect 117750 658760 117860 659000
rect 118100 658760 118190 659000
rect 118430 658760 118520 659000
rect 118760 658760 118850 659000
rect 119090 658760 119200 659000
rect 119440 658760 119530 659000
rect 119770 658760 119860 659000
rect 120100 658760 120190 659000
rect 120430 658760 120540 659000
rect 120780 658760 120870 659000
rect 121110 658760 121200 659000
rect 121440 658760 121530 659000
rect 121770 658760 122190 659000
rect 122430 658760 122540 659000
rect 122780 658760 122870 659000
rect 123110 658760 123200 659000
rect 123440 658760 123530 659000
rect 123770 658760 123880 659000
rect 124120 658760 124210 659000
rect 124450 658760 124540 659000
rect 124780 658760 124870 659000
rect 125110 658760 125220 659000
rect 125460 658760 125550 659000
rect 125790 658760 125880 659000
rect 126120 658760 126210 659000
rect 126450 658760 126560 659000
rect 126800 658760 126890 659000
rect 127130 658760 127220 659000
rect 127460 658760 127550 659000
rect 127790 658760 127900 659000
rect 128140 658760 128230 659000
rect 128470 658760 128560 659000
rect 128800 658760 128890 659000
rect 129130 658760 129240 659000
rect 129480 658760 129570 659000
rect 129810 658760 129900 659000
rect 130140 658760 130230 659000
rect 130470 658760 130580 659000
rect 130820 658760 130910 659000
rect 131150 658760 131240 659000
rect 131480 658760 131570 659000
rect 131810 658760 131920 659000
rect 132160 658760 132250 659000
rect 132490 658760 132580 659000
rect 132820 658760 132910 659000
rect 133150 658760 133570 659000
rect 133810 658760 133920 659000
rect 134160 658760 134250 659000
rect 134490 658760 134580 659000
rect 134820 658760 134910 659000
rect 135150 658760 135260 659000
rect 135500 658760 135590 659000
rect 135830 658760 135920 659000
rect 136160 658760 136250 659000
rect 136490 658760 136600 659000
rect 136840 658760 136930 659000
rect 137170 658760 137260 659000
rect 137500 658760 137590 659000
rect 137830 658760 137940 659000
rect 138180 658760 138270 659000
rect 138510 658760 138600 659000
rect 138840 658760 138930 659000
rect 139170 658760 139280 659000
rect 139520 658760 139610 659000
rect 139850 658760 139940 659000
rect 140180 658760 140270 659000
rect 140510 658760 140620 659000
rect 140860 658760 140950 659000
rect 141190 658760 141280 659000
rect 141520 658760 141610 659000
rect 141850 658760 141960 659000
rect 142200 658760 142290 659000
rect 142530 658760 142620 659000
rect 142860 658760 142950 659000
rect 143190 658760 143300 659000
rect 143540 658760 143630 659000
rect 143870 658760 143960 659000
rect 144200 658760 144290 659000
rect 144530 658760 144950 659000
rect 145190 658760 145300 659000
rect 145540 658760 145630 659000
rect 145870 658760 145960 659000
rect 146200 658760 146290 659000
rect 146530 658760 146640 659000
rect 146880 658760 146970 659000
rect 147210 658760 147300 659000
rect 147540 658760 147630 659000
rect 147870 658760 147980 659000
rect 148220 658760 148310 659000
rect 148550 658760 148640 659000
rect 148880 658760 148970 659000
rect 149210 658760 149320 659000
rect 149560 658760 149650 659000
rect 149890 658760 149980 659000
rect 150220 658760 150310 659000
rect 150550 658760 150660 659000
rect 150900 658760 150990 659000
rect 151230 658760 151320 659000
rect 151560 658760 151650 659000
rect 151890 658760 152000 659000
rect 152240 658760 152330 659000
rect 152570 658760 152660 659000
rect 152900 658760 152990 659000
rect 153230 658760 153340 659000
rect 153580 658760 153670 659000
rect 153910 658760 154000 659000
rect 154240 658760 154330 659000
rect 154570 658760 154680 659000
rect 154920 658760 155010 659000
rect 155250 658760 155340 659000
rect 155580 658760 155670 659000
rect 155910 658760 155960 659000
rect 110760 658670 155960 658760
rect 110760 658430 110810 658670
rect 111050 658430 111160 658670
rect 111400 658430 111490 658670
rect 111730 658430 111820 658670
rect 112060 658430 112150 658670
rect 112390 658430 112500 658670
rect 112740 658430 112830 658670
rect 113070 658430 113160 658670
rect 113400 658430 113490 658670
rect 113730 658430 113840 658670
rect 114080 658430 114170 658670
rect 114410 658430 114500 658670
rect 114740 658430 114830 658670
rect 115070 658430 115180 658670
rect 115420 658430 115510 658670
rect 115750 658430 115840 658670
rect 116080 658430 116170 658670
rect 116410 658430 116520 658670
rect 116760 658430 116850 658670
rect 117090 658430 117180 658670
rect 117420 658430 117510 658670
rect 117750 658430 117860 658670
rect 118100 658430 118190 658670
rect 118430 658430 118520 658670
rect 118760 658430 118850 658670
rect 119090 658430 119200 658670
rect 119440 658430 119530 658670
rect 119770 658430 119860 658670
rect 120100 658430 120190 658670
rect 120430 658430 120540 658670
rect 120780 658430 120870 658670
rect 121110 658430 121200 658670
rect 121440 658430 121530 658670
rect 121770 658430 122190 658670
rect 122430 658430 122540 658670
rect 122780 658430 122870 658670
rect 123110 658430 123200 658670
rect 123440 658430 123530 658670
rect 123770 658430 123880 658670
rect 124120 658430 124210 658670
rect 124450 658430 124540 658670
rect 124780 658430 124870 658670
rect 125110 658430 125220 658670
rect 125460 658430 125550 658670
rect 125790 658430 125880 658670
rect 126120 658430 126210 658670
rect 126450 658430 126560 658670
rect 126800 658430 126890 658670
rect 127130 658430 127220 658670
rect 127460 658430 127550 658670
rect 127790 658430 127900 658670
rect 128140 658430 128230 658670
rect 128470 658430 128560 658670
rect 128800 658430 128890 658670
rect 129130 658430 129240 658670
rect 129480 658430 129570 658670
rect 129810 658430 129900 658670
rect 130140 658430 130230 658670
rect 130470 658430 130580 658670
rect 130820 658430 130910 658670
rect 131150 658430 131240 658670
rect 131480 658430 131570 658670
rect 131810 658430 131920 658670
rect 132160 658430 132250 658670
rect 132490 658430 132580 658670
rect 132820 658430 132910 658670
rect 133150 658430 133570 658670
rect 133810 658430 133920 658670
rect 134160 658430 134250 658670
rect 134490 658430 134580 658670
rect 134820 658430 134910 658670
rect 135150 658430 135260 658670
rect 135500 658430 135590 658670
rect 135830 658430 135920 658670
rect 136160 658430 136250 658670
rect 136490 658430 136600 658670
rect 136840 658430 136930 658670
rect 137170 658430 137260 658670
rect 137500 658430 137590 658670
rect 137830 658430 137940 658670
rect 138180 658430 138270 658670
rect 138510 658430 138600 658670
rect 138840 658430 138930 658670
rect 139170 658430 139280 658670
rect 139520 658430 139610 658670
rect 139850 658430 139940 658670
rect 140180 658430 140270 658670
rect 140510 658430 140620 658670
rect 140860 658430 140950 658670
rect 141190 658430 141280 658670
rect 141520 658430 141610 658670
rect 141850 658430 141960 658670
rect 142200 658430 142290 658670
rect 142530 658430 142620 658670
rect 142860 658430 142950 658670
rect 143190 658430 143300 658670
rect 143540 658430 143630 658670
rect 143870 658430 143960 658670
rect 144200 658430 144290 658670
rect 144530 658430 144950 658670
rect 145190 658430 145300 658670
rect 145540 658430 145630 658670
rect 145870 658430 145960 658670
rect 146200 658430 146290 658670
rect 146530 658430 146640 658670
rect 146880 658430 146970 658670
rect 147210 658430 147300 658670
rect 147540 658430 147630 658670
rect 147870 658430 147980 658670
rect 148220 658430 148310 658670
rect 148550 658430 148640 658670
rect 148880 658430 148970 658670
rect 149210 658430 149320 658670
rect 149560 658430 149650 658670
rect 149890 658430 149980 658670
rect 150220 658430 150310 658670
rect 150550 658430 150660 658670
rect 150900 658430 150990 658670
rect 151230 658430 151320 658670
rect 151560 658430 151650 658670
rect 151890 658430 152000 658670
rect 152240 658430 152330 658670
rect 152570 658430 152660 658670
rect 152900 658430 152990 658670
rect 153230 658430 153340 658670
rect 153580 658430 153670 658670
rect 153910 658430 154000 658670
rect 154240 658430 154330 658670
rect 154570 658430 154680 658670
rect 154920 658430 155010 658670
rect 155250 658430 155340 658670
rect 155580 658430 155670 658670
rect 155910 658430 155960 658670
rect 110760 658340 155960 658430
rect 110760 658100 110810 658340
rect 111050 658100 111160 658340
rect 111400 658100 111490 658340
rect 111730 658100 111820 658340
rect 112060 658100 112150 658340
rect 112390 658100 112500 658340
rect 112740 658100 112830 658340
rect 113070 658100 113160 658340
rect 113400 658100 113490 658340
rect 113730 658100 113840 658340
rect 114080 658100 114170 658340
rect 114410 658100 114500 658340
rect 114740 658100 114830 658340
rect 115070 658100 115180 658340
rect 115420 658100 115510 658340
rect 115750 658100 115840 658340
rect 116080 658100 116170 658340
rect 116410 658100 116520 658340
rect 116760 658100 116850 658340
rect 117090 658100 117180 658340
rect 117420 658100 117510 658340
rect 117750 658100 117860 658340
rect 118100 658100 118190 658340
rect 118430 658100 118520 658340
rect 118760 658100 118850 658340
rect 119090 658100 119200 658340
rect 119440 658100 119530 658340
rect 119770 658100 119860 658340
rect 120100 658100 120190 658340
rect 120430 658100 120540 658340
rect 120780 658100 120870 658340
rect 121110 658100 121200 658340
rect 121440 658100 121530 658340
rect 121770 658100 122190 658340
rect 122430 658100 122540 658340
rect 122780 658100 122870 658340
rect 123110 658100 123200 658340
rect 123440 658100 123530 658340
rect 123770 658100 123880 658340
rect 124120 658100 124210 658340
rect 124450 658100 124540 658340
rect 124780 658100 124870 658340
rect 125110 658100 125220 658340
rect 125460 658100 125550 658340
rect 125790 658100 125880 658340
rect 126120 658100 126210 658340
rect 126450 658100 126560 658340
rect 126800 658100 126890 658340
rect 127130 658100 127220 658340
rect 127460 658100 127550 658340
rect 127790 658100 127900 658340
rect 128140 658100 128230 658340
rect 128470 658100 128560 658340
rect 128800 658100 128890 658340
rect 129130 658100 129240 658340
rect 129480 658100 129570 658340
rect 129810 658100 129900 658340
rect 130140 658100 130230 658340
rect 130470 658100 130580 658340
rect 130820 658100 130910 658340
rect 131150 658100 131240 658340
rect 131480 658100 131570 658340
rect 131810 658100 131920 658340
rect 132160 658100 132250 658340
rect 132490 658100 132580 658340
rect 132820 658100 132910 658340
rect 133150 658100 133570 658340
rect 133810 658100 133920 658340
rect 134160 658100 134250 658340
rect 134490 658100 134580 658340
rect 134820 658100 134910 658340
rect 135150 658100 135260 658340
rect 135500 658100 135590 658340
rect 135830 658100 135920 658340
rect 136160 658100 136250 658340
rect 136490 658100 136600 658340
rect 136840 658100 136930 658340
rect 137170 658100 137260 658340
rect 137500 658100 137590 658340
rect 137830 658100 137940 658340
rect 138180 658100 138270 658340
rect 138510 658100 138600 658340
rect 138840 658100 138930 658340
rect 139170 658100 139280 658340
rect 139520 658100 139610 658340
rect 139850 658100 139940 658340
rect 140180 658100 140270 658340
rect 140510 658100 140620 658340
rect 140860 658100 140950 658340
rect 141190 658100 141280 658340
rect 141520 658100 141610 658340
rect 141850 658100 141960 658340
rect 142200 658100 142290 658340
rect 142530 658100 142620 658340
rect 142860 658100 142950 658340
rect 143190 658100 143300 658340
rect 143540 658100 143630 658340
rect 143870 658100 143960 658340
rect 144200 658100 144290 658340
rect 144530 658100 144950 658340
rect 145190 658100 145300 658340
rect 145540 658100 145630 658340
rect 145870 658100 145960 658340
rect 146200 658100 146290 658340
rect 146530 658100 146640 658340
rect 146880 658100 146970 658340
rect 147210 658100 147300 658340
rect 147540 658100 147630 658340
rect 147870 658100 147980 658340
rect 148220 658100 148310 658340
rect 148550 658100 148640 658340
rect 148880 658100 148970 658340
rect 149210 658100 149320 658340
rect 149560 658100 149650 658340
rect 149890 658100 149980 658340
rect 150220 658100 150310 658340
rect 150550 658100 150660 658340
rect 150900 658100 150990 658340
rect 151230 658100 151320 658340
rect 151560 658100 151650 658340
rect 151890 658100 152000 658340
rect 152240 658100 152330 658340
rect 152570 658100 152660 658340
rect 152900 658100 152990 658340
rect 153230 658100 153340 658340
rect 153580 658100 153670 658340
rect 153910 658100 154000 658340
rect 154240 658100 154330 658340
rect 154570 658100 154680 658340
rect 154920 658100 155010 658340
rect 155250 658100 155340 658340
rect 155580 658100 155670 658340
rect 155910 658100 155960 658340
rect 110760 658010 155960 658100
rect 110760 657770 110810 658010
rect 111050 657770 111160 658010
rect 111400 657770 111490 658010
rect 111730 657770 111820 658010
rect 112060 657770 112150 658010
rect 112390 657770 112500 658010
rect 112740 657770 112830 658010
rect 113070 657770 113160 658010
rect 113400 657770 113490 658010
rect 113730 657770 113840 658010
rect 114080 657770 114170 658010
rect 114410 657770 114500 658010
rect 114740 657770 114830 658010
rect 115070 657770 115180 658010
rect 115420 657770 115510 658010
rect 115750 657770 115840 658010
rect 116080 657770 116170 658010
rect 116410 657770 116520 658010
rect 116760 657770 116850 658010
rect 117090 657770 117180 658010
rect 117420 657770 117510 658010
rect 117750 657770 117860 658010
rect 118100 657770 118190 658010
rect 118430 657770 118520 658010
rect 118760 657770 118850 658010
rect 119090 657770 119200 658010
rect 119440 657770 119530 658010
rect 119770 657770 119860 658010
rect 120100 657770 120190 658010
rect 120430 657770 120540 658010
rect 120780 657770 120870 658010
rect 121110 657770 121200 658010
rect 121440 657770 121530 658010
rect 121770 657770 122190 658010
rect 122430 657770 122540 658010
rect 122780 657770 122870 658010
rect 123110 657770 123200 658010
rect 123440 657770 123530 658010
rect 123770 657770 123880 658010
rect 124120 657770 124210 658010
rect 124450 657770 124540 658010
rect 124780 657770 124870 658010
rect 125110 657770 125220 658010
rect 125460 657770 125550 658010
rect 125790 657770 125880 658010
rect 126120 657770 126210 658010
rect 126450 657770 126560 658010
rect 126800 657770 126890 658010
rect 127130 657770 127220 658010
rect 127460 657770 127550 658010
rect 127790 657770 127900 658010
rect 128140 657770 128230 658010
rect 128470 657770 128560 658010
rect 128800 657770 128890 658010
rect 129130 657770 129240 658010
rect 129480 657770 129570 658010
rect 129810 657770 129900 658010
rect 130140 657770 130230 658010
rect 130470 657770 130580 658010
rect 130820 657770 130910 658010
rect 131150 657770 131240 658010
rect 131480 657770 131570 658010
rect 131810 657770 131920 658010
rect 132160 657770 132250 658010
rect 132490 657770 132580 658010
rect 132820 657770 132910 658010
rect 133150 657770 133570 658010
rect 133810 657770 133920 658010
rect 134160 657770 134250 658010
rect 134490 657770 134580 658010
rect 134820 657770 134910 658010
rect 135150 657770 135260 658010
rect 135500 657770 135590 658010
rect 135830 657770 135920 658010
rect 136160 657770 136250 658010
rect 136490 657770 136600 658010
rect 136840 657770 136930 658010
rect 137170 657770 137260 658010
rect 137500 657770 137590 658010
rect 137830 657770 137940 658010
rect 138180 657770 138270 658010
rect 138510 657770 138600 658010
rect 138840 657770 138930 658010
rect 139170 657770 139280 658010
rect 139520 657770 139610 658010
rect 139850 657770 139940 658010
rect 140180 657770 140270 658010
rect 140510 657770 140620 658010
rect 140860 657770 140950 658010
rect 141190 657770 141280 658010
rect 141520 657770 141610 658010
rect 141850 657770 141960 658010
rect 142200 657770 142290 658010
rect 142530 657770 142620 658010
rect 142860 657770 142950 658010
rect 143190 657770 143300 658010
rect 143540 657770 143630 658010
rect 143870 657770 143960 658010
rect 144200 657770 144290 658010
rect 144530 657770 144950 658010
rect 145190 657770 145300 658010
rect 145540 657770 145630 658010
rect 145870 657770 145960 658010
rect 146200 657770 146290 658010
rect 146530 657770 146640 658010
rect 146880 657770 146970 658010
rect 147210 657770 147300 658010
rect 147540 657770 147630 658010
rect 147870 657770 147980 658010
rect 148220 657770 148310 658010
rect 148550 657770 148640 658010
rect 148880 657770 148970 658010
rect 149210 657770 149320 658010
rect 149560 657770 149650 658010
rect 149890 657770 149980 658010
rect 150220 657770 150310 658010
rect 150550 657770 150660 658010
rect 150900 657770 150990 658010
rect 151230 657770 151320 658010
rect 151560 657770 151650 658010
rect 151890 657770 152000 658010
rect 152240 657770 152330 658010
rect 152570 657770 152660 658010
rect 152900 657770 152990 658010
rect 153230 657770 153340 658010
rect 153580 657770 153670 658010
rect 153910 657770 154000 658010
rect 154240 657770 154330 658010
rect 154570 657770 154680 658010
rect 154920 657770 155010 658010
rect 155250 657770 155340 658010
rect 155580 657770 155670 658010
rect 155910 657770 155960 658010
rect 110760 657660 155960 657770
rect 110760 657627 110810 657660
rect 103643 657420 110810 657627
rect 111050 657420 111160 657660
rect 111400 657420 111490 657660
rect 111730 657420 111820 657660
rect 112060 657420 112150 657660
rect 112390 657420 112500 657660
rect 112740 657420 112830 657660
rect 113070 657420 113160 657660
rect 113400 657420 113490 657660
rect 113730 657420 113840 657660
rect 114080 657420 114170 657660
rect 114410 657420 114500 657660
rect 114740 657420 114830 657660
rect 115070 657420 115180 657660
rect 115420 657420 115510 657660
rect 115750 657420 115840 657660
rect 116080 657420 116170 657660
rect 116410 657420 116520 657660
rect 116760 657420 116850 657660
rect 117090 657420 117180 657660
rect 117420 657420 117510 657660
rect 117750 657420 117860 657660
rect 118100 657420 118190 657660
rect 118430 657420 118520 657660
rect 118760 657420 118850 657660
rect 119090 657420 119200 657660
rect 119440 657420 119530 657660
rect 119770 657420 119860 657660
rect 120100 657420 120190 657660
rect 120430 657420 120540 657660
rect 120780 657420 120870 657660
rect 121110 657420 121200 657660
rect 121440 657420 121530 657660
rect 121770 657420 122190 657660
rect 122430 657420 122540 657660
rect 122780 657420 122870 657660
rect 123110 657420 123200 657660
rect 123440 657420 123530 657660
rect 123770 657420 123880 657660
rect 124120 657420 124210 657660
rect 124450 657420 124540 657660
rect 124780 657420 124870 657660
rect 125110 657420 125220 657660
rect 125460 657420 125550 657660
rect 125790 657420 125880 657660
rect 126120 657420 126210 657660
rect 126450 657420 126560 657660
rect 126800 657420 126890 657660
rect 127130 657420 127220 657660
rect 127460 657420 127550 657660
rect 127790 657420 127900 657660
rect 128140 657420 128230 657660
rect 128470 657420 128560 657660
rect 128800 657420 128890 657660
rect 129130 657420 129240 657660
rect 129480 657420 129570 657660
rect 129810 657420 129900 657660
rect 130140 657420 130230 657660
rect 130470 657420 130580 657660
rect 130820 657420 130910 657660
rect 131150 657420 131240 657660
rect 131480 657420 131570 657660
rect 131810 657420 131920 657660
rect 132160 657420 132250 657660
rect 132490 657420 132580 657660
rect 132820 657420 132910 657660
rect 133150 657420 133570 657660
rect 133810 657420 133920 657660
rect 134160 657420 134250 657660
rect 134490 657420 134580 657660
rect 134820 657420 134910 657660
rect 135150 657420 135260 657660
rect 135500 657420 135590 657660
rect 135830 657420 135920 657660
rect 136160 657420 136250 657660
rect 136490 657420 136600 657660
rect 136840 657420 136930 657660
rect 137170 657420 137260 657660
rect 137500 657420 137590 657660
rect 137830 657420 137940 657660
rect 138180 657420 138270 657660
rect 138510 657420 138600 657660
rect 138840 657420 138930 657660
rect 139170 657420 139280 657660
rect 139520 657420 139610 657660
rect 139850 657420 139940 657660
rect 140180 657420 140270 657660
rect 140510 657420 140620 657660
rect 140860 657420 140950 657660
rect 141190 657420 141280 657660
rect 141520 657420 141610 657660
rect 141850 657420 141960 657660
rect 142200 657420 142290 657660
rect 142530 657420 142620 657660
rect 142860 657420 142950 657660
rect 143190 657420 143300 657660
rect 143540 657420 143630 657660
rect 143870 657420 143960 657660
rect 144200 657420 144290 657660
rect 144530 657420 144950 657660
rect 145190 657420 145300 657660
rect 145540 657420 145630 657660
rect 145870 657420 145960 657660
rect 146200 657420 146290 657660
rect 146530 657420 146640 657660
rect 146880 657420 146970 657660
rect 147210 657420 147300 657660
rect 147540 657420 147630 657660
rect 147870 657420 147980 657660
rect 148220 657420 148310 657660
rect 148550 657420 148640 657660
rect 148880 657420 148970 657660
rect 149210 657420 149320 657660
rect 149560 657420 149650 657660
rect 149890 657420 149980 657660
rect 150220 657420 150310 657660
rect 150550 657420 150660 657660
rect 150900 657420 150990 657660
rect 151230 657420 151320 657660
rect 151560 657420 151650 657660
rect 151890 657420 152000 657660
rect 152240 657420 152330 657660
rect 152570 657420 152660 657660
rect 152900 657420 152990 657660
rect 153230 657420 153340 657660
rect 153580 657420 153670 657660
rect 153910 657420 154000 657660
rect 154240 657420 154330 657660
rect 154570 657420 154680 657660
rect 154920 657420 155010 657660
rect 155250 657420 155340 657660
rect 155580 657420 155670 657660
rect 155910 657627 155960 657660
rect 157440 657627 162436 674152
rect 467200 660850 467520 703060
rect 222414 660530 467520 660850
rect 569580 702870 569900 702890
rect 569580 702800 569600 702870
rect 569670 702800 569700 702870
rect 569770 702800 569800 702870
rect 569870 702800 569900 702870
rect 569580 702770 569900 702800
rect 569580 702700 569600 702770
rect 569670 702700 569700 702770
rect 569770 702700 569800 702770
rect 569870 702700 569900 702770
rect 569580 702670 569900 702700
rect 569580 702600 569600 702670
rect 569670 702600 569700 702670
rect 569770 702600 569800 702670
rect 569870 702600 569900 702670
rect 155910 657420 162436 657627
rect 103643 657330 162436 657420
rect 103643 657090 110810 657330
rect 111050 657090 111160 657330
rect 111400 657090 111490 657330
rect 111730 657090 111820 657330
rect 112060 657090 112150 657330
rect 112390 657090 112500 657330
rect 112740 657090 112830 657330
rect 113070 657090 113160 657330
rect 113400 657090 113490 657330
rect 113730 657090 113840 657330
rect 114080 657090 114170 657330
rect 114410 657090 114500 657330
rect 114740 657090 114830 657330
rect 115070 657090 115180 657330
rect 115420 657090 115510 657330
rect 115750 657090 115840 657330
rect 116080 657090 116170 657330
rect 116410 657090 116520 657330
rect 116760 657090 116850 657330
rect 117090 657090 117180 657330
rect 117420 657090 117510 657330
rect 117750 657090 117860 657330
rect 118100 657090 118190 657330
rect 118430 657090 118520 657330
rect 118760 657090 118850 657330
rect 119090 657090 119200 657330
rect 119440 657090 119530 657330
rect 119770 657090 119860 657330
rect 120100 657090 120190 657330
rect 120430 657090 120540 657330
rect 120780 657090 120870 657330
rect 121110 657090 121200 657330
rect 121440 657090 121530 657330
rect 121770 657090 122190 657330
rect 122430 657090 122540 657330
rect 122780 657090 122870 657330
rect 123110 657090 123200 657330
rect 123440 657090 123530 657330
rect 123770 657090 123880 657330
rect 124120 657090 124210 657330
rect 124450 657090 124540 657330
rect 124780 657090 124870 657330
rect 125110 657090 125220 657330
rect 125460 657090 125550 657330
rect 125790 657090 125880 657330
rect 126120 657090 126210 657330
rect 126450 657090 126560 657330
rect 126800 657090 126890 657330
rect 127130 657090 127220 657330
rect 127460 657090 127550 657330
rect 127790 657090 127900 657330
rect 128140 657090 128230 657330
rect 128470 657090 128560 657330
rect 128800 657090 128890 657330
rect 129130 657090 129240 657330
rect 129480 657090 129570 657330
rect 129810 657090 129900 657330
rect 130140 657090 130230 657330
rect 130470 657090 130580 657330
rect 130820 657090 130910 657330
rect 131150 657090 131240 657330
rect 131480 657090 131570 657330
rect 131810 657090 131920 657330
rect 132160 657090 132250 657330
rect 132490 657090 132580 657330
rect 132820 657090 132910 657330
rect 133150 657090 133570 657330
rect 133810 657090 133920 657330
rect 134160 657090 134250 657330
rect 134490 657090 134580 657330
rect 134820 657090 134910 657330
rect 135150 657090 135260 657330
rect 135500 657090 135590 657330
rect 135830 657090 135920 657330
rect 136160 657090 136250 657330
rect 136490 657090 136600 657330
rect 136840 657090 136930 657330
rect 137170 657090 137260 657330
rect 137500 657090 137590 657330
rect 137830 657090 137940 657330
rect 138180 657090 138270 657330
rect 138510 657090 138600 657330
rect 138840 657090 138930 657330
rect 139170 657090 139280 657330
rect 139520 657090 139610 657330
rect 139850 657090 139940 657330
rect 140180 657090 140270 657330
rect 140510 657090 140620 657330
rect 140860 657090 140950 657330
rect 141190 657090 141280 657330
rect 141520 657090 141610 657330
rect 141850 657090 141960 657330
rect 142200 657090 142290 657330
rect 142530 657090 142620 657330
rect 142860 657090 142950 657330
rect 143190 657090 143300 657330
rect 143540 657090 143630 657330
rect 143870 657090 143960 657330
rect 144200 657090 144290 657330
rect 144530 657090 144950 657330
rect 145190 657090 145300 657330
rect 145540 657090 145630 657330
rect 145870 657090 145960 657330
rect 146200 657090 146290 657330
rect 146530 657090 146640 657330
rect 146880 657090 146970 657330
rect 147210 657090 147300 657330
rect 147540 657090 147630 657330
rect 147870 657090 147980 657330
rect 148220 657090 148310 657330
rect 148550 657090 148640 657330
rect 148880 657090 148970 657330
rect 149210 657090 149320 657330
rect 149560 657090 149650 657330
rect 149890 657090 149980 657330
rect 150220 657090 150310 657330
rect 150550 657090 150660 657330
rect 150900 657090 150990 657330
rect 151230 657090 151320 657330
rect 151560 657090 151650 657330
rect 151890 657090 152000 657330
rect 152240 657090 152330 657330
rect 152570 657090 152660 657330
rect 152900 657090 152990 657330
rect 153230 657090 153340 657330
rect 153580 657090 153670 657330
rect 153910 657090 154000 657330
rect 154240 657090 154330 657330
rect 154570 657090 154680 657330
rect 154920 657090 155010 657330
rect 155250 657090 155340 657330
rect 155580 657090 155670 657330
rect 155910 657090 162436 657330
rect 103643 657000 162436 657090
rect 103643 656760 110810 657000
rect 111050 656760 111160 657000
rect 111400 656760 111490 657000
rect 111730 656760 111820 657000
rect 112060 656760 112150 657000
rect 112390 656760 112500 657000
rect 112740 656760 112830 657000
rect 113070 656760 113160 657000
rect 113400 656760 113490 657000
rect 113730 656760 113840 657000
rect 114080 656760 114170 657000
rect 114410 656760 114500 657000
rect 114740 656760 114830 657000
rect 115070 656760 115180 657000
rect 115420 656760 115510 657000
rect 115750 656760 115840 657000
rect 116080 656760 116170 657000
rect 116410 656760 116520 657000
rect 116760 656760 116850 657000
rect 117090 656760 117180 657000
rect 117420 656760 117510 657000
rect 117750 656760 117860 657000
rect 118100 656760 118190 657000
rect 118430 656760 118520 657000
rect 118760 656760 118850 657000
rect 119090 656760 119200 657000
rect 119440 656760 119530 657000
rect 119770 656760 119860 657000
rect 120100 656760 120190 657000
rect 120430 656760 120540 657000
rect 120780 656760 120870 657000
rect 121110 656760 121200 657000
rect 121440 656760 121530 657000
rect 121770 656760 122190 657000
rect 122430 656760 122540 657000
rect 122780 656760 122870 657000
rect 123110 656760 123200 657000
rect 123440 656760 123530 657000
rect 123770 656760 123880 657000
rect 124120 656760 124210 657000
rect 124450 656760 124540 657000
rect 124780 656760 124870 657000
rect 125110 656760 125220 657000
rect 125460 656760 125550 657000
rect 125790 656760 125880 657000
rect 126120 656760 126210 657000
rect 126450 656760 126560 657000
rect 126800 656760 126890 657000
rect 127130 656760 127220 657000
rect 127460 656760 127550 657000
rect 127790 656760 127900 657000
rect 128140 656760 128230 657000
rect 128470 656760 128560 657000
rect 128800 656760 128890 657000
rect 129130 656760 129240 657000
rect 129480 656760 129570 657000
rect 129810 656760 129900 657000
rect 130140 656760 130230 657000
rect 130470 656760 130580 657000
rect 130820 656760 130910 657000
rect 131150 656760 131240 657000
rect 131480 656760 131570 657000
rect 131810 656760 131920 657000
rect 132160 656760 132250 657000
rect 132490 656760 132580 657000
rect 132820 656760 132910 657000
rect 133150 656760 133570 657000
rect 133810 656760 133920 657000
rect 134160 656760 134250 657000
rect 134490 656760 134580 657000
rect 134820 656760 134910 657000
rect 135150 656760 135260 657000
rect 135500 656760 135590 657000
rect 135830 656760 135920 657000
rect 136160 656760 136250 657000
rect 136490 656760 136600 657000
rect 136840 656760 136930 657000
rect 137170 656760 137260 657000
rect 137500 656760 137590 657000
rect 137830 656760 137940 657000
rect 138180 656760 138270 657000
rect 138510 656760 138600 657000
rect 138840 656760 138930 657000
rect 139170 656760 139280 657000
rect 139520 656760 139610 657000
rect 139850 656760 139940 657000
rect 140180 656760 140270 657000
rect 140510 656760 140620 657000
rect 140860 656760 140950 657000
rect 141190 656760 141280 657000
rect 141520 656760 141610 657000
rect 141850 656760 141960 657000
rect 142200 656760 142290 657000
rect 142530 656760 142620 657000
rect 142860 656760 142950 657000
rect 143190 656760 143300 657000
rect 143540 656760 143630 657000
rect 143870 656760 143960 657000
rect 144200 656760 144290 657000
rect 144530 656760 144950 657000
rect 145190 656760 145300 657000
rect 145540 656760 145630 657000
rect 145870 656760 145960 657000
rect 146200 656760 146290 657000
rect 146530 656760 146640 657000
rect 146880 656760 146970 657000
rect 147210 656760 147300 657000
rect 147540 656760 147630 657000
rect 147870 656760 147980 657000
rect 148220 656760 148310 657000
rect 148550 656760 148640 657000
rect 148880 656760 148970 657000
rect 149210 656760 149320 657000
rect 149560 656760 149650 657000
rect 149890 656760 149980 657000
rect 150220 656760 150310 657000
rect 150550 656760 150660 657000
rect 150900 656760 150990 657000
rect 151230 656760 151320 657000
rect 151560 656760 151650 657000
rect 151890 656760 152000 657000
rect 152240 656760 152330 657000
rect 152570 656760 152660 657000
rect 152900 656760 152990 657000
rect 153230 656760 153340 657000
rect 153580 656760 153670 657000
rect 153910 656760 154000 657000
rect 154240 656760 154330 657000
rect 154570 656760 154680 657000
rect 154920 656760 155010 657000
rect 155250 656760 155340 657000
rect 155580 656760 155670 657000
rect 155910 656760 162436 657000
rect 103643 656670 162436 656760
rect 103643 656430 110810 656670
rect 111050 656430 111160 656670
rect 111400 656430 111490 656670
rect 111730 656430 111820 656670
rect 112060 656430 112150 656670
rect 112390 656430 112500 656670
rect 112740 656430 112830 656670
rect 113070 656430 113160 656670
rect 113400 656430 113490 656670
rect 113730 656430 113840 656670
rect 114080 656430 114170 656670
rect 114410 656430 114500 656670
rect 114740 656430 114830 656670
rect 115070 656430 115180 656670
rect 115420 656430 115510 656670
rect 115750 656430 115840 656670
rect 116080 656430 116170 656670
rect 116410 656430 116520 656670
rect 116760 656430 116850 656670
rect 117090 656430 117180 656670
rect 117420 656430 117510 656670
rect 117750 656430 117860 656670
rect 118100 656430 118190 656670
rect 118430 656430 118520 656670
rect 118760 656430 118850 656670
rect 119090 656430 119200 656670
rect 119440 656430 119530 656670
rect 119770 656430 119860 656670
rect 120100 656430 120190 656670
rect 120430 656430 120540 656670
rect 120780 656430 120870 656670
rect 121110 656430 121200 656670
rect 121440 656430 121530 656670
rect 121770 656430 122190 656670
rect 122430 656430 122540 656670
rect 122780 656430 122870 656670
rect 123110 656430 123200 656670
rect 123440 656430 123530 656670
rect 123770 656430 123880 656670
rect 124120 656430 124210 656670
rect 124450 656430 124540 656670
rect 124780 656430 124870 656670
rect 125110 656430 125220 656670
rect 125460 656430 125550 656670
rect 125790 656430 125880 656670
rect 126120 656430 126210 656670
rect 126450 656430 126560 656670
rect 126800 656430 126890 656670
rect 127130 656430 127220 656670
rect 127460 656430 127550 656670
rect 127790 656430 127900 656670
rect 128140 656430 128230 656670
rect 128470 656430 128560 656670
rect 128800 656430 128890 656670
rect 129130 656430 129240 656670
rect 129480 656430 129570 656670
rect 129810 656430 129900 656670
rect 130140 656430 130230 656670
rect 130470 656430 130580 656670
rect 130820 656430 130910 656670
rect 131150 656430 131240 656670
rect 131480 656430 131570 656670
rect 131810 656430 131920 656670
rect 132160 656430 132250 656670
rect 132490 656430 132580 656670
rect 132820 656430 132910 656670
rect 133150 656430 133570 656670
rect 133810 656430 133920 656670
rect 134160 656430 134250 656670
rect 134490 656430 134580 656670
rect 134820 656430 134910 656670
rect 135150 656430 135260 656670
rect 135500 656430 135590 656670
rect 135830 656430 135920 656670
rect 136160 656430 136250 656670
rect 136490 656430 136600 656670
rect 136840 656430 136930 656670
rect 137170 656430 137260 656670
rect 137500 656430 137590 656670
rect 137830 656430 137940 656670
rect 138180 656430 138270 656670
rect 138510 656430 138600 656670
rect 138840 656430 138930 656670
rect 139170 656430 139280 656670
rect 139520 656430 139610 656670
rect 139850 656430 139940 656670
rect 140180 656430 140270 656670
rect 140510 656430 140620 656670
rect 140860 656430 140950 656670
rect 141190 656430 141280 656670
rect 141520 656430 141610 656670
rect 141850 656430 141960 656670
rect 142200 656430 142290 656670
rect 142530 656430 142620 656670
rect 142860 656430 142950 656670
rect 143190 656430 143300 656670
rect 143540 656430 143630 656670
rect 143870 656430 143960 656670
rect 144200 656430 144290 656670
rect 144530 656430 144950 656670
rect 145190 656430 145300 656670
rect 145540 656430 145630 656670
rect 145870 656430 145960 656670
rect 146200 656430 146290 656670
rect 146530 656430 146640 656670
rect 146880 656430 146970 656670
rect 147210 656430 147300 656670
rect 147540 656430 147630 656670
rect 147870 656430 147980 656670
rect 148220 656430 148310 656670
rect 148550 656430 148640 656670
rect 148880 656430 148970 656670
rect 149210 656430 149320 656670
rect 149560 656430 149650 656670
rect 149890 656430 149980 656670
rect 150220 656430 150310 656670
rect 150550 656430 150660 656670
rect 150900 656430 150990 656670
rect 151230 656430 151320 656670
rect 151560 656430 151650 656670
rect 151890 656430 152000 656670
rect 152240 656430 152330 656670
rect 152570 656430 152660 656670
rect 152900 656430 152990 656670
rect 153230 656430 153340 656670
rect 153580 656430 153670 656670
rect 153910 656430 154000 656670
rect 154240 656430 154330 656670
rect 154570 656430 154680 656670
rect 154920 656430 155010 656670
rect 155250 656430 155340 656670
rect 155580 656430 155670 656670
rect 155910 656430 162436 656670
rect 103643 656320 162436 656430
rect 103643 656080 110810 656320
rect 111050 656080 111160 656320
rect 111400 656080 111490 656320
rect 111730 656080 111820 656320
rect 112060 656080 112150 656320
rect 112390 656080 112500 656320
rect 112740 656080 112830 656320
rect 113070 656080 113160 656320
rect 113400 656080 113490 656320
rect 113730 656080 113840 656320
rect 114080 656080 114170 656320
rect 114410 656080 114500 656320
rect 114740 656080 114830 656320
rect 115070 656080 115180 656320
rect 115420 656080 115510 656320
rect 115750 656080 115840 656320
rect 116080 656080 116170 656320
rect 116410 656080 116520 656320
rect 116760 656080 116850 656320
rect 117090 656080 117180 656320
rect 117420 656080 117510 656320
rect 117750 656080 117860 656320
rect 118100 656080 118190 656320
rect 118430 656080 118520 656320
rect 118760 656080 118850 656320
rect 119090 656080 119200 656320
rect 119440 656080 119530 656320
rect 119770 656080 119860 656320
rect 120100 656080 120190 656320
rect 120430 656080 120540 656320
rect 120780 656080 120870 656320
rect 121110 656080 121200 656320
rect 121440 656080 121530 656320
rect 121770 656080 122190 656320
rect 122430 656080 122540 656320
rect 122780 656080 122870 656320
rect 123110 656080 123200 656320
rect 123440 656080 123530 656320
rect 123770 656080 123880 656320
rect 124120 656080 124210 656320
rect 124450 656080 124540 656320
rect 124780 656080 124870 656320
rect 125110 656080 125220 656320
rect 125460 656080 125550 656320
rect 125790 656080 125880 656320
rect 126120 656080 126210 656320
rect 126450 656080 126560 656320
rect 126800 656080 126890 656320
rect 127130 656080 127220 656320
rect 127460 656080 127550 656320
rect 127790 656080 127900 656320
rect 128140 656080 128230 656320
rect 128470 656080 128560 656320
rect 128800 656080 128890 656320
rect 129130 656080 129240 656320
rect 129480 656080 129570 656320
rect 129810 656080 129900 656320
rect 130140 656080 130230 656320
rect 130470 656080 130580 656320
rect 130820 656080 130910 656320
rect 131150 656080 131240 656320
rect 131480 656080 131570 656320
rect 131810 656080 131920 656320
rect 132160 656080 132250 656320
rect 132490 656080 132580 656320
rect 132820 656080 132910 656320
rect 133150 656080 133570 656320
rect 133810 656080 133920 656320
rect 134160 656080 134250 656320
rect 134490 656080 134580 656320
rect 134820 656080 134910 656320
rect 135150 656080 135260 656320
rect 135500 656080 135590 656320
rect 135830 656080 135920 656320
rect 136160 656080 136250 656320
rect 136490 656080 136600 656320
rect 136840 656080 136930 656320
rect 137170 656080 137260 656320
rect 137500 656080 137590 656320
rect 137830 656080 137940 656320
rect 138180 656080 138270 656320
rect 138510 656080 138600 656320
rect 138840 656080 138930 656320
rect 139170 656080 139280 656320
rect 139520 656080 139610 656320
rect 139850 656080 139940 656320
rect 140180 656080 140270 656320
rect 140510 656080 140620 656320
rect 140860 656080 140950 656320
rect 141190 656080 141280 656320
rect 141520 656080 141610 656320
rect 141850 656080 141960 656320
rect 142200 656080 142290 656320
rect 142530 656080 142620 656320
rect 142860 656080 142950 656320
rect 143190 656080 143300 656320
rect 143540 656080 143630 656320
rect 143870 656080 143960 656320
rect 144200 656080 144290 656320
rect 144530 656080 144950 656320
rect 145190 656080 145300 656320
rect 145540 656080 145630 656320
rect 145870 656080 145960 656320
rect 146200 656080 146290 656320
rect 146530 656080 146640 656320
rect 146880 656080 146970 656320
rect 147210 656080 147300 656320
rect 147540 656080 147630 656320
rect 147870 656080 147980 656320
rect 148220 656080 148310 656320
rect 148550 656080 148640 656320
rect 148880 656080 148970 656320
rect 149210 656080 149320 656320
rect 149560 656080 149650 656320
rect 149890 656080 149980 656320
rect 150220 656080 150310 656320
rect 150550 656080 150660 656320
rect 150900 656080 150990 656320
rect 151230 656080 151320 656320
rect 151560 656080 151650 656320
rect 151890 656080 152000 656320
rect 152240 656080 152330 656320
rect 152570 656080 152660 656320
rect 152900 656080 152990 656320
rect 153230 656080 153340 656320
rect 153580 656080 153670 656320
rect 153910 656080 154000 656320
rect 154240 656080 154330 656320
rect 154570 656080 154680 656320
rect 154920 656080 155010 656320
rect 155250 656080 155340 656320
rect 155580 656080 155670 656320
rect 155910 656080 162436 656320
rect 103643 655990 162436 656080
rect 103643 655750 110810 655990
rect 111050 655750 111160 655990
rect 111400 655750 111490 655990
rect 111730 655750 111820 655990
rect 112060 655750 112150 655990
rect 112390 655750 112500 655990
rect 112740 655750 112830 655990
rect 113070 655750 113160 655990
rect 113400 655750 113490 655990
rect 113730 655750 113840 655990
rect 114080 655750 114170 655990
rect 114410 655750 114500 655990
rect 114740 655750 114830 655990
rect 115070 655750 115180 655990
rect 115420 655750 115510 655990
rect 115750 655750 115840 655990
rect 116080 655750 116170 655990
rect 116410 655750 116520 655990
rect 116760 655750 116850 655990
rect 117090 655750 117180 655990
rect 117420 655750 117510 655990
rect 117750 655750 117860 655990
rect 118100 655750 118190 655990
rect 118430 655750 118520 655990
rect 118760 655750 118850 655990
rect 119090 655750 119200 655990
rect 119440 655750 119530 655990
rect 119770 655750 119860 655990
rect 120100 655750 120190 655990
rect 120430 655750 120540 655990
rect 120780 655750 120870 655990
rect 121110 655750 121200 655990
rect 121440 655750 121530 655990
rect 121770 655750 122190 655990
rect 122430 655750 122540 655990
rect 122780 655750 122870 655990
rect 123110 655750 123200 655990
rect 123440 655750 123530 655990
rect 123770 655750 123880 655990
rect 124120 655750 124210 655990
rect 124450 655750 124540 655990
rect 124780 655750 124870 655990
rect 125110 655750 125220 655990
rect 125460 655750 125550 655990
rect 125790 655750 125880 655990
rect 126120 655750 126210 655990
rect 126450 655750 126560 655990
rect 126800 655750 126890 655990
rect 127130 655750 127220 655990
rect 127460 655750 127550 655990
rect 127790 655750 127900 655990
rect 128140 655750 128230 655990
rect 128470 655750 128560 655990
rect 128800 655750 128890 655990
rect 129130 655750 129240 655990
rect 129480 655750 129570 655990
rect 129810 655750 129900 655990
rect 130140 655750 130230 655990
rect 130470 655750 130580 655990
rect 130820 655750 130910 655990
rect 131150 655750 131240 655990
rect 131480 655750 131570 655990
rect 131810 655750 131920 655990
rect 132160 655750 132250 655990
rect 132490 655750 132580 655990
rect 132820 655750 132910 655990
rect 133150 655750 133570 655990
rect 133810 655750 133920 655990
rect 134160 655750 134250 655990
rect 134490 655750 134580 655990
rect 134820 655750 134910 655990
rect 135150 655750 135260 655990
rect 135500 655750 135590 655990
rect 135830 655750 135920 655990
rect 136160 655750 136250 655990
rect 136490 655750 136600 655990
rect 136840 655750 136930 655990
rect 137170 655750 137260 655990
rect 137500 655750 137590 655990
rect 137830 655750 137940 655990
rect 138180 655750 138270 655990
rect 138510 655750 138600 655990
rect 138840 655750 138930 655990
rect 139170 655750 139280 655990
rect 139520 655750 139610 655990
rect 139850 655750 139940 655990
rect 140180 655750 140270 655990
rect 140510 655750 140620 655990
rect 140860 655750 140950 655990
rect 141190 655750 141280 655990
rect 141520 655750 141610 655990
rect 141850 655750 141960 655990
rect 142200 655750 142290 655990
rect 142530 655750 142620 655990
rect 142860 655750 142950 655990
rect 143190 655750 143300 655990
rect 143540 655750 143630 655990
rect 143870 655750 143960 655990
rect 144200 655750 144290 655990
rect 144530 655750 144950 655990
rect 145190 655750 145300 655990
rect 145540 655750 145630 655990
rect 145870 655750 145960 655990
rect 146200 655750 146290 655990
rect 146530 655750 146640 655990
rect 146880 655750 146970 655990
rect 147210 655750 147300 655990
rect 147540 655750 147630 655990
rect 147870 655750 147980 655990
rect 148220 655750 148310 655990
rect 148550 655750 148640 655990
rect 148880 655750 148970 655990
rect 149210 655750 149320 655990
rect 149560 655750 149650 655990
rect 149890 655750 149980 655990
rect 150220 655750 150310 655990
rect 150550 655750 150660 655990
rect 150900 655750 150990 655990
rect 151230 655750 151320 655990
rect 151560 655750 151650 655990
rect 151890 655750 152000 655990
rect 152240 655750 152330 655990
rect 152570 655750 152660 655990
rect 152900 655750 152990 655990
rect 153230 655750 153340 655990
rect 153580 655750 153670 655990
rect 153910 655750 154000 655990
rect 154240 655750 154330 655990
rect 154570 655750 154680 655990
rect 154920 655750 155010 655990
rect 155250 655750 155340 655990
rect 155580 655750 155670 655990
rect 155910 655750 162436 655990
rect 103643 655660 162436 655750
rect 103643 655420 110810 655660
rect 111050 655420 111160 655660
rect 111400 655420 111490 655660
rect 111730 655420 111820 655660
rect 112060 655420 112150 655660
rect 112390 655420 112500 655660
rect 112740 655420 112830 655660
rect 113070 655420 113160 655660
rect 113400 655420 113490 655660
rect 113730 655420 113840 655660
rect 114080 655420 114170 655660
rect 114410 655420 114500 655660
rect 114740 655420 114830 655660
rect 115070 655420 115180 655660
rect 115420 655420 115510 655660
rect 115750 655420 115840 655660
rect 116080 655420 116170 655660
rect 116410 655420 116520 655660
rect 116760 655420 116850 655660
rect 117090 655420 117180 655660
rect 117420 655420 117510 655660
rect 117750 655420 117860 655660
rect 118100 655420 118190 655660
rect 118430 655420 118520 655660
rect 118760 655420 118850 655660
rect 119090 655420 119200 655660
rect 119440 655420 119530 655660
rect 119770 655420 119860 655660
rect 120100 655420 120190 655660
rect 120430 655420 120540 655660
rect 120780 655420 120870 655660
rect 121110 655420 121200 655660
rect 121440 655420 121530 655660
rect 121770 655420 122190 655660
rect 122430 655420 122540 655660
rect 122780 655420 122870 655660
rect 123110 655420 123200 655660
rect 123440 655420 123530 655660
rect 123770 655420 123880 655660
rect 124120 655420 124210 655660
rect 124450 655420 124540 655660
rect 124780 655420 124870 655660
rect 125110 655420 125220 655660
rect 125460 655420 125550 655660
rect 125790 655420 125880 655660
rect 126120 655420 126210 655660
rect 126450 655420 126560 655660
rect 126800 655420 126890 655660
rect 127130 655420 127220 655660
rect 127460 655420 127550 655660
rect 127790 655420 127900 655660
rect 128140 655420 128230 655660
rect 128470 655420 128560 655660
rect 128800 655420 128890 655660
rect 129130 655420 129240 655660
rect 129480 655420 129570 655660
rect 129810 655420 129900 655660
rect 130140 655420 130230 655660
rect 130470 655420 130580 655660
rect 130820 655420 130910 655660
rect 131150 655420 131240 655660
rect 131480 655420 131570 655660
rect 131810 655420 131920 655660
rect 132160 655420 132250 655660
rect 132490 655420 132580 655660
rect 132820 655420 132910 655660
rect 133150 655420 133570 655660
rect 133810 655420 133920 655660
rect 134160 655420 134250 655660
rect 134490 655420 134580 655660
rect 134820 655420 134910 655660
rect 135150 655420 135260 655660
rect 135500 655420 135590 655660
rect 135830 655420 135920 655660
rect 136160 655420 136250 655660
rect 136490 655420 136600 655660
rect 136840 655420 136930 655660
rect 137170 655420 137260 655660
rect 137500 655420 137590 655660
rect 137830 655420 137940 655660
rect 138180 655420 138270 655660
rect 138510 655420 138600 655660
rect 138840 655420 138930 655660
rect 139170 655420 139280 655660
rect 139520 655420 139610 655660
rect 139850 655420 139940 655660
rect 140180 655420 140270 655660
rect 140510 655420 140620 655660
rect 140860 655420 140950 655660
rect 141190 655420 141280 655660
rect 141520 655420 141610 655660
rect 141850 655420 141960 655660
rect 142200 655420 142290 655660
rect 142530 655420 142620 655660
rect 142860 655420 142950 655660
rect 143190 655420 143300 655660
rect 143540 655420 143630 655660
rect 143870 655420 143960 655660
rect 144200 655420 144290 655660
rect 144530 655420 144950 655660
rect 145190 655420 145300 655660
rect 145540 655420 145630 655660
rect 145870 655420 145960 655660
rect 146200 655420 146290 655660
rect 146530 655420 146640 655660
rect 146880 655420 146970 655660
rect 147210 655420 147300 655660
rect 147540 655420 147630 655660
rect 147870 655420 147980 655660
rect 148220 655420 148310 655660
rect 148550 655420 148640 655660
rect 148880 655420 148970 655660
rect 149210 655420 149320 655660
rect 149560 655420 149650 655660
rect 149890 655420 149980 655660
rect 150220 655420 150310 655660
rect 150550 655420 150660 655660
rect 150900 655420 150990 655660
rect 151230 655420 151320 655660
rect 151560 655420 151650 655660
rect 151890 655420 152000 655660
rect 152240 655420 152330 655660
rect 152570 655420 152660 655660
rect 152900 655420 152990 655660
rect 153230 655420 153340 655660
rect 153580 655420 153670 655660
rect 153910 655420 154000 655660
rect 154240 655420 154330 655660
rect 154570 655420 154680 655660
rect 154920 655420 155010 655660
rect 155250 655420 155340 655660
rect 155580 655420 155670 655660
rect 155910 655420 162436 655660
rect 103643 655330 162436 655420
rect 103643 655090 110810 655330
rect 111050 655090 111160 655330
rect 111400 655090 111490 655330
rect 111730 655090 111820 655330
rect 112060 655090 112150 655330
rect 112390 655090 112500 655330
rect 112740 655090 112830 655330
rect 113070 655090 113160 655330
rect 113400 655090 113490 655330
rect 113730 655090 113840 655330
rect 114080 655090 114170 655330
rect 114410 655090 114500 655330
rect 114740 655090 114830 655330
rect 115070 655090 115180 655330
rect 115420 655090 115510 655330
rect 115750 655090 115840 655330
rect 116080 655090 116170 655330
rect 116410 655090 116520 655330
rect 116760 655090 116850 655330
rect 117090 655090 117180 655330
rect 117420 655090 117510 655330
rect 117750 655090 117860 655330
rect 118100 655090 118190 655330
rect 118430 655090 118520 655330
rect 118760 655090 118850 655330
rect 119090 655090 119200 655330
rect 119440 655090 119530 655330
rect 119770 655090 119860 655330
rect 120100 655090 120190 655330
rect 120430 655090 120540 655330
rect 120780 655090 120870 655330
rect 121110 655090 121200 655330
rect 121440 655090 121530 655330
rect 121770 655090 122190 655330
rect 122430 655090 122540 655330
rect 122780 655090 122870 655330
rect 123110 655090 123200 655330
rect 123440 655090 123530 655330
rect 123770 655090 123880 655330
rect 124120 655090 124210 655330
rect 124450 655090 124540 655330
rect 124780 655090 124870 655330
rect 125110 655090 125220 655330
rect 125460 655090 125550 655330
rect 125790 655090 125880 655330
rect 126120 655090 126210 655330
rect 126450 655090 126560 655330
rect 126800 655090 126890 655330
rect 127130 655090 127220 655330
rect 127460 655090 127550 655330
rect 127790 655090 127900 655330
rect 128140 655090 128230 655330
rect 128470 655090 128560 655330
rect 128800 655090 128890 655330
rect 129130 655090 129240 655330
rect 129480 655090 129570 655330
rect 129810 655090 129900 655330
rect 130140 655090 130230 655330
rect 130470 655090 130580 655330
rect 130820 655090 130910 655330
rect 131150 655090 131240 655330
rect 131480 655090 131570 655330
rect 131810 655090 131920 655330
rect 132160 655090 132250 655330
rect 132490 655090 132580 655330
rect 132820 655090 132910 655330
rect 133150 655090 133570 655330
rect 133810 655090 133920 655330
rect 134160 655090 134250 655330
rect 134490 655090 134580 655330
rect 134820 655090 134910 655330
rect 135150 655090 135260 655330
rect 135500 655090 135590 655330
rect 135830 655090 135920 655330
rect 136160 655090 136250 655330
rect 136490 655090 136600 655330
rect 136840 655090 136930 655330
rect 137170 655090 137260 655330
rect 137500 655090 137590 655330
rect 137830 655090 137940 655330
rect 138180 655090 138270 655330
rect 138510 655090 138600 655330
rect 138840 655090 138930 655330
rect 139170 655090 139280 655330
rect 139520 655090 139610 655330
rect 139850 655090 139940 655330
rect 140180 655090 140270 655330
rect 140510 655090 140620 655330
rect 140860 655090 140950 655330
rect 141190 655090 141280 655330
rect 141520 655090 141610 655330
rect 141850 655090 141960 655330
rect 142200 655090 142290 655330
rect 142530 655090 142620 655330
rect 142860 655090 142950 655330
rect 143190 655090 143300 655330
rect 143540 655090 143630 655330
rect 143870 655090 143960 655330
rect 144200 655090 144290 655330
rect 144530 655090 144950 655330
rect 145190 655090 145300 655330
rect 145540 655090 145630 655330
rect 145870 655090 145960 655330
rect 146200 655090 146290 655330
rect 146530 655090 146640 655330
rect 146880 655090 146970 655330
rect 147210 655090 147300 655330
rect 147540 655090 147630 655330
rect 147870 655090 147980 655330
rect 148220 655090 148310 655330
rect 148550 655090 148640 655330
rect 148880 655090 148970 655330
rect 149210 655090 149320 655330
rect 149560 655090 149650 655330
rect 149890 655090 149980 655330
rect 150220 655090 150310 655330
rect 150550 655090 150660 655330
rect 150900 655090 150990 655330
rect 151230 655090 151320 655330
rect 151560 655090 151650 655330
rect 151890 655090 152000 655330
rect 152240 655090 152330 655330
rect 152570 655090 152660 655330
rect 152900 655090 152990 655330
rect 153230 655090 153340 655330
rect 153580 655090 153670 655330
rect 153910 655090 154000 655330
rect 154240 655090 154330 655330
rect 154570 655090 154680 655330
rect 154920 655090 155010 655330
rect 155250 655090 155340 655330
rect 155580 655090 155670 655330
rect 155910 655090 162436 655330
rect 103643 654980 162436 655090
rect 569580 654990 569900 702600
rect 103643 654740 110810 654980
rect 111050 654740 111160 654980
rect 111400 654740 111490 654980
rect 111730 654740 111820 654980
rect 112060 654740 112150 654980
rect 112390 654740 112500 654980
rect 112740 654740 112830 654980
rect 113070 654740 113160 654980
rect 113400 654740 113490 654980
rect 113730 654740 113840 654980
rect 114080 654740 114170 654980
rect 114410 654740 114500 654980
rect 114740 654740 114830 654980
rect 115070 654740 115180 654980
rect 115420 654740 115510 654980
rect 115750 654740 115840 654980
rect 116080 654740 116170 654980
rect 116410 654740 116520 654980
rect 116760 654740 116850 654980
rect 117090 654740 117180 654980
rect 117420 654740 117510 654980
rect 117750 654740 117860 654980
rect 118100 654740 118190 654980
rect 118430 654740 118520 654980
rect 118760 654740 118850 654980
rect 119090 654740 119200 654980
rect 119440 654740 119530 654980
rect 119770 654740 119860 654980
rect 120100 654740 120190 654980
rect 120430 654740 120540 654980
rect 120780 654740 120870 654980
rect 121110 654740 121200 654980
rect 121440 654740 121530 654980
rect 121770 654740 122190 654980
rect 122430 654740 122540 654980
rect 122780 654740 122870 654980
rect 123110 654740 123200 654980
rect 123440 654740 123530 654980
rect 123770 654740 123880 654980
rect 124120 654740 124210 654980
rect 124450 654740 124540 654980
rect 124780 654740 124870 654980
rect 125110 654740 125220 654980
rect 125460 654740 125550 654980
rect 125790 654740 125880 654980
rect 126120 654740 126210 654980
rect 126450 654740 126560 654980
rect 126800 654740 126890 654980
rect 127130 654740 127220 654980
rect 127460 654740 127550 654980
rect 127790 654740 127900 654980
rect 128140 654740 128230 654980
rect 128470 654740 128560 654980
rect 128800 654740 128890 654980
rect 129130 654740 129240 654980
rect 129480 654740 129570 654980
rect 129810 654740 129900 654980
rect 130140 654740 130230 654980
rect 130470 654740 130580 654980
rect 130820 654740 130910 654980
rect 131150 654740 131240 654980
rect 131480 654740 131570 654980
rect 131810 654740 131920 654980
rect 132160 654740 132250 654980
rect 132490 654740 132580 654980
rect 132820 654740 132910 654980
rect 133150 654740 133570 654980
rect 133810 654740 133920 654980
rect 134160 654740 134250 654980
rect 134490 654740 134580 654980
rect 134820 654740 134910 654980
rect 135150 654740 135260 654980
rect 135500 654740 135590 654980
rect 135830 654740 135920 654980
rect 136160 654740 136250 654980
rect 136490 654740 136600 654980
rect 136840 654740 136930 654980
rect 137170 654740 137260 654980
rect 137500 654740 137590 654980
rect 137830 654740 137940 654980
rect 138180 654740 138270 654980
rect 138510 654740 138600 654980
rect 138840 654740 138930 654980
rect 139170 654740 139280 654980
rect 139520 654740 139610 654980
rect 139850 654740 139940 654980
rect 140180 654740 140270 654980
rect 140510 654740 140620 654980
rect 140860 654740 140950 654980
rect 141190 654740 141280 654980
rect 141520 654740 141610 654980
rect 141850 654740 141960 654980
rect 142200 654740 142290 654980
rect 142530 654740 142620 654980
rect 142860 654740 142950 654980
rect 143190 654740 143300 654980
rect 143540 654740 143630 654980
rect 143870 654740 143960 654980
rect 144200 654740 144290 654980
rect 144530 654740 144950 654980
rect 145190 654740 145300 654980
rect 145540 654740 145630 654980
rect 145870 654740 145960 654980
rect 146200 654740 146290 654980
rect 146530 654740 146640 654980
rect 146880 654740 146970 654980
rect 147210 654740 147300 654980
rect 147540 654740 147630 654980
rect 147870 654740 147980 654980
rect 148220 654740 148310 654980
rect 148550 654740 148640 654980
rect 148880 654740 148970 654980
rect 149210 654740 149320 654980
rect 149560 654740 149650 654980
rect 149890 654740 149980 654980
rect 150220 654740 150310 654980
rect 150550 654740 150660 654980
rect 150900 654740 150990 654980
rect 151230 654740 151320 654980
rect 151560 654740 151650 654980
rect 151890 654740 152000 654980
rect 152240 654740 152330 654980
rect 152570 654740 152660 654980
rect 152900 654740 152990 654980
rect 153230 654740 153340 654980
rect 153580 654740 153670 654980
rect 153910 654740 154000 654980
rect 154240 654740 154330 654980
rect 154570 654740 154680 654980
rect 154920 654740 155010 654980
rect 155250 654740 155340 654980
rect 155580 654740 155670 654980
rect 155910 654740 162436 654980
rect 103643 654650 162436 654740
rect 222254 654670 569900 654990
rect 576129 679930 583240 679960
rect 576129 679860 582950 679930
rect 583020 679860 583050 679930
rect 583120 679860 583150 679930
rect 583220 679860 583240 679930
rect 576129 679830 583240 679860
rect 576129 679760 582950 679830
rect 583020 679760 583050 679830
rect 583120 679760 583150 679830
rect 583220 679760 583240 679830
rect 576129 679730 583240 679760
rect 576129 679660 582950 679730
rect 583020 679660 583050 679730
rect 583120 679660 583150 679730
rect 583220 679660 583240 679730
rect 576129 679639 583240 679660
rect 103643 654410 110810 654650
rect 111050 654410 111160 654650
rect 111400 654410 111490 654650
rect 111730 654410 111820 654650
rect 112060 654410 112150 654650
rect 112390 654410 112500 654650
rect 112740 654410 112830 654650
rect 113070 654410 113160 654650
rect 113400 654410 113490 654650
rect 113730 654410 113840 654650
rect 114080 654410 114170 654650
rect 114410 654410 114500 654650
rect 114740 654410 114830 654650
rect 115070 654410 115180 654650
rect 115420 654410 115510 654650
rect 115750 654410 115840 654650
rect 116080 654410 116170 654650
rect 116410 654410 116520 654650
rect 116760 654410 116850 654650
rect 117090 654410 117180 654650
rect 117420 654410 117510 654650
rect 117750 654410 117860 654650
rect 118100 654410 118190 654650
rect 118430 654410 118520 654650
rect 118760 654410 118850 654650
rect 119090 654410 119200 654650
rect 119440 654410 119530 654650
rect 119770 654410 119860 654650
rect 120100 654410 120190 654650
rect 120430 654410 120540 654650
rect 120780 654410 120870 654650
rect 121110 654410 121200 654650
rect 121440 654410 121530 654650
rect 121770 654410 122190 654650
rect 122430 654410 122540 654650
rect 122780 654410 122870 654650
rect 123110 654410 123200 654650
rect 123440 654410 123530 654650
rect 123770 654410 123880 654650
rect 124120 654410 124210 654650
rect 124450 654410 124540 654650
rect 124780 654410 124870 654650
rect 125110 654410 125220 654650
rect 125460 654410 125550 654650
rect 125790 654410 125880 654650
rect 126120 654410 126210 654650
rect 126450 654410 126560 654650
rect 126800 654410 126890 654650
rect 127130 654410 127220 654650
rect 127460 654410 127550 654650
rect 127790 654410 127900 654650
rect 128140 654410 128230 654650
rect 128470 654410 128560 654650
rect 128800 654410 128890 654650
rect 129130 654410 129240 654650
rect 129480 654410 129570 654650
rect 129810 654410 129900 654650
rect 130140 654410 130230 654650
rect 130470 654410 130580 654650
rect 130820 654410 130910 654650
rect 131150 654410 131240 654650
rect 131480 654410 131570 654650
rect 131810 654410 131920 654650
rect 132160 654410 132250 654650
rect 132490 654410 132580 654650
rect 132820 654410 132910 654650
rect 133150 654410 133570 654650
rect 133810 654410 133920 654650
rect 134160 654410 134250 654650
rect 134490 654410 134580 654650
rect 134820 654410 134910 654650
rect 135150 654410 135260 654650
rect 135500 654410 135590 654650
rect 135830 654410 135920 654650
rect 136160 654410 136250 654650
rect 136490 654410 136600 654650
rect 136840 654410 136930 654650
rect 137170 654410 137260 654650
rect 137500 654410 137590 654650
rect 137830 654410 137940 654650
rect 138180 654410 138270 654650
rect 138510 654410 138600 654650
rect 138840 654410 138930 654650
rect 139170 654410 139280 654650
rect 139520 654410 139610 654650
rect 139850 654410 139940 654650
rect 140180 654410 140270 654650
rect 140510 654410 140620 654650
rect 140860 654410 140950 654650
rect 141190 654410 141280 654650
rect 141520 654410 141610 654650
rect 141850 654410 141960 654650
rect 142200 654410 142290 654650
rect 142530 654410 142620 654650
rect 142860 654410 142950 654650
rect 143190 654410 143300 654650
rect 143540 654410 143630 654650
rect 143870 654410 143960 654650
rect 144200 654410 144290 654650
rect 144530 654410 144950 654650
rect 145190 654410 145300 654650
rect 145540 654410 145630 654650
rect 145870 654410 145960 654650
rect 146200 654410 146290 654650
rect 146530 654410 146640 654650
rect 146880 654410 146970 654650
rect 147210 654410 147300 654650
rect 147540 654410 147630 654650
rect 147870 654410 147980 654650
rect 148220 654410 148310 654650
rect 148550 654410 148640 654650
rect 148880 654410 148970 654650
rect 149210 654410 149320 654650
rect 149560 654410 149650 654650
rect 149890 654410 149980 654650
rect 150220 654410 150310 654650
rect 150550 654410 150660 654650
rect 150900 654410 150990 654650
rect 151230 654410 151320 654650
rect 151560 654410 151650 654650
rect 151890 654410 152000 654650
rect 152240 654410 152330 654650
rect 152570 654410 152660 654650
rect 152900 654410 152990 654650
rect 153230 654410 153340 654650
rect 153580 654410 153670 654650
rect 153910 654410 154000 654650
rect 154240 654410 154330 654650
rect 154570 654410 154680 654650
rect 154920 654410 155010 654650
rect 155250 654410 155340 654650
rect 155580 654410 155670 654650
rect 155910 654410 162436 654650
rect 103643 654320 162436 654410
rect 103643 654080 110810 654320
rect 111050 654080 111160 654320
rect 111400 654080 111490 654320
rect 111730 654080 111820 654320
rect 112060 654080 112150 654320
rect 112390 654080 112500 654320
rect 112740 654080 112830 654320
rect 113070 654080 113160 654320
rect 113400 654080 113490 654320
rect 113730 654080 113840 654320
rect 114080 654080 114170 654320
rect 114410 654080 114500 654320
rect 114740 654080 114830 654320
rect 115070 654080 115180 654320
rect 115420 654080 115510 654320
rect 115750 654080 115840 654320
rect 116080 654080 116170 654320
rect 116410 654080 116520 654320
rect 116760 654080 116850 654320
rect 117090 654080 117180 654320
rect 117420 654080 117510 654320
rect 117750 654080 117860 654320
rect 118100 654080 118190 654320
rect 118430 654080 118520 654320
rect 118760 654080 118850 654320
rect 119090 654080 119200 654320
rect 119440 654080 119530 654320
rect 119770 654080 119860 654320
rect 120100 654080 120190 654320
rect 120430 654080 120540 654320
rect 120780 654080 120870 654320
rect 121110 654080 121200 654320
rect 121440 654080 121530 654320
rect 121770 654080 122190 654320
rect 122430 654080 122540 654320
rect 122780 654080 122870 654320
rect 123110 654080 123200 654320
rect 123440 654080 123530 654320
rect 123770 654080 123880 654320
rect 124120 654080 124210 654320
rect 124450 654080 124540 654320
rect 124780 654080 124870 654320
rect 125110 654080 125220 654320
rect 125460 654080 125550 654320
rect 125790 654080 125880 654320
rect 126120 654080 126210 654320
rect 126450 654080 126560 654320
rect 126800 654080 126890 654320
rect 127130 654080 127220 654320
rect 127460 654080 127550 654320
rect 127790 654080 127900 654320
rect 128140 654080 128230 654320
rect 128470 654080 128560 654320
rect 128800 654080 128890 654320
rect 129130 654080 129240 654320
rect 129480 654080 129570 654320
rect 129810 654080 129900 654320
rect 130140 654080 130230 654320
rect 130470 654080 130580 654320
rect 130820 654080 130910 654320
rect 131150 654080 131240 654320
rect 131480 654080 131570 654320
rect 131810 654080 131920 654320
rect 132160 654080 132250 654320
rect 132490 654080 132580 654320
rect 132820 654080 132910 654320
rect 133150 654080 133570 654320
rect 133810 654080 133920 654320
rect 134160 654080 134250 654320
rect 134490 654080 134580 654320
rect 134820 654080 134910 654320
rect 135150 654080 135260 654320
rect 135500 654080 135590 654320
rect 135830 654080 135920 654320
rect 136160 654080 136250 654320
rect 136490 654080 136600 654320
rect 136840 654080 136930 654320
rect 137170 654080 137260 654320
rect 137500 654080 137590 654320
rect 137830 654080 137940 654320
rect 138180 654080 138270 654320
rect 138510 654080 138600 654320
rect 138840 654080 138930 654320
rect 139170 654080 139280 654320
rect 139520 654080 139610 654320
rect 139850 654080 139940 654320
rect 140180 654080 140270 654320
rect 140510 654080 140620 654320
rect 140860 654080 140950 654320
rect 141190 654080 141280 654320
rect 141520 654080 141610 654320
rect 141850 654080 141960 654320
rect 142200 654080 142290 654320
rect 142530 654080 142620 654320
rect 142860 654080 142950 654320
rect 143190 654080 143300 654320
rect 143540 654080 143630 654320
rect 143870 654080 143960 654320
rect 144200 654080 144290 654320
rect 144530 654080 144950 654320
rect 145190 654080 145300 654320
rect 145540 654080 145630 654320
rect 145870 654080 145960 654320
rect 146200 654080 146290 654320
rect 146530 654080 146640 654320
rect 146880 654080 146970 654320
rect 147210 654080 147300 654320
rect 147540 654080 147630 654320
rect 147870 654080 147980 654320
rect 148220 654080 148310 654320
rect 148550 654080 148640 654320
rect 148880 654080 148970 654320
rect 149210 654080 149320 654320
rect 149560 654080 149650 654320
rect 149890 654080 149980 654320
rect 150220 654080 150310 654320
rect 150550 654080 150660 654320
rect 150900 654080 150990 654320
rect 151230 654080 151320 654320
rect 151560 654080 151650 654320
rect 151890 654080 152000 654320
rect 152240 654080 152330 654320
rect 152570 654080 152660 654320
rect 152900 654080 152990 654320
rect 153230 654080 153340 654320
rect 153580 654080 153670 654320
rect 153910 654080 154000 654320
rect 154240 654080 154330 654320
rect 154570 654080 154680 654320
rect 154920 654080 155010 654320
rect 155250 654080 155340 654320
rect 155580 654080 155670 654320
rect 155910 654080 162436 654320
rect 103643 653990 162436 654080
rect 103643 653750 110810 653990
rect 111050 653750 111160 653990
rect 111400 653750 111490 653990
rect 111730 653750 111820 653990
rect 112060 653750 112150 653990
rect 112390 653750 112500 653990
rect 112740 653750 112830 653990
rect 113070 653750 113160 653990
rect 113400 653750 113490 653990
rect 113730 653750 113840 653990
rect 114080 653750 114170 653990
rect 114410 653750 114500 653990
rect 114740 653750 114830 653990
rect 115070 653750 115180 653990
rect 115420 653750 115510 653990
rect 115750 653750 115840 653990
rect 116080 653750 116170 653990
rect 116410 653750 116520 653990
rect 116760 653750 116850 653990
rect 117090 653750 117180 653990
rect 117420 653750 117510 653990
rect 117750 653750 117860 653990
rect 118100 653750 118190 653990
rect 118430 653750 118520 653990
rect 118760 653750 118850 653990
rect 119090 653750 119200 653990
rect 119440 653750 119530 653990
rect 119770 653750 119860 653990
rect 120100 653750 120190 653990
rect 120430 653750 120540 653990
rect 120780 653750 120870 653990
rect 121110 653750 121200 653990
rect 121440 653750 121530 653990
rect 121770 653750 122190 653990
rect 122430 653750 122540 653990
rect 122780 653750 122870 653990
rect 123110 653750 123200 653990
rect 123440 653750 123530 653990
rect 123770 653750 123880 653990
rect 124120 653750 124210 653990
rect 124450 653750 124540 653990
rect 124780 653750 124870 653990
rect 125110 653750 125220 653990
rect 125460 653750 125550 653990
rect 125790 653750 125880 653990
rect 126120 653750 126210 653990
rect 126450 653750 126560 653990
rect 126800 653750 126890 653990
rect 127130 653750 127220 653990
rect 127460 653750 127550 653990
rect 127790 653750 127900 653990
rect 128140 653750 128230 653990
rect 128470 653750 128560 653990
rect 128800 653750 128890 653990
rect 129130 653750 129240 653990
rect 129480 653750 129570 653990
rect 129810 653750 129900 653990
rect 130140 653750 130230 653990
rect 130470 653750 130580 653990
rect 130820 653750 130910 653990
rect 131150 653750 131240 653990
rect 131480 653750 131570 653990
rect 131810 653750 131920 653990
rect 132160 653750 132250 653990
rect 132490 653750 132580 653990
rect 132820 653750 132910 653990
rect 133150 653750 133570 653990
rect 133810 653750 133920 653990
rect 134160 653750 134250 653990
rect 134490 653750 134580 653990
rect 134820 653750 134910 653990
rect 135150 653750 135260 653990
rect 135500 653750 135590 653990
rect 135830 653750 135920 653990
rect 136160 653750 136250 653990
rect 136490 653750 136600 653990
rect 136840 653750 136930 653990
rect 137170 653750 137260 653990
rect 137500 653750 137590 653990
rect 137830 653750 137940 653990
rect 138180 653750 138270 653990
rect 138510 653750 138600 653990
rect 138840 653750 138930 653990
rect 139170 653750 139280 653990
rect 139520 653750 139610 653990
rect 139850 653750 139940 653990
rect 140180 653750 140270 653990
rect 140510 653750 140620 653990
rect 140860 653750 140950 653990
rect 141190 653750 141280 653990
rect 141520 653750 141610 653990
rect 141850 653750 141960 653990
rect 142200 653750 142290 653990
rect 142530 653750 142620 653990
rect 142860 653750 142950 653990
rect 143190 653750 143300 653990
rect 143540 653750 143630 653990
rect 143870 653750 143960 653990
rect 144200 653750 144290 653990
rect 144530 653750 144950 653990
rect 145190 653750 145300 653990
rect 145540 653750 145630 653990
rect 145870 653750 145960 653990
rect 146200 653750 146290 653990
rect 146530 653750 146640 653990
rect 146880 653750 146970 653990
rect 147210 653750 147300 653990
rect 147540 653750 147630 653990
rect 147870 653750 147980 653990
rect 148220 653750 148310 653990
rect 148550 653750 148640 653990
rect 148880 653750 148970 653990
rect 149210 653750 149320 653990
rect 149560 653750 149650 653990
rect 149890 653750 149980 653990
rect 150220 653750 150310 653990
rect 150550 653750 150660 653990
rect 150900 653750 150990 653990
rect 151230 653750 151320 653990
rect 151560 653750 151650 653990
rect 151890 653750 152000 653990
rect 152240 653750 152330 653990
rect 152570 653750 152660 653990
rect 152900 653750 152990 653990
rect 153230 653750 153340 653990
rect 153580 653750 153670 653990
rect 153910 653750 154000 653990
rect 154240 653750 154330 653990
rect 154570 653750 154680 653990
rect 154920 653750 155010 653990
rect 155250 653750 155340 653990
rect 155580 653750 155670 653990
rect 155910 653750 162436 653990
rect 103643 653640 162436 653750
rect 103643 653400 110810 653640
rect 111050 653400 111160 653640
rect 111400 653400 111490 653640
rect 111730 653400 111820 653640
rect 112060 653400 112150 653640
rect 112390 653400 112500 653640
rect 112740 653400 112830 653640
rect 113070 653400 113160 653640
rect 113400 653400 113490 653640
rect 113730 653400 113840 653640
rect 114080 653400 114170 653640
rect 114410 653400 114500 653640
rect 114740 653400 114830 653640
rect 115070 653400 115180 653640
rect 115420 653400 115510 653640
rect 115750 653400 115840 653640
rect 116080 653400 116170 653640
rect 116410 653400 116520 653640
rect 116760 653400 116850 653640
rect 117090 653400 117180 653640
rect 117420 653400 117510 653640
rect 117750 653400 117860 653640
rect 118100 653400 118190 653640
rect 118430 653400 118520 653640
rect 118760 653400 118850 653640
rect 119090 653400 119200 653640
rect 119440 653400 119530 653640
rect 119770 653400 119860 653640
rect 120100 653400 120190 653640
rect 120430 653400 120540 653640
rect 120780 653400 120870 653640
rect 121110 653400 121200 653640
rect 121440 653400 121530 653640
rect 121770 653400 122190 653640
rect 122430 653400 122540 653640
rect 122780 653400 122870 653640
rect 123110 653400 123200 653640
rect 123440 653400 123530 653640
rect 123770 653400 123880 653640
rect 124120 653400 124210 653640
rect 124450 653400 124540 653640
rect 124780 653400 124870 653640
rect 125110 653400 125220 653640
rect 125460 653400 125550 653640
rect 125790 653400 125880 653640
rect 126120 653400 126210 653640
rect 126450 653400 126560 653640
rect 126800 653400 126890 653640
rect 127130 653400 127220 653640
rect 127460 653400 127550 653640
rect 127790 653400 127900 653640
rect 128140 653400 128230 653640
rect 128470 653400 128560 653640
rect 128800 653400 128890 653640
rect 129130 653400 129240 653640
rect 129480 653400 129570 653640
rect 129810 653400 129900 653640
rect 130140 653400 130230 653640
rect 130470 653400 130580 653640
rect 130820 653400 130910 653640
rect 131150 653400 131240 653640
rect 131480 653400 131570 653640
rect 131810 653400 131920 653640
rect 132160 653400 132250 653640
rect 132490 653400 132580 653640
rect 132820 653400 132910 653640
rect 133150 653400 133570 653640
rect 133810 653400 133920 653640
rect 134160 653400 134250 653640
rect 134490 653400 134580 653640
rect 134820 653400 134910 653640
rect 135150 653400 135260 653640
rect 135500 653400 135590 653640
rect 135830 653400 135920 653640
rect 136160 653400 136250 653640
rect 136490 653400 136600 653640
rect 136840 653400 136930 653640
rect 137170 653400 137260 653640
rect 137500 653400 137590 653640
rect 137830 653400 137940 653640
rect 138180 653400 138270 653640
rect 138510 653400 138600 653640
rect 138840 653400 138930 653640
rect 139170 653400 139280 653640
rect 139520 653400 139610 653640
rect 139850 653400 139940 653640
rect 140180 653400 140270 653640
rect 140510 653400 140620 653640
rect 140860 653400 140950 653640
rect 141190 653400 141280 653640
rect 141520 653400 141610 653640
rect 141850 653400 141960 653640
rect 142200 653400 142290 653640
rect 142530 653400 142620 653640
rect 142860 653400 142950 653640
rect 143190 653400 143300 653640
rect 143540 653400 143630 653640
rect 143870 653400 143960 653640
rect 144200 653400 144290 653640
rect 144530 653400 144950 653640
rect 145190 653400 145300 653640
rect 145540 653400 145630 653640
rect 145870 653400 145960 653640
rect 146200 653400 146290 653640
rect 146530 653400 146640 653640
rect 146880 653400 146970 653640
rect 147210 653400 147300 653640
rect 147540 653400 147630 653640
rect 147870 653400 147980 653640
rect 148220 653400 148310 653640
rect 148550 653400 148640 653640
rect 148880 653400 148970 653640
rect 149210 653400 149320 653640
rect 149560 653400 149650 653640
rect 149890 653400 149980 653640
rect 150220 653400 150310 653640
rect 150550 653400 150660 653640
rect 150900 653400 150990 653640
rect 151230 653400 151320 653640
rect 151560 653400 151650 653640
rect 151890 653400 152000 653640
rect 152240 653400 152330 653640
rect 152570 653400 152660 653640
rect 152900 653400 152990 653640
rect 153230 653400 153340 653640
rect 153580 653400 153670 653640
rect 153910 653400 154000 653640
rect 154240 653400 154330 653640
rect 154570 653400 154680 653640
rect 154920 653400 155010 653640
rect 155250 653400 155340 653640
rect 155580 653400 155670 653640
rect 155910 653400 162436 653640
rect 103643 653310 162436 653400
rect 103643 653070 110810 653310
rect 111050 653070 111160 653310
rect 111400 653070 111490 653310
rect 111730 653070 111820 653310
rect 112060 653070 112150 653310
rect 112390 653070 112500 653310
rect 112740 653070 112830 653310
rect 113070 653070 113160 653310
rect 113400 653070 113490 653310
rect 113730 653070 113840 653310
rect 114080 653070 114170 653310
rect 114410 653070 114500 653310
rect 114740 653070 114830 653310
rect 115070 653070 115180 653310
rect 115420 653070 115510 653310
rect 115750 653070 115840 653310
rect 116080 653070 116170 653310
rect 116410 653070 116520 653310
rect 116760 653070 116850 653310
rect 117090 653070 117180 653310
rect 117420 653070 117510 653310
rect 117750 653070 117860 653310
rect 118100 653070 118190 653310
rect 118430 653070 118520 653310
rect 118760 653070 118850 653310
rect 119090 653070 119200 653310
rect 119440 653070 119530 653310
rect 119770 653070 119860 653310
rect 120100 653070 120190 653310
rect 120430 653070 120540 653310
rect 120780 653070 120870 653310
rect 121110 653070 121200 653310
rect 121440 653070 121530 653310
rect 121770 653070 122190 653310
rect 122430 653070 122540 653310
rect 122780 653070 122870 653310
rect 123110 653070 123200 653310
rect 123440 653070 123530 653310
rect 123770 653070 123880 653310
rect 124120 653070 124210 653310
rect 124450 653070 124540 653310
rect 124780 653070 124870 653310
rect 125110 653070 125220 653310
rect 125460 653070 125550 653310
rect 125790 653070 125880 653310
rect 126120 653070 126210 653310
rect 126450 653070 126560 653310
rect 126800 653070 126890 653310
rect 127130 653070 127220 653310
rect 127460 653070 127550 653310
rect 127790 653070 127900 653310
rect 128140 653070 128230 653310
rect 128470 653070 128560 653310
rect 128800 653070 128890 653310
rect 129130 653070 129240 653310
rect 129480 653070 129570 653310
rect 129810 653070 129900 653310
rect 130140 653070 130230 653310
rect 130470 653070 130580 653310
rect 130820 653070 130910 653310
rect 131150 653070 131240 653310
rect 131480 653070 131570 653310
rect 131810 653070 131920 653310
rect 132160 653070 132250 653310
rect 132490 653070 132580 653310
rect 132820 653070 132910 653310
rect 133150 653070 133570 653310
rect 133810 653070 133920 653310
rect 134160 653070 134250 653310
rect 134490 653070 134580 653310
rect 134820 653070 134910 653310
rect 135150 653070 135260 653310
rect 135500 653070 135590 653310
rect 135830 653070 135920 653310
rect 136160 653070 136250 653310
rect 136490 653070 136600 653310
rect 136840 653070 136930 653310
rect 137170 653070 137260 653310
rect 137500 653070 137590 653310
rect 137830 653070 137940 653310
rect 138180 653070 138270 653310
rect 138510 653070 138600 653310
rect 138840 653070 138930 653310
rect 139170 653070 139280 653310
rect 139520 653070 139610 653310
rect 139850 653070 139940 653310
rect 140180 653070 140270 653310
rect 140510 653070 140620 653310
rect 140860 653070 140950 653310
rect 141190 653070 141280 653310
rect 141520 653070 141610 653310
rect 141850 653070 141960 653310
rect 142200 653070 142290 653310
rect 142530 653070 142620 653310
rect 142860 653070 142950 653310
rect 143190 653070 143300 653310
rect 143540 653070 143630 653310
rect 143870 653070 143960 653310
rect 144200 653070 144290 653310
rect 144530 653070 144950 653310
rect 145190 653070 145300 653310
rect 145540 653070 145630 653310
rect 145870 653070 145960 653310
rect 146200 653070 146290 653310
rect 146530 653070 146640 653310
rect 146880 653070 146970 653310
rect 147210 653070 147300 653310
rect 147540 653070 147630 653310
rect 147870 653070 147980 653310
rect 148220 653070 148310 653310
rect 148550 653070 148640 653310
rect 148880 653070 148970 653310
rect 149210 653070 149320 653310
rect 149560 653070 149650 653310
rect 149890 653070 149980 653310
rect 150220 653070 150310 653310
rect 150550 653070 150660 653310
rect 150900 653070 150990 653310
rect 151230 653070 151320 653310
rect 151560 653070 151650 653310
rect 151890 653070 152000 653310
rect 152240 653070 152330 653310
rect 152570 653070 152660 653310
rect 152900 653070 152990 653310
rect 153230 653070 153340 653310
rect 153580 653070 153670 653310
rect 153910 653070 154000 653310
rect 154240 653070 154330 653310
rect 154570 653070 154680 653310
rect 154920 653070 155010 653310
rect 155250 653070 155340 653310
rect 155580 653070 155670 653310
rect 155910 653070 162436 653310
rect 103643 652980 162436 653070
rect 103643 652740 110810 652980
rect 111050 652740 111160 652980
rect 111400 652740 111490 652980
rect 111730 652740 111820 652980
rect 112060 652740 112150 652980
rect 112390 652740 112500 652980
rect 112740 652740 112830 652980
rect 113070 652740 113160 652980
rect 113400 652740 113490 652980
rect 113730 652740 113840 652980
rect 114080 652740 114170 652980
rect 114410 652740 114500 652980
rect 114740 652740 114830 652980
rect 115070 652740 115180 652980
rect 115420 652740 115510 652980
rect 115750 652740 115840 652980
rect 116080 652740 116170 652980
rect 116410 652740 116520 652980
rect 116760 652740 116850 652980
rect 117090 652740 117180 652980
rect 117420 652740 117510 652980
rect 117750 652740 117860 652980
rect 118100 652740 118190 652980
rect 118430 652740 118520 652980
rect 118760 652740 118850 652980
rect 119090 652740 119200 652980
rect 119440 652740 119530 652980
rect 119770 652740 119860 652980
rect 120100 652740 120190 652980
rect 120430 652740 120540 652980
rect 120780 652740 120870 652980
rect 121110 652740 121200 652980
rect 121440 652740 121530 652980
rect 121770 652740 122190 652980
rect 122430 652740 122540 652980
rect 122780 652740 122870 652980
rect 123110 652740 123200 652980
rect 123440 652740 123530 652980
rect 123770 652740 123880 652980
rect 124120 652740 124210 652980
rect 124450 652740 124540 652980
rect 124780 652740 124870 652980
rect 125110 652740 125220 652980
rect 125460 652740 125550 652980
rect 125790 652740 125880 652980
rect 126120 652740 126210 652980
rect 126450 652740 126560 652980
rect 126800 652740 126890 652980
rect 127130 652740 127220 652980
rect 127460 652740 127550 652980
rect 127790 652740 127900 652980
rect 128140 652740 128230 652980
rect 128470 652740 128560 652980
rect 128800 652740 128890 652980
rect 129130 652740 129240 652980
rect 129480 652740 129570 652980
rect 129810 652740 129900 652980
rect 130140 652740 130230 652980
rect 130470 652740 130580 652980
rect 130820 652740 130910 652980
rect 131150 652740 131240 652980
rect 131480 652740 131570 652980
rect 131810 652740 131920 652980
rect 132160 652740 132250 652980
rect 132490 652740 132580 652980
rect 132820 652740 132910 652980
rect 133150 652740 133570 652980
rect 133810 652740 133920 652980
rect 134160 652740 134250 652980
rect 134490 652740 134580 652980
rect 134820 652740 134910 652980
rect 135150 652740 135260 652980
rect 135500 652740 135590 652980
rect 135830 652740 135920 652980
rect 136160 652740 136250 652980
rect 136490 652740 136600 652980
rect 136840 652740 136930 652980
rect 137170 652740 137260 652980
rect 137500 652740 137590 652980
rect 137830 652740 137940 652980
rect 138180 652740 138270 652980
rect 138510 652740 138600 652980
rect 138840 652740 138930 652980
rect 139170 652740 139280 652980
rect 139520 652740 139610 652980
rect 139850 652740 139940 652980
rect 140180 652740 140270 652980
rect 140510 652740 140620 652980
rect 140860 652740 140950 652980
rect 141190 652740 141280 652980
rect 141520 652740 141610 652980
rect 141850 652740 141960 652980
rect 142200 652740 142290 652980
rect 142530 652740 142620 652980
rect 142860 652740 142950 652980
rect 143190 652740 143300 652980
rect 143540 652740 143630 652980
rect 143870 652740 143960 652980
rect 144200 652740 144290 652980
rect 144530 652740 144950 652980
rect 145190 652740 145300 652980
rect 145540 652740 145630 652980
rect 145870 652740 145960 652980
rect 146200 652740 146290 652980
rect 146530 652740 146640 652980
rect 146880 652740 146970 652980
rect 147210 652740 147300 652980
rect 147540 652740 147630 652980
rect 147870 652740 147980 652980
rect 148220 652740 148310 652980
rect 148550 652740 148640 652980
rect 148880 652740 148970 652980
rect 149210 652740 149320 652980
rect 149560 652740 149650 652980
rect 149890 652740 149980 652980
rect 150220 652740 150310 652980
rect 150550 652740 150660 652980
rect 150900 652740 150990 652980
rect 151230 652740 151320 652980
rect 151560 652740 151650 652980
rect 151890 652740 152000 652980
rect 152240 652740 152330 652980
rect 152570 652740 152660 652980
rect 152900 652740 152990 652980
rect 153230 652740 153340 652980
rect 153580 652740 153670 652980
rect 153910 652740 154000 652980
rect 154240 652740 154330 652980
rect 154570 652740 154680 652980
rect 154920 652740 155010 652980
rect 155250 652740 155340 652980
rect 155580 652740 155670 652980
rect 155910 652740 162436 652980
rect 103643 652650 162436 652740
rect 103643 652631 110810 652650
rect 110760 652410 110810 652631
rect 111050 652410 111160 652650
rect 111400 652410 111490 652650
rect 111730 652410 111820 652650
rect 112060 652410 112150 652650
rect 112390 652410 112500 652650
rect 112740 652410 112830 652650
rect 113070 652410 113160 652650
rect 113400 652410 113490 652650
rect 113730 652410 113840 652650
rect 114080 652410 114170 652650
rect 114410 652410 114500 652650
rect 114740 652410 114830 652650
rect 115070 652410 115180 652650
rect 115420 652410 115510 652650
rect 115750 652410 115840 652650
rect 116080 652410 116170 652650
rect 116410 652410 116520 652650
rect 116760 652410 116850 652650
rect 117090 652410 117180 652650
rect 117420 652410 117510 652650
rect 117750 652410 117860 652650
rect 118100 652410 118190 652650
rect 118430 652410 118520 652650
rect 118760 652410 118850 652650
rect 119090 652410 119200 652650
rect 119440 652410 119530 652650
rect 119770 652410 119860 652650
rect 120100 652410 120190 652650
rect 120430 652410 120540 652650
rect 120780 652410 120870 652650
rect 121110 652410 121200 652650
rect 121440 652410 121530 652650
rect 121770 652410 122190 652650
rect 122430 652410 122540 652650
rect 122780 652410 122870 652650
rect 123110 652410 123200 652650
rect 123440 652410 123530 652650
rect 123770 652410 123880 652650
rect 124120 652410 124210 652650
rect 124450 652410 124540 652650
rect 124780 652410 124870 652650
rect 125110 652410 125220 652650
rect 125460 652410 125550 652650
rect 125790 652410 125880 652650
rect 126120 652410 126210 652650
rect 126450 652410 126560 652650
rect 126800 652410 126890 652650
rect 127130 652410 127220 652650
rect 127460 652410 127550 652650
rect 127790 652410 127900 652650
rect 128140 652410 128230 652650
rect 128470 652410 128560 652650
rect 128800 652410 128890 652650
rect 129130 652410 129240 652650
rect 129480 652410 129570 652650
rect 129810 652410 129900 652650
rect 130140 652410 130230 652650
rect 130470 652410 130580 652650
rect 130820 652410 130910 652650
rect 131150 652410 131240 652650
rect 131480 652410 131570 652650
rect 131810 652410 131920 652650
rect 132160 652410 132250 652650
rect 132490 652410 132580 652650
rect 132820 652410 132910 652650
rect 133150 652410 133570 652650
rect 133810 652410 133920 652650
rect 134160 652410 134250 652650
rect 134490 652410 134580 652650
rect 134820 652410 134910 652650
rect 135150 652410 135260 652650
rect 135500 652410 135590 652650
rect 135830 652410 135920 652650
rect 136160 652410 136250 652650
rect 136490 652410 136600 652650
rect 136840 652410 136930 652650
rect 137170 652410 137260 652650
rect 137500 652410 137590 652650
rect 137830 652410 137940 652650
rect 138180 652410 138270 652650
rect 138510 652410 138600 652650
rect 138840 652410 138930 652650
rect 139170 652410 139280 652650
rect 139520 652410 139610 652650
rect 139850 652410 139940 652650
rect 140180 652410 140270 652650
rect 140510 652410 140620 652650
rect 140860 652410 140950 652650
rect 141190 652410 141280 652650
rect 141520 652410 141610 652650
rect 141850 652410 141960 652650
rect 142200 652410 142290 652650
rect 142530 652410 142620 652650
rect 142860 652410 142950 652650
rect 143190 652410 143300 652650
rect 143540 652410 143630 652650
rect 143870 652410 143960 652650
rect 144200 652410 144290 652650
rect 144530 652410 144950 652650
rect 145190 652410 145300 652650
rect 145540 652410 145630 652650
rect 145870 652410 145960 652650
rect 146200 652410 146290 652650
rect 146530 652410 146640 652650
rect 146880 652410 146970 652650
rect 147210 652410 147300 652650
rect 147540 652410 147630 652650
rect 147870 652410 147980 652650
rect 148220 652410 148310 652650
rect 148550 652410 148640 652650
rect 148880 652410 148970 652650
rect 149210 652410 149320 652650
rect 149560 652410 149650 652650
rect 149890 652410 149980 652650
rect 150220 652410 150310 652650
rect 150550 652410 150660 652650
rect 150900 652410 150990 652650
rect 151230 652410 151320 652650
rect 151560 652410 151650 652650
rect 151890 652410 152000 652650
rect 152240 652410 152330 652650
rect 152570 652410 152660 652650
rect 152900 652410 152990 652650
rect 153230 652410 153340 652650
rect 153580 652410 153670 652650
rect 153910 652410 154000 652650
rect 154240 652410 154330 652650
rect 154570 652410 154680 652650
rect 154920 652410 155010 652650
rect 155250 652410 155340 652650
rect 155580 652410 155670 652650
rect 155910 652631 162436 652650
rect 155910 652410 155960 652631
rect 110760 652300 155960 652410
rect 110760 652060 110810 652300
rect 111050 652060 111160 652300
rect 111400 652060 111490 652300
rect 111730 652060 111820 652300
rect 112060 652060 112150 652300
rect 112390 652060 112500 652300
rect 112740 652060 112830 652300
rect 113070 652060 113160 652300
rect 113400 652060 113490 652300
rect 113730 652060 113840 652300
rect 114080 652060 114170 652300
rect 114410 652060 114500 652300
rect 114740 652060 114830 652300
rect 115070 652060 115180 652300
rect 115420 652060 115510 652300
rect 115750 652060 115840 652300
rect 116080 652060 116170 652300
rect 116410 652060 116520 652300
rect 116760 652060 116850 652300
rect 117090 652060 117180 652300
rect 117420 652060 117510 652300
rect 117750 652060 117860 652300
rect 118100 652060 118190 652300
rect 118430 652060 118520 652300
rect 118760 652060 118850 652300
rect 119090 652060 119200 652300
rect 119440 652060 119530 652300
rect 119770 652060 119860 652300
rect 120100 652060 120190 652300
rect 120430 652060 120540 652300
rect 120780 652060 120870 652300
rect 121110 652060 121200 652300
rect 121440 652060 121530 652300
rect 121770 652060 122190 652300
rect 122430 652060 122540 652300
rect 122780 652060 122870 652300
rect 123110 652060 123200 652300
rect 123440 652060 123530 652300
rect 123770 652060 123880 652300
rect 124120 652060 124210 652300
rect 124450 652060 124540 652300
rect 124780 652060 124870 652300
rect 125110 652060 125220 652300
rect 125460 652060 125550 652300
rect 125790 652060 125880 652300
rect 126120 652060 126210 652300
rect 126450 652060 126560 652300
rect 126800 652060 126890 652300
rect 127130 652060 127220 652300
rect 127460 652060 127550 652300
rect 127790 652060 127900 652300
rect 128140 652060 128230 652300
rect 128470 652060 128560 652300
rect 128800 652060 128890 652300
rect 129130 652060 129240 652300
rect 129480 652060 129570 652300
rect 129810 652060 129900 652300
rect 130140 652060 130230 652300
rect 130470 652060 130580 652300
rect 130820 652060 130910 652300
rect 131150 652060 131240 652300
rect 131480 652060 131570 652300
rect 131810 652060 131920 652300
rect 132160 652060 132250 652300
rect 132490 652060 132580 652300
rect 132820 652060 132910 652300
rect 133150 652060 133570 652300
rect 133810 652060 133920 652300
rect 134160 652060 134250 652300
rect 134490 652060 134580 652300
rect 134820 652060 134910 652300
rect 135150 652060 135260 652300
rect 135500 652060 135590 652300
rect 135830 652060 135920 652300
rect 136160 652060 136250 652300
rect 136490 652060 136600 652300
rect 136840 652060 136930 652300
rect 137170 652060 137260 652300
rect 137500 652060 137590 652300
rect 137830 652060 137940 652300
rect 138180 652060 138270 652300
rect 138510 652060 138600 652300
rect 138840 652060 138930 652300
rect 139170 652060 139280 652300
rect 139520 652060 139610 652300
rect 139850 652060 139940 652300
rect 140180 652060 140270 652300
rect 140510 652060 140620 652300
rect 140860 652060 140950 652300
rect 141190 652060 141280 652300
rect 141520 652060 141610 652300
rect 141850 652060 141960 652300
rect 142200 652060 142290 652300
rect 142530 652060 142620 652300
rect 142860 652060 142950 652300
rect 143190 652060 143300 652300
rect 143540 652060 143630 652300
rect 143870 652060 143960 652300
rect 144200 652060 144290 652300
rect 144530 652060 144950 652300
rect 145190 652060 145300 652300
rect 145540 652060 145630 652300
rect 145870 652060 145960 652300
rect 146200 652060 146290 652300
rect 146530 652060 146640 652300
rect 146880 652060 146970 652300
rect 147210 652060 147300 652300
rect 147540 652060 147630 652300
rect 147870 652060 147980 652300
rect 148220 652060 148310 652300
rect 148550 652060 148640 652300
rect 148880 652060 148970 652300
rect 149210 652060 149320 652300
rect 149560 652060 149650 652300
rect 149890 652060 149980 652300
rect 150220 652060 150310 652300
rect 150550 652060 150660 652300
rect 150900 652060 150990 652300
rect 151230 652060 151320 652300
rect 151560 652060 151650 652300
rect 151890 652060 152000 652300
rect 152240 652060 152330 652300
rect 152570 652060 152660 652300
rect 152900 652060 152990 652300
rect 153230 652060 153340 652300
rect 153580 652060 153670 652300
rect 153910 652060 154000 652300
rect 154240 652060 154330 652300
rect 154570 652060 154680 652300
rect 154920 652060 155010 652300
rect 155250 652060 155340 652300
rect 155580 652060 155670 652300
rect 155910 652060 155960 652300
rect 110760 651970 155960 652060
rect 110760 651730 110810 651970
rect 111050 651730 111160 651970
rect 111400 651730 111490 651970
rect 111730 651730 111820 651970
rect 112060 651730 112150 651970
rect 112390 651730 112500 651970
rect 112740 651730 112830 651970
rect 113070 651730 113160 651970
rect 113400 651730 113490 651970
rect 113730 651730 113840 651970
rect 114080 651730 114170 651970
rect 114410 651730 114500 651970
rect 114740 651730 114830 651970
rect 115070 651730 115180 651970
rect 115420 651730 115510 651970
rect 115750 651730 115840 651970
rect 116080 651730 116170 651970
rect 116410 651730 116520 651970
rect 116760 651730 116850 651970
rect 117090 651730 117180 651970
rect 117420 651730 117510 651970
rect 117750 651730 117860 651970
rect 118100 651730 118190 651970
rect 118430 651730 118520 651970
rect 118760 651730 118850 651970
rect 119090 651730 119200 651970
rect 119440 651730 119530 651970
rect 119770 651730 119860 651970
rect 120100 651730 120190 651970
rect 120430 651730 120540 651970
rect 120780 651730 120870 651970
rect 121110 651730 121200 651970
rect 121440 651730 121530 651970
rect 121770 651730 122190 651970
rect 122430 651730 122540 651970
rect 122780 651730 122870 651970
rect 123110 651730 123200 651970
rect 123440 651730 123530 651970
rect 123770 651730 123880 651970
rect 124120 651730 124210 651970
rect 124450 651730 124540 651970
rect 124780 651730 124870 651970
rect 125110 651730 125220 651970
rect 125460 651730 125550 651970
rect 125790 651730 125880 651970
rect 126120 651730 126210 651970
rect 126450 651730 126560 651970
rect 126800 651730 126890 651970
rect 127130 651730 127220 651970
rect 127460 651730 127550 651970
rect 127790 651730 127900 651970
rect 128140 651730 128230 651970
rect 128470 651730 128560 651970
rect 128800 651730 128890 651970
rect 129130 651730 129240 651970
rect 129480 651730 129570 651970
rect 129810 651730 129900 651970
rect 130140 651730 130230 651970
rect 130470 651730 130580 651970
rect 130820 651730 130910 651970
rect 131150 651730 131240 651970
rect 131480 651730 131570 651970
rect 131810 651730 131920 651970
rect 132160 651730 132250 651970
rect 132490 651730 132580 651970
rect 132820 651730 132910 651970
rect 133150 651730 133570 651970
rect 133810 651730 133920 651970
rect 134160 651730 134250 651970
rect 134490 651730 134580 651970
rect 134820 651730 134910 651970
rect 135150 651730 135260 651970
rect 135500 651730 135590 651970
rect 135830 651730 135920 651970
rect 136160 651730 136250 651970
rect 136490 651730 136600 651970
rect 136840 651730 136930 651970
rect 137170 651730 137260 651970
rect 137500 651730 137590 651970
rect 137830 651730 137940 651970
rect 138180 651730 138270 651970
rect 138510 651730 138600 651970
rect 138840 651730 138930 651970
rect 139170 651730 139280 651970
rect 139520 651730 139610 651970
rect 139850 651730 139940 651970
rect 140180 651730 140270 651970
rect 140510 651730 140620 651970
rect 140860 651730 140950 651970
rect 141190 651730 141280 651970
rect 141520 651730 141610 651970
rect 141850 651730 141960 651970
rect 142200 651730 142290 651970
rect 142530 651730 142620 651970
rect 142860 651730 142950 651970
rect 143190 651730 143300 651970
rect 143540 651730 143630 651970
rect 143870 651730 143960 651970
rect 144200 651730 144290 651970
rect 144530 651730 144950 651970
rect 145190 651730 145300 651970
rect 145540 651730 145630 651970
rect 145870 651730 145960 651970
rect 146200 651730 146290 651970
rect 146530 651730 146640 651970
rect 146880 651730 146970 651970
rect 147210 651730 147300 651970
rect 147540 651730 147630 651970
rect 147870 651730 147980 651970
rect 148220 651730 148310 651970
rect 148550 651730 148640 651970
rect 148880 651730 148970 651970
rect 149210 651730 149320 651970
rect 149560 651730 149650 651970
rect 149890 651730 149980 651970
rect 150220 651730 150310 651970
rect 150550 651730 150660 651970
rect 150900 651730 150990 651970
rect 151230 651730 151320 651970
rect 151560 651730 151650 651970
rect 151890 651730 152000 651970
rect 152240 651730 152330 651970
rect 152570 651730 152660 651970
rect 152900 651730 152990 651970
rect 153230 651730 153340 651970
rect 153580 651730 153670 651970
rect 153910 651730 154000 651970
rect 154240 651730 154330 651970
rect 154570 651730 154680 651970
rect 154920 651730 155010 651970
rect 155250 651730 155340 651970
rect 155580 651730 155670 651970
rect 155910 651730 155960 651970
rect 110760 651640 155960 651730
rect 110760 651400 110810 651640
rect 111050 651400 111160 651640
rect 111400 651400 111490 651640
rect 111730 651400 111820 651640
rect 112060 651400 112150 651640
rect 112390 651400 112500 651640
rect 112740 651400 112830 651640
rect 113070 651400 113160 651640
rect 113400 651400 113490 651640
rect 113730 651400 113840 651640
rect 114080 651400 114170 651640
rect 114410 651400 114500 651640
rect 114740 651400 114830 651640
rect 115070 651400 115180 651640
rect 115420 651400 115510 651640
rect 115750 651400 115840 651640
rect 116080 651400 116170 651640
rect 116410 651400 116520 651640
rect 116760 651400 116850 651640
rect 117090 651400 117180 651640
rect 117420 651400 117510 651640
rect 117750 651400 117860 651640
rect 118100 651400 118190 651640
rect 118430 651400 118520 651640
rect 118760 651400 118850 651640
rect 119090 651400 119200 651640
rect 119440 651400 119530 651640
rect 119770 651400 119860 651640
rect 120100 651400 120190 651640
rect 120430 651400 120540 651640
rect 120780 651400 120870 651640
rect 121110 651400 121200 651640
rect 121440 651400 121530 651640
rect 121770 651400 122190 651640
rect 122430 651400 122540 651640
rect 122780 651400 122870 651640
rect 123110 651400 123200 651640
rect 123440 651400 123530 651640
rect 123770 651400 123880 651640
rect 124120 651400 124210 651640
rect 124450 651400 124540 651640
rect 124780 651400 124870 651640
rect 125110 651400 125220 651640
rect 125460 651400 125550 651640
rect 125790 651400 125880 651640
rect 126120 651400 126210 651640
rect 126450 651400 126560 651640
rect 126800 651400 126890 651640
rect 127130 651400 127220 651640
rect 127460 651400 127550 651640
rect 127790 651400 127900 651640
rect 128140 651400 128230 651640
rect 128470 651400 128560 651640
rect 128800 651400 128890 651640
rect 129130 651400 129240 651640
rect 129480 651400 129570 651640
rect 129810 651400 129900 651640
rect 130140 651400 130230 651640
rect 130470 651400 130580 651640
rect 130820 651400 130910 651640
rect 131150 651400 131240 651640
rect 131480 651400 131570 651640
rect 131810 651400 131920 651640
rect 132160 651400 132250 651640
rect 132490 651400 132580 651640
rect 132820 651400 132910 651640
rect 133150 651400 133570 651640
rect 133810 651400 133920 651640
rect 134160 651400 134250 651640
rect 134490 651400 134580 651640
rect 134820 651400 134910 651640
rect 135150 651400 135260 651640
rect 135500 651400 135590 651640
rect 135830 651400 135920 651640
rect 136160 651400 136250 651640
rect 136490 651400 136600 651640
rect 136840 651400 136930 651640
rect 137170 651400 137260 651640
rect 137500 651400 137590 651640
rect 137830 651400 137940 651640
rect 138180 651400 138270 651640
rect 138510 651400 138600 651640
rect 138840 651400 138930 651640
rect 139170 651400 139280 651640
rect 139520 651400 139610 651640
rect 139850 651400 139940 651640
rect 140180 651400 140270 651640
rect 140510 651400 140620 651640
rect 140860 651400 140950 651640
rect 141190 651400 141280 651640
rect 141520 651400 141610 651640
rect 141850 651400 141960 651640
rect 142200 651400 142290 651640
rect 142530 651400 142620 651640
rect 142860 651400 142950 651640
rect 143190 651400 143300 651640
rect 143540 651400 143630 651640
rect 143870 651400 143960 651640
rect 144200 651400 144290 651640
rect 144530 651400 144950 651640
rect 145190 651400 145300 651640
rect 145540 651400 145630 651640
rect 145870 651400 145960 651640
rect 146200 651400 146290 651640
rect 146530 651400 146640 651640
rect 146880 651400 146970 651640
rect 147210 651400 147300 651640
rect 147540 651400 147630 651640
rect 147870 651400 147980 651640
rect 148220 651400 148310 651640
rect 148550 651400 148640 651640
rect 148880 651400 148970 651640
rect 149210 651400 149320 651640
rect 149560 651400 149650 651640
rect 149890 651400 149980 651640
rect 150220 651400 150310 651640
rect 150550 651400 150660 651640
rect 150900 651400 150990 651640
rect 151230 651400 151320 651640
rect 151560 651400 151650 651640
rect 151890 651400 152000 651640
rect 152240 651400 152330 651640
rect 152570 651400 152660 651640
rect 152900 651400 152990 651640
rect 153230 651400 153340 651640
rect 153580 651400 153670 651640
rect 153910 651400 154000 651640
rect 154240 651400 154330 651640
rect 154570 651400 154680 651640
rect 154920 651400 155010 651640
rect 155250 651400 155340 651640
rect 155580 651400 155670 651640
rect 155910 651400 155960 651640
rect 110760 651310 155960 651400
rect 110760 651070 110810 651310
rect 111050 651070 111160 651310
rect 111400 651070 111490 651310
rect 111730 651070 111820 651310
rect 112060 651070 112150 651310
rect 112390 651070 112500 651310
rect 112740 651070 112830 651310
rect 113070 651070 113160 651310
rect 113400 651070 113490 651310
rect 113730 651070 113840 651310
rect 114080 651070 114170 651310
rect 114410 651070 114500 651310
rect 114740 651070 114830 651310
rect 115070 651070 115180 651310
rect 115420 651070 115510 651310
rect 115750 651070 115840 651310
rect 116080 651070 116170 651310
rect 116410 651070 116520 651310
rect 116760 651070 116850 651310
rect 117090 651070 117180 651310
rect 117420 651070 117510 651310
rect 117750 651070 117860 651310
rect 118100 651070 118190 651310
rect 118430 651070 118520 651310
rect 118760 651070 118850 651310
rect 119090 651070 119200 651310
rect 119440 651070 119530 651310
rect 119770 651070 119860 651310
rect 120100 651070 120190 651310
rect 120430 651070 120540 651310
rect 120780 651070 120870 651310
rect 121110 651070 121200 651310
rect 121440 651070 121530 651310
rect 121770 651070 122190 651310
rect 122430 651070 122540 651310
rect 122780 651070 122870 651310
rect 123110 651070 123200 651310
rect 123440 651070 123530 651310
rect 123770 651070 123880 651310
rect 124120 651070 124210 651310
rect 124450 651070 124540 651310
rect 124780 651070 124870 651310
rect 125110 651070 125220 651310
rect 125460 651070 125550 651310
rect 125790 651070 125880 651310
rect 126120 651070 126210 651310
rect 126450 651070 126560 651310
rect 126800 651070 126890 651310
rect 127130 651070 127220 651310
rect 127460 651070 127550 651310
rect 127790 651070 127900 651310
rect 128140 651070 128230 651310
rect 128470 651070 128560 651310
rect 128800 651070 128890 651310
rect 129130 651070 129240 651310
rect 129480 651070 129570 651310
rect 129810 651070 129900 651310
rect 130140 651070 130230 651310
rect 130470 651070 130580 651310
rect 130820 651070 130910 651310
rect 131150 651070 131240 651310
rect 131480 651070 131570 651310
rect 131810 651070 131920 651310
rect 132160 651070 132250 651310
rect 132490 651070 132580 651310
rect 132820 651070 132910 651310
rect 133150 651070 133570 651310
rect 133810 651070 133920 651310
rect 134160 651070 134250 651310
rect 134490 651070 134580 651310
rect 134820 651070 134910 651310
rect 135150 651070 135260 651310
rect 135500 651070 135590 651310
rect 135830 651070 135920 651310
rect 136160 651070 136250 651310
rect 136490 651070 136600 651310
rect 136840 651070 136930 651310
rect 137170 651070 137260 651310
rect 137500 651070 137590 651310
rect 137830 651070 137940 651310
rect 138180 651070 138270 651310
rect 138510 651070 138600 651310
rect 138840 651070 138930 651310
rect 139170 651070 139280 651310
rect 139520 651070 139610 651310
rect 139850 651070 139940 651310
rect 140180 651070 140270 651310
rect 140510 651070 140620 651310
rect 140860 651070 140950 651310
rect 141190 651070 141280 651310
rect 141520 651070 141610 651310
rect 141850 651070 141960 651310
rect 142200 651070 142290 651310
rect 142530 651070 142620 651310
rect 142860 651070 142950 651310
rect 143190 651070 143300 651310
rect 143540 651070 143630 651310
rect 143870 651070 143960 651310
rect 144200 651070 144290 651310
rect 144530 651070 144950 651310
rect 145190 651070 145300 651310
rect 145540 651070 145630 651310
rect 145870 651070 145960 651310
rect 146200 651070 146290 651310
rect 146530 651070 146640 651310
rect 146880 651070 146970 651310
rect 147210 651070 147300 651310
rect 147540 651070 147630 651310
rect 147870 651070 147980 651310
rect 148220 651070 148310 651310
rect 148550 651070 148640 651310
rect 148880 651070 148970 651310
rect 149210 651070 149320 651310
rect 149560 651070 149650 651310
rect 149890 651070 149980 651310
rect 150220 651070 150310 651310
rect 150550 651070 150660 651310
rect 150900 651070 150990 651310
rect 151230 651070 151320 651310
rect 151560 651070 151650 651310
rect 151890 651070 152000 651310
rect 152240 651070 152330 651310
rect 152570 651070 152660 651310
rect 152900 651070 152990 651310
rect 153230 651070 153340 651310
rect 153580 651070 153670 651310
rect 153910 651070 154000 651310
rect 154240 651070 154330 651310
rect 154570 651070 154680 651310
rect 154920 651070 155010 651310
rect 155250 651070 155340 651310
rect 155580 651070 155670 651310
rect 155910 651070 155960 651310
rect 110760 650960 155960 651070
rect 110760 650720 110810 650960
rect 111050 650720 111160 650960
rect 111400 650720 111490 650960
rect 111730 650720 111820 650960
rect 112060 650720 112150 650960
rect 112390 650720 112500 650960
rect 112740 650720 112830 650960
rect 113070 650720 113160 650960
rect 113400 650720 113490 650960
rect 113730 650720 113840 650960
rect 114080 650720 114170 650960
rect 114410 650720 114500 650960
rect 114740 650720 114830 650960
rect 115070 650720 115180 650960
rect 115420 650720 115510 650960
rect 115750 650720 115840 650960
rect 116080 650720 116170 650960
rect 116410 650720 116520 650960
rect 116760 650720 116850 650960
rect 117090 650720 117180 650960
rect 117420 650720 117510 650960
rect 117750 650720 117860 650960
rect 118100 650720 118190 650960
rect 118430 650720 118520 650960
rect 118760 650720 118850 650960
rect 119090 650720 119200 650960
rect 119440 650720 119530 650960
rect 119770 650720 119860 650960
rect 120100 650720 120190 650960
rect 120430 650720 120540 650960
rect 120780 650720 120870 650960
rect 121110 650720 121200 650960
rect 121440 650720 121530 650960
rect 121770 650720 122190 650960
rect 122430 650720 122540 650960
rect 122780 650720 122870 650960
rect 123110 650720 123200 650960
rect 123440 650720 123530 650960
rect 123770 650720 123880 650960
rect 124120 650720 124210 650960
rect 124450 650720 124540 650960
rect 124780 650720 124870 650960
rect 125110 650720 125220 650960
rect 125460 650720 125550 650960
rect 125790 650720 125880 650960
rect 126120 650720 126210 650960
rect 126450 650720 126560 650960
rect 126800 650720 126890 650960
rect 127130 650720 127220 650960
rect 127460 650720 127550 650960
rect 127790 650720 127900 650960
rect 128140 650720 128230 650960
rect 128470 650720 128560 650960
rect 128800 650720 128890 650960
rect 129130 650720 129240 650960
rect 129480 650720 129570 650960
rect 129810 650720 129900 650960
rect 130140 650720 130230 650960
rect 130470 650720 130580 650960
rect 130820 650720 130910 650960
rect 131150 650720 131240 650960
rect 131480 650720 131570 650960
rect 131810 650720 131920 650960
rect 132160 650720 132250 650960
rect 132490 650720 132580 650960
rect 132820 650720 132910 650960
rect 133150 650720 133570 650960
rect 133810 650720 133920 650960
rect 134160 650720 134250 650960
rect 134490 650720 134580 650960
rect 134820 650720 134910 650960
rect 135150 650720 135260 650960
rect 135500 650720 135590 650960
rect 135830 650720 135920 650960
rect 136160 650720 136250 650960
rect 136490 650720 136600 650960
rect 136840 650720 136930 650960
rect 137170 650720 137260 650960
rect 137500 650720 137590 650960
rect 137830 650720 137940 650960
rect 138180 650720 138270 650960
rect 138510 650720 138600 650960
rect 138840 650720 138930 650960
rect 139170 650720 139280 650960
rect 139520 650720 139610 650960
rect 139850 650720 139940 650960
rect 140180 650720 140270 650960
rect 140510 650720 140620 650960
rect 140860 650720 140950 650960
rect 141190 650720 141280 650960
rect 141520 650720 141610 650960
rect 141850 650720 141960 650960
rect 142200 650720 142290 650960
rect 142530 650720 142620 650960
rect 142860 650720 142950 650960
rect 143190 650720 143300 650960
rect 143540 650720 143630 650960
rect 143870 650720 143960 650960
rect 144200 650720 144290 650960
rect 144530 650720 144950 650960
rect 145190 650720 145300 650960
rect 145540 650720 145630 650960
rect 145870 650720 145960 650960
rect 146200 650720 146290 650960
rect 146530 650720 146640 650960
rect 146880 650720 146970 650960
rect 147210 650720 147300 650960
rect 147540 650720 147630 650960
rect 147870 650720 147980 650960
rect 148220 650720 148310 650960
rect 148550 650720 148640 650960
rect 148880 650720 148970 650960
rect 149210 650720 149320 650960
rect 149560 650720 149650 650960
rect 149890 650720 149980 650960
rect 150220 650720 150310 650960
rect 150550 650720 150660 650960
rect 150900 650720 150990 650960
rect 151230 650720 151320 650960
rect 151560 650720 151650 650960
rect 151890 650720 152000 650960
rect 152240 650720 152330 650960
rect 152570 650720 152660 650960
rect 152900 650720 152990 650960
rect 153230 650720 153340 650960
rect 153580 650720 153670 650960
rect 153910 650720 154000 650960
rect 154240 650720 154330 650960
rect 154570 650720 154680 650960
rect 154920 650720 155010 650960
rect 155250 650720 155340 650960
rect 155580 650720 155670 650960
rect 155910 650720 155960 650960
rect 110760 650630 155960 650720
rect 110760 650390 110810 650630
rect 111050 650390 111160 650630
rect 111400 650390 111490 650630
rect 111730 650390 111820 650630
rect 112060 650390 112150 650630
rect 112390 650390 112500 650630
rect 112740 650390 112830 650630
rect 113070 650390 113160 650630
rect 113400 650390 113490 650630
rect 113730 650390 113840 650630
rect 114080 650390 114170 650630
rect 114410 650390 114500 650630
rect 114740 650390 114830 650630
rect 115070 650390 115180 650630
rect 115420 650390 115510 650630
rect 115750 650390 115840 650630
rect 116080 650390 116170 650630
rect 116410 650390 116520 650630
rect 116760 650390 116850 650630
rect 117090 650390 117180 650630
rect 117420 650390 117510 650630
rect 117750 650390 117860 650630
rect 118100 650390 118190 650630
rect 118430 650390 118520 650630
rect 118760 650390 118850 650630
rect 119090 650390 119200 650630
rect 119440 650390 119530 650630
rect 119770 650390 119860 650630
rect 120100 650390 120190 650630
rect 120430 650390 120540 650630
rect 120780 650390 120870 650630
rect 121110 650390 121200 650630
rect 121440 650390 121530 650630
rect 121770 650390 122190 650630
rect 122430 650390 122540 650630
rect 122780 650390 122870 650630
rect 123110 650390 123200 650630
rect 123440 650390 123530 650630
rect 123770 650390 123880 650630
rect 124120 650390 124210 650630
rect 124450 650390 124540 650630
rect 124780 650390 124870 650630
rect 125110 650390 125220 650630
rect 125460 650390 125550 650630
rect 125790 650390 125880 650630
rect 126120 650390 126210 650630
rect 126450 650390 126560 650630
rect 126800 650390 126890 650630
rect 127130 650390 127220 650630
rect 127460 650390 127550 650630
rect 127790 650390 127900 650630
rect 128140 650390 128230 650630
rect 128470 650390 128560 650630
rect 128800 650390 128890 650630
rect 129130 650390 129240 650630
rect 129480 650390 129570 650630
rect 129810 650390 129900 650630
rect 130140 650390 130230 650630
rect 130470 650390 130580 650630
rect 130820 650390 130910 650630
rect 131150 650390 131240 650630
rect 131480 650390 131570 650630
rect 131810 650390 131920 650630
rect 132160 650390 132250 650630
rect 132490 650390 132580 650630
rect 132820 650390 132910 650630
rect 133150 650390 133570 650630
rect 133810 650390 133920 650630
rect 134160 650390 134250 650630
rect 134490 650390 134580 650630
rect 134820 650390 134910 650630
rect 135150 650390 135260 650630
rect 135500 650390 135590 650630
rect 135830 650390 135920 650630
rect 136160 650390 136250 650630
rect 136490 650390 136600 650630
rect 136840 650390 136930 650630
rect 137170 650390 137260 650630
rect 137500 650390 137590 650630
rect 137830 650390 137940 650630
rect 138180 650390 138270 650630
rect 138510 650390 138600 650630
rect 138840 650390 138930 650630
rect 139170 650390 139280 650630
rect 139520 650390 139610 650630
rect 139850 650390 139940 650630
rect 140180 650390 140270 650630
rect 140510 650390 140620 650630
rect 140860 650390 140950 650630
rect 141190 650390 141280 650630
rect 141520 650390 141610 650630
rect 141850 650390 141960 650630
rect 142200 650390 142290 650630
rect 142530 650390 142620 650630
rect 142860 650390 142950 650630
rect 143190 650390 143300 650630
rect 143540 650390 143630 650630
rect 143870 650390 143960 650630
rect 144200 650390 144290 650630
rect 144530 650390 144950 650630
rect 145190 650390 145300 650630
rect 145540 650390 145630 650630
rect 145870 650390 145960 650630
rect 146200 650390 146290 650630
rect 146530 650390 146640 650630
rect 146880 650390 146970 650630
rect 147210 650390 147300 650630
rect 147540 650390 147630 650630
rect 147870 650390 147980 650630
rect 148220 650390 148310 650630
rect 148550 650390 148640 650630
rect 148880 650390 148970 650630
rect 149210 650390 149320 650630
rect 149560 650390 149650 650630
rect 149890 650390 149980 650630
rect 150220 650390 150310 650630
rect 150550 650390 150660 650630
rect 150900 650390 150990 650630
rect 151230 650390 151320 650630
rect 151560 650390 151650 650630
rect 151890 650390 152000 650630
rect 152240 650390 152330 650630
rect 152570 650390 152660 650630
rect 152900 650390 152990 650630
rect 153230 650390 153340 650630
rect 153580 650390 153670 650630
rect 153910 650390 154000 650630
rect 154240 650390 154330 650630
rect 154570 650390 154680 650630
rect 154920 650390 155010 650630
rect 155250 650390 155340 650630
rect 155580 650390 155670 650630
rect 155910 650390 155960 650630
rect 110760 650300 155960 650390
rect 110760 650060 110810 650300
rect 111050 650060 111160 650300
rect 111400 650060 111490 650300
rect 111730 650060 111820 650300
rect 112060 650060 112150 650300
rect 112390 650060 112500 650300
rect 112740 650060 112830 650300
rect 113070 650060 113160 650300
rect 113400 650060 113490 650300
rect 113730 650060 113840 650300
rect 114080 650060 114170 650300
rect 114410 650060 114500 650300
rect 114740 650060 114830 650300
rect 115070 650060 115180 650300
rect 115420 650060 115510 650300
rect 115750 650060 115840 650300
rect 116080 650060 116170 650300
rect 116410 650060 116520 650300
rect 116760 650060 116850 650300
rect 117090 650060 117180 650300
rect 117420 650060 117510 650300
rect 117750 650060 117860 650300
rect 118100 650060 118190 650300
rect 118430 650060 118520 650300
rect 118760 650060 118850 650300
rect 119090 650060 119200 650300
rect 119440 650060 119530 650300
rect 119770 650060 119860 650300
rect 120100 650060 120190 650300
rect 120430 650060 120540 650300
rect 120780 650060 120870 650300
rect 121110 650060 121200 650300
rect 121440 650060 121530 650300
rect 121770 650060 122190 650300
rect 122430 650060 122540 650300
rect 122780 650060 122870 650300
rect 123110 650060 123200 650300
rect 123440 650060 123530 650300
rect 123770 650060 123880 650300
rect 124120 650060 124210 650300
rect 124450 650060 124540 650300
rect 124780 650060 124870 650300
rect 125110 650060 125220 650300
rect 125460 650060 125550 650300
rect 125790 650060 125880 650300
rect 126120 650060 126210 650300
rect 126450 650060 126560 650300
rect 126800 650060 126890 650300
rect 127130 650060 127220 650300
rect 127460 650060 127550 650300
rect 127790 650060 127900 650300
rect 128140 650060 128230 650300
rect 128470 650060 128560 650300
rect 128800 650060 128890 650300
rect 129130 650060 129240 650300
rect 129480 650060 129570 650300
rect 129810 650060 129900 650300
rect 130140 650060 130230 650300
rect 130470 650060 130580 650300
rect 130820 650060 130910 650300
rect 131150 650060 131240 650300
rect 131480 650060 131570 650300
rect 131810 650060 131920 650300
rect 132160 650060 132250 650300
rect 132490 650060 132580 650300
rect 132820 650060 132910 650300
rect 133150 650060 133570 650300
rect 133810 650060 133920 650300
rect 134160 650060 134250 650300
rect 134490 650060 134580 650300
rect 134820 650060 134910 650300
rect 135150 650060 135260 650300
rect 135500 650060 135590 650300
rect 135830 650060 135920 650300
rect 136160 650060 136250 650300
rect 136490 650060 136600 650300
rect 136840 650060 136930 650300
rect 137170 650060 137260 650300
rect 137500 650060 137590 650300
rect 137830 650060 137940 650300
rect 138180 650060 138270 650300
rect 138510 650060 138600 650300
rect 138840 650060 138930 650300
rect 139170 650060 139280 650300
rect 139520 650060 139610 650300
rect 139850 650060 139940 650300
rect 140180 650060 140270 650300
rect 140510 650060 140620 650300
rect 140860 650060 140950 650300
rect 141190 650060 141280 650300
rect 141520 650060 141610 650300
rect 141850 650060 141960 650300
rect 142200 650060 142290 650300
rect 142530 650060 142620 650300
rect 142860 650060 142950 650300
rect 143190 650060 143300 650300
rect 143540 650060 143630 650300
rect 143870 650060 143960 650300
rect 144200 650060 144290 650300
rect 144530 650060 144950 650300
rect 145190 650060 145300 650300
rect 145540 650060 145630 650300
rect 145870 650060 145960 650300
rect 146200 650060 146290 650300
rect 146530 650060 146640 650300
rect 146880 650060 146970 650300
rect 147210 650060 147300 650300
rect 147540 650060 147630 650300
rect 147870 650060 147980 650300
rect 148220 650060 148310 650300
rect 148550 650060 148640 650300
rect 148880 650060 148970 650300
rect 149210 650060 149320 650300
rect 149560 650060 149650 650300
rect 149890 650060 149980 650300
rect 150220 650060 150310 650300
rect 150550 650060 150660 650300
rect 150900 650060 150990 650300
rect 151230 650060 151320 650300
rect 151560 650060 151650 650300
rect 151890 650060 152000 650300
rect 152240 650060 152330 650300
rect 152570 650060 152660 650300
rect 152900 650060 152990 650300
rect 153230 650060 153340 650300
rect 153580 650060 153670 650300
rect 153910 650060 154000 650300
rect 154240 650060 154330 650300
rect 154570 650060 154680 650300
rect 154920 650060 155010 650300
rect 155250 650060 155340 650300
rect 155580 650060 155670 650300
rect 155910 650060 155960 650300
rect 110760 649970 155960 650060
rect 110760 649730 110810 649970
rect 111050 649730 111160 649970
rect 111400 649730 111490 649970
rect 111730 649730 111820 649970
rect 112060 649730 112150 649970
rect 112390 649730 112500 649970
rect 112740 649730 112830 649970
rect 113070 649730 113160 649970
rect 113400 649730 113490 649970
rect 113730 649730 113840 649970
rect 114080 649730 114170 649970
rect 114410 649730 114500 649970
rect 114740 649730 114830 649970
rect 115070 649730 115180 649970
rect 115420 649730 115510 649970
rect 115750 649730 115840 649970
rect 116080 649730 116170 649970
rect 116410 649730 116520 649970
rect 116760 649730 116850 649970
rect 117090 649730 117180 649970
rect 117420 649730 117510 649970
rect 117750 649730 117860 649970
rect 118100 649730 118190 649970
rect 118430 649730 118520 649970
rect 118760 649730 118850 649970
rect 119090 649730 119200 649970
rect 119440 649730 119530 649970
rect 119770 649730 119860 649970
rect 120100 649730 120190 649970
rect 120430 649730 120540 649970
rect 120780 649730 120870 649970
rect 121110 649730 121200 649970
rect 121440 649730 121530 649970
rect 121770 649730 122190 649970
rect 122430 649730 122540 649970
rect 122780 649730 122870 649970
rect 123110 649730 123200 649970
rect 123440 649730 123530 649970
rect 123770 649730 123880 649970
rect 124120 649730 124210 649970
rect 124450 649730 124540 649970
rect 124780 649730 124870 649970
rect 125110 649730 125220 649970
rect 125460 649730 125550 649970
rect 125790 649730 125880 649970
rect 126120 649730 126210 649970
rect 126450 649730 126560 649970
rect 126800 649730 126890 649970
rect 127130 649730 127220 649970
rect 127460 649730 127550 649970
rect 127790 649730 127900 649970
rect 128140 649730 128230 649970
rect 128470 649730 128560 649970
rect 128800 649730 128890 649970
rect 129130 649730 129240 649970
rect 129480 649730 129570 649970
rect 129810 649730 129900 649970
rect 130140 649730 130230 649970
rect 130470 649730 130580 649970
rect 130820 649730 130910 649970
rect 131150 649730 131240 649970
rect 131480 649730 131570 649970
rect 131810 649730 131920 649970
rect 132160 649730 132250 649970
rect 132490 649730 132580 649970
rect 132820 649730 132910 649970
rect 133150 649730 133570 649970
rect 133810 649730 133920 649970
rect 134160 649730 134250 649970
rect 134490 649730 134580 649970
rect 134820 649730 134910 649970
rect 135150 649730 135260 649970
rect 135500 649730 135590 649970
rect 135830 649730 135920 649970
rect 136160 649730 136250 649970
rect 136490 649730 136600 649970
rect 136840 649730 136930 649970
rect 137170 649730 137260 649970
rect 137500 649730 137590 649970
rect 137830 649730 137940 649970
rect 138180 649730 138270 649970
rect 138510 649730 138600 649970
rect 138840 649730 138930 649970
rect 139170 649730 139280 649970
rect 139520 649730 139610 649970
rect 139850 649730 139940 649970
rect 140180 649730 140270 649970
rect 140510 649730 140620 649970
rect 140860 649730 140950 649970
rect 141190 649730 141280 649970
rect 141520 649730 141610 649970
rect 141850 649730 141960 649970
rect 142200 649730 142290 649970
rect 142530 649730 142620 649970
rect 142860 649730 142950 649970
rect 143190 649730 143300 649970
rect 143540 649730 143630 649970
rect 143870 649730 143960 649970
rect 144200 649730 144290 649970
rect 144530 649730 144950 649970
rect 145190 649730 145300 649970
rect 145540 649730 145630 649970
rect 145870 649730 145960 649970
rect 146200 649730 146290 649970
rect 146530 649730 146640 649970
rect 146880 649730 146970 649970
rect 147210 649730 147300 649970
rect 147540 649730 147630 649970
rect 147870 649730 147980 649970
rect 148220 649730 148310 649970
rect 148550 649730 148640 649970
rect 148880 649730 148970 649970
rect 149210 649730 149320 649970
rect 149560 649730 149650 649970
rect 149890 649730 149980 649970
rect 150220 649730 150310 649970
rect 150550 649730 150660 649970
rect 150900 649730 150990 649970
rect 151230 649730 151320 649970
rect 151560 649730 151650 649970
rect 151890 649730 152000 649970
rect 152240 649730 152330 649970
rect 152570 649730 152660 649970
rect 152900 649730 152990 649970
rect 153230 649730 153340 649970
rect 153580 649730 153670 649970
rect 153910 649730 154000 649970
rect 154240 649730 154330 649970
rect 154570 649730 154680 649970
rect 154920 649730 155010 649970
rect 155250 649730 155340 649970
rect 155580 649730 155670 649970
rect 155910 649730 155960 649970
rect 110760 649620 155960 649730
rect 110760 649380 110810 649620
rect 111050 649380 111160 649620
rect 111400 649380 111490 649620
rect 111730 649380 111820 649620
rect 112060 649380 112150 649620
rect 112390 649380 112500 649620
rect 112740 649380 112830 649620
rect 113070 649380 113160 649620
rect 113400 649380 113490 649620
rect 113730 649380 113840 649620
rect 114080 649380 114170 649620
rect 114410 649380 114500 649620
rect 114740 649380 114830 649620
rect 115070 649380 115180 649620
rect 115420 649380 115510 649620
rect 115750 649380 115840 649620
rect 116080 649380 116170 649620
rect 116410 649380 116520 649620
rect 116760 649380 116850 649620
rect 117090 649380 117180 649620
rect 117420 649380 117510 649620
rect 117750 649380 117860 649620
rect 118100 649380 118190 649620
rect 118430 649380 118520 649620
rect 118760 649380 118850 649620
rect 119090 649380 119200 649620
rect 119440 649380 119530 649620
rect 119770 649380 119860 649620
rect 120100 649380 120190 649620
rect 120430 649380 120540 649620
rect 120780 649380 120870 649620
rect 121110 649380 121200 649620
rect 121440 649380 121530 649620
rect 121770 649380 122190 649620
rect 122430 649380 122540 649620
rect 122780 649380 122870 649620
rect 123110 649380 123200 649620
rect 123440 649380 123530 649620
rect 123770 649380 123880 649620
rect 124120 649380 124210 649620
rect 124450 649380 124540 649620
rect 124780 649380 124870 649620
rect 125110 649380 125220 649620
rect 125460 649380 125550 649620
rect 125790 649380 125880 649620
rect 126120 649380 126210 649620
rect 126450 649380 126560 649620
rect 126800 649380 126890 649620
rect 127130 649380 127220 649620
rect 127460 649380 127550 649620
rect 127790 649380 127900 649620
rect 128140 649380 128230 649620
rect 128470 649380 128560 649620
rect 128800 649380 128890 649620
rect 129130 649380 129240 649620
rect 129480 649380 129570 649620
rect 129810 649380 129900 649620
rect 130140 649380 130230 649620
rect 130470 649380 130580 649620
rect 130820 649380 130910 649620
rect 131150 649380 131240 649620
rect 131480 649380 131570 649620
rect 131810 649380 131920 649620
rect 132160 649380 132250 649620
rect 132490 649380 132580 649620
rect 132820 649380 132910 649620
rect 133150 649380 133570 649620
rect 133810 649380 133920 649620
rect 134160 649380 134250 649620
rect 134490 649380 134580 649620
rect 134820 649380 134910 649620
rect 135150 649380 135260 649620
rect 135500 649380 135590 649620
rect 135830 649380 135920 649620
rect 136160 649380 136250 649620
rect 136490 649380 136600 649620
rect 136840 649380 136930 649620
rect 137170 649380 137260 649620
rect 137500 649380 137590 649620
rect 137830 649380 137940 649620
rect 138180 649380 138270 649620
rect 138510 649380 138600 649620
rect 138840 649380 138930 649620
rect 139170 649380 139280 649620
rect 139520 649380 139610 649620
rect 139850 649380 139940 649620
rect 140180 649380 140270 649620
rect 140510 649380 140620 649620
rect 140860 649380 140950 649620
rect 141190 649380 141280 649620
rect 141520 649380 141610 649620
rect 141850 649380 141960 649620
rect 142200 649380 142290 649620
rect 142530 649380 142620 649620
rect 142860 649380 142950 649620
rect 143190 649380 143300 649620
rect 143540 649380 143630 649620
rect 143870 649380 143960 649620
rect 144200 649380 144290 649620
rect 144530 649380 144950 649620
rect 145190 649380 145300 649620
rect 145540 649380 145630 649620
rect 145870 649380 145960 649620
rect 146200 649380 146290 649620
rect 146530 649380 146640 649620
rect 146880 649380 146970 649620
rect 147210 649380 147300 649620
rect 147540 649380 147630 649620
rect 147870 649380 147980 649620
rect 148220 649380 148310 649620
rect 148550 649380 148640 649620
rect 148880 649380 148970 649620
rect 149210 649380 149320 649620
rect 149560 649380 149650 649620
rect 149890 649380 149980 649620
rect 150220 649380 150310 649620
rect 150550 649380 150660 649620
rect 150900 649380 150990 649620
rect 151230 649380 151320 649620
rect 151560 649380 151650 649620
rect 151890 649380 152000 649620
rect 152240 649380 152330 649620
rect 152570 649380 152660 649620
rect 152900 649380 152990 649620
rect 153230 649380 153340 649620
rect 153580 649380 153670 649620
rect 153910 649380 154000 649620
rect 154240 649380 154330 649620
rect 154570 649380 154680 649620
rect 154920 649380 155010 649620
rect 155250 649380 155340 649620
rect 155580 649380 155670 649620
rect 155910 649380 155960 649620
rect 110760 649330 155960 649380
rect 576129 649131 576450 679639
rect 221900 648810 576450 649131
rect 196200 647380 197220 647400
rect 196200 647310 196680 647380
rect 196750 647310 196780 647380
rect 196850 647310 196880 647380
rect 196950 647310 197220 647380
rect 196200 647290 197220 647310
rect 196200 647220 196680 647290
rect 196750 647220 196780 647290
rect 196850 647220 196880 647290
rect 196950 647220 197220 647290
rect 196200 645944 197220 647220
rect 98509 644924 197220 645944
rect 200788 647380 201808 647400
rect 200788 647310 201238 647380
rect 201308 647310 201338 647380
rect 201408 647310 201438 647380
rect 201508 647310 201808 647380
rect 200788 647290 201808 647310
rect 200788 647220 201238 647290
rect 201308 647220 201338 647290
rect 201408 647220 201438 647290
rect 201508 647220 201808 647290
rect 200788 643561 201808 647220
rect 94338 642541 201808 643561
<< via4 >>
rect 16352 703500 16652 703800
rect 16852 703500 17152 703800
rect 17352 703500 17652 703800
rect 17852 703500 18152 703800
rect 18352 703500 18652 703800
rect 18852 703500 19152 703800
rect 19352 703500 19652 703800
rect 19852 703500 20152 703800
rect 20352 703500 20652 703800
rect 20852 703500 21152 703800
rect 16352 703000 16652 703300
rect 16852 703000 17152 703300
rect 17352 703000 17652 703300
rect 17852 703000 18152 703300
rect 18352 703000 18652 703300
rect 18852 703000 19152 703300
rect 19352 703000 19652 703300
rect 19852 703000 20152 703300
rect 20352 703000 20652 703300
rect 20852 703000 21152 703300
rect 16352 702500 16652 702800
rect 16852 702500 17152 702800
rect 17352 702500 17652 702800
rect 17852 702500 18152 702800
rect 18352 702500 18652 702800
rect 18852 702500 19152 702800
rect 19352 702500 19652 702800
rect 19852 702500 20152 702800
rect 20352 702500 20652 702800
rect 20852 702500 21152 702800
rect 200 684900 500 685200
rect 700 684900 1000 685200
rect 1200 684900 1500 685200
rect 200 684400 500 684700
rect 700 684400 1000 684700
rect 1200 684400 1500 684700
rect 200 683900 500 684200
rect 700 683900 1000 684200
rect 1200 683900 1500 684200
rect 200 683400 500 683700
rect 700 683400 1000 683700
rect 1200 683400 1500 683700
rect 200 682900 500 683200
rect 700 682900 1000 683200
rect 1200 682900 1500 683200
rect 200 682400 500 682700
rect 700 682400 1000 682700
rect 1200 682400 1500 682700
rect 200 681900 500 682200
rect 700 681900 1000 682200
rect 1200 681900 1500 682200
rect 200 681400 500 681700
rect 700 681400 1000 681700
rect 1200 681400 1500 681700
rect 200 680900 500 681200
rect 700 680900 1000 681200
rect 1200 680900 1500 681200
rect 200 680400 500 680700
rect 700 680400 1000 680700
rect 1200 680400 1500 680700
rect 110890 683460 111130 683700
rect 111220 683460 111460 683700
rect 111550 683460 111790 683700
rect 111880 683460 112120 683700
rect 112210 683460 112450 683700
rect 112540 683460 112780 683700
rect 112870 683460 113110 683700
rect 113200 683460 113440 683700
rect 113530 683460 113770 683700
rect 113860 683460 114100 683700
rect 114190 683460 114430 683700
rect 114520 683460 114760 683700
rect 114850 683460 115090 683700
rect 115180 683460 115420 683700
rect 115510 683460 115750 683700
rect 115840 683460 116080 683700
rect 116170 683460 116410 683700
rect 116500 683460 116740 683700
rect 116830 683460 117070 683700
rect 117160 683460 117400 683700
rect 117490 683460 117730 683700
rect 117820 683460 118060 683700
rect 118150 683460 118390 683700
rect 118480 683460 118720 683700
rect 118810 683460 119050 683700
rect 119140 683460 119380 683700
rect 119470 683460 119710 683700
rect 119800 683460 120040 683700
rect 120130 683460 120370 683700
rect 120460 683460 120700 683700
rect 120790 683460 121030 683700
rect 121120 683460 121360 683700
rect 121450 683460 121690 683700
rect 122270 683460 122510 683700
rect 122600 683460 122840 683700
rect 122930 683460 123170 683700
rect 123260 683460 123500 683700
rect 123590 683460 123830 683700
rect 123920 683460 124160 683700
rect 124250 683460 124490 683700
rect 124580 683460 124820 683700
rect 124910 683460 125150 683700
rect 125240 683460 125480 683700
rect 125570 683460 125810 683700
rect 125900 683460 126140 683700
rect 126230 683460 126470 683700
rect 126560 683460 126800 683700
rect 126890 683460 127130 683700
rect 127220 683460 127460 683700
rect 127550 683460 127790 683700
rect 127880 683460 128120 683700
rect 128210 683460 128450 683700
rect 128540 683460 128780 683700
rect 128870 683460 129110 683700
rect 129200 683460 129440 683700
rect 129530 683460 129770 683700
rect 129860 683460 130100 683700
rect 130190 683460 130430 683700
rect 130520 683460 130760 683700
rect 130850 683460 131090 683700
rect 131180 683460 131420 683700
rect 131510 683460 131750 683700
rect 131840 683460 132080 683700
rect 132170 683460 132410 683700
rect 132500 683460 132740 683700
rect 132830 683460 133070 683700
rect 133650 683460 133890 683700
rect 133980 683460 134220 683700
rect 134310 683460 134550 683700
rect 134640 683460 134880 683700
rect 134970 683460 135210 683700
rect 135300 683460 135540 683700
rect 135630 683460 135870 683700
rect 135960 683460 136200 683700
rect 136290 683460 136530 683700
rect 136620 683460 136860 683700
rect 136950 683460 137190 683700
rect 137280 683460 137520 683700
rect 137610 683460 137850 683700
rect 137940 683460 138180 683700
rect 138270 683460 138510 683700
rect 138600 683460 138840 683700
rect 138930 683460 139170 683700
rect 139260 683460 139500 683700
rect 139590 683460 139830 683700
rect 139920 683460 140160 683700
rect 140250 683460 140490 683700
rect 140580 683460 140820 683700
rect 140910 683460 141150 683700
rect 141240 683460 141480 683700
rect 141570 683460 141810 683700
rect 141900 683460 142140 683700
rect 142230 683460 142470 683700
rect 142560 683460 142800 683700
rect 142890 683460 143130 683700
rect 143220 683460 143460 683700
rect 143550 683460 143790 683700
rect 143880 683460 144120 683700
rect 144210 683460 144450 683700
rect 145030 683460 145270 683700
rect 145360 683460 145600 683700
rect 145690 683460 145930 683700
rect 146020 683460 146260 683700
rect 146350 683460 146590 683700
rect 146680 683460 146920 683700
rect 147010 683460 147250 683700
rect 147340 683460 147580 683700
rect 147670 683460 147910 683700
rect 148000 683460 148240 683700
rect 148330 683460 148570 683700
rect 148660 683460 148900 683700
rect 148990 683460 149230 683700
rect 149320 683460 149560 683700
rect 149650 683460 149890 683700
rect 149980 683460 150220 683700
rect 150310 683460 150550 683700
rect 150640 683460 150880 683700
rect 150970 683460 151210 683700
rect 151300 683460 151540 683700
rect 151630 683460 151870 683700
rect 151960 683460 152200 683700
rect 152290 683460 152530 683700
rect 152620 683460 152860 683700
rect 152950 683460 153190 683700
rect 153280 683460 153520 683700
rect 153610 683460 153850 683700
rect 153940 683460 154180 683700
rect 154270 683460 154510 683700
rect 154600 683460 154840 683700
rect 154930 683460 155170 683700
rect 155260 683460 155500 683700
rect 155590 683460 155830 683700
rect 107220 678740 107480 678980
rect 107580 678740 107840 678980
rect 107940 678740 108200 678980
rect 108300 678740 108560 678980
rect 157520 678739 157780 678979
rect 157880 678739 158140 678979
rect 158240 678739 158500 678979
rect 158600 678739 158860 678979
rect 107220 678400 107480 678640
rect 107580 678400 107840 678640
rect 107940 678400 108200 678640
rect 108300 678400 108560 678640
rect 157520 678399 157780 678639
rect 157880 678399 158140 678639
rect 158240 678399 158500 678639
rect 158600 678399 158860 678639
rect 107220 678060 107480 678300
rect 107580 678060 107840 678300
rect 107940 678060 108200 678300
rect 108300 678060 108560 678300
rect 157520 678059 157780 678299
rect 157880 678059 158140 678299
rect 158240 678059 158500 678299
rect 158600 678059 158860 678299
rect 107220 677720 107480 677960
rect 107580 677720 107840 677960
rect 107940 677720 108200 677960
rect 108300 677720 108560 677960
rect 157520 677719 157780 677959
rect 157880 677719 158140 677959
rect 158240 677719 158500 677959
rect 158600 677719 158860 677959
rect 107220 677380 107480 677620
rect 107580 677380 107840 677620
rect 107940 677380 108200 677620
rect 108300 677380 108560 677620
rect 157520 677379 157780 677619
rect 157880 677379 158140 677619
rect 158240 677379 158500 677619
rect 158600 677379 158860 677619
rect 107220 677040 107480 677280
rect 107580 677040 107840 677280
rect 107940 677040 108200 677280
rect 108300 677040 108560 677280
rect 157520 677039 157780 677279
rect 157880 677039 158140 677279
rect 158240 677039 158500 677279
rect 158600 677039 158860 677279
rect 107220 676700 107480 676940
rect 107580 676700 107840 676940
rect 107940 676700 108200 676940
rect 108300 676700 108560 676940
rect 157520 676699 157780 676939
rect 157880 676699 158140 676939
rect 158240 676699 158500 676939
rect 158600 676699 158860 676939
rect 107220 676360 107480 676600
rect 107580 676360 107840 676600
rect 107940 676360 108200 676600
rect 108300 676360 108560 676600
rect 157520 676359 157780 676599
rect 157880 676359 158140 676599
rect 158240 676359 158500 676599
rect 158600 676359 158860 676599
rect 107220 676020 107480 676260
rect 107580 676020 107840 676260
rect 107940 676020 108200 676260
rect 108300 676020 108560 676260
rect 157520 676019 157780 676259
rect 157880 676019 158140 676259
rect 158240 676019 158500 676259
rect 158600 676019 158860 676259
rect 107220 675680 107480 675920
rect 107580 675680 107840 675920
rect 107940 675680 108200 675920
rect 108300 675680 108560 675920
rect 157520 675679 157780 675919
rect 157880 675679 158140 675919
rect 158240 675679 158500 675919
rect 158600 675679 158860 675919
rect 107220 675340 107480 675580
rect 107580 675340 107840 675580
rect 107940 675340 108200 675580
rect 108300 675340 108560 675580
rect 157520 675339 157780 675579
rect 157880 675339 158140 675579
rect 158240 675339 158500 675579
rect 158600 675339 158860 675579
rect 107220 675000 107480 675240
rect 107580 675000 107840 675240
rect 107940 675000 108200 675240
rect 108300 675000 108560 675240
rect 157520 674999 157780 675239
rect 157880 674999 158140 675239
rect 158240 674999 158500 675239
rect 158600 674999 158860 675239
rect 107220 674660 107480 674900
rect 107580 674660 107840 674900
rect 107940 674660 108200 674900
rect 108300 674660 108560 674900
rect 157520 674659 157780 674899
rect 157880 674659 158140 674899
rect 158240 674659 158500 674899
rect 158600 674659 158860 674899
rect 107220 674320 107480 674560
rect 107580 674320 107840 674560
rect 107940 674320 108200 674560
rect 108300 674320 108560 674560
rect 157520 674319 157780 674559
rect 157880 674319 158140 674559
rect 158240 674319 158500 674559
rect 158600 674319 158860 674559
rect 110890 660520 111130 660760
rect 111220 660520 111460 660760
rect 111550 660520 111790 660760
rect 111880 660520 112120 660760
rect 112210 660520 112450 660760
rect 112540 660520 112780 660760
rect 112870 660520 113110 660760
rect 113200 660520 113440 660760
rect 113530 660520 113770 660760
rect 113860 660520 114100 660760
rect 114190 660520 114430 660760
rect 114520 660520 114760 660760
rect 114850 660520 115090 660760
rect 115180 660520 115420 660760
rect 115510 660520 115750 660760
rect 115840 660520 116080 660760
rect 116170 660520 116410 660760
rect 116500 660520 116740 660760
rect 116830 660520 117070 660760
rect 117160 660520 117400 660760
rect 117490 660520 117730 660760
rect 117820 660520 118060 660760
rect 118150 660520 118390 660760
rect 118480 660520 118720 660760
rect 118810 660520 119050 660760
rect 119140 660520 119380 660760
rect 119470 660520 119710 660760
rect 119800 660520 120040 660760
rect 120130 660520 120370 660760
rect 120460 660520 120700 660760
rect 120790 660520 121030 660760
rect 121120 660520 121360 660760
rect 121450 660520 121690 660760
rect 122270 660520 122510 660760
rect 122600 660520 122840 660760
rect 122930 660520 123170 660760
rect 123260 660520 123500 660760
rect 123590 660520 123830 660760
rect 123920 660520 124160 660760
rect 124250 660520 124490 660760
rect 124580 660520 124820 660760
rect 124910 660520 125150 660760
rect 125240 660520 125480 660760
rect 125570 660520 125810 660760
rect 125900 660520 126140 660760
rect 126230 660520 126470 660760
rect 126560 660520 126800 660760
rect 126890 660520 127130 660760
rect 127220 660520 127460 660760
rect 127550 660520 127790 660760
rect 127880 660520 128120 660760
rect 128210 660520 128450 660760
rect 128540 660520 128780 660760
rect 128870 660520 129110 660760
rect 129200 660520 129440 660760
rect 129530 660520 129770 660760
rect 129860 660520 130100 660760
rect 130190 660520 130430 660760
rect 130520 660520 130760 660760
rect 130850 660520 131090 660760
rect 131180 660520 131420 660760
rect 131510 660520 131750 660760
rect 131840 660520 132080 660760
rect 132170 660520 132410 660760
rect 132500 660520 132740 660760
rect 132830 660520 133070 660760
rect 133650 660520 133890 660760
rect 133980 660520 134220 660760
rect 134310 660520 134550 660760
rect 134640 660520 134880 660760
rect 134970 660520 135210 660760
rect 135300 660520 135540 660760
rect 135630 660520 135870 660760
rect 135960 660520 136200 660760
rect 136290 660520 136530 660760
rect 136620 660520 136860 660760
rect 136950 660520 137190 660760
rect 137280 660520 137520 660760
rect 137610 660520 137850 660760
rect 137940 660520 138180 660760
rect 138270 660520 138510 660760
rect 138600 660520 138840 660760
rect 138930 660520 139170 660760
rect 139260 660520 139500 660760
rect 139590 660520 139830 660760
rect 139920 660520 140160 660760
rect 140250 660520 140490 660760
rect 140580 660520 140820 660760
rect 140910 660520 141150 660760
rect 141240 660520 141480 660760
rect 141570 660520 141810 660760
rect 141900 660520 142140 660760
rect 142230 660520 142470 660760
rect 142560 660520 142800 660760
rect 142890 660520 143130 660760
rect 143220 660520 143460 660760
rect 143550 660520 143790 660760
rect 143880 660520 144120 660760
rect 144210 660520 144450 660760
rect 145030 660520 145270 660760
rect 145360 660520 145600 660760
rect 145690 660520 145930 660760
rect 146020 660520 146260 660760
rect 146350 660520 146590 660760
rect 146680 660520 146920 660760
rect 147010 660520 147250 660760
rect 147340 660520 147580 660760
rect 147670 660520 147910 660760
rect 148000 660520 148240 660760
rect 148330 660520 148570 660760
rect 148660 660520 148900 660760
rect 148990 660520 149230 660760
rect 149320 660520 149560 660760
rect 149650 660520 149890 660760
rect 149980 660520 150220 660760
rect 150310 660520 150550 660760
rect 150640 660520 150880 660760
rect 150970 660520 151210 660760
rect 151300 660520 151540 660760
rect 151630 660520 151870 660760
rect 151960 660520 152200 660760
rect 152290 660520 152530 660760
rect 152620 660520 152860 660760
rect 152950 660520 153190 660760
rect 153280 660520 153520 660760
rect 153610 660520 153850 660760
rect 153940 660520 154180 660760
rect 154270 660520 154510 660760
rect 154600 660520 154840 660760
rect 154930 660520 155170 660760
rect 155260 660520 155500 660760
rect 155590 660520 155830 660760
<< mimcap2 >>
rect 110790 694840 121790 694860
rect 110790 694600 110810 694840
rect 111050 694600 111140 694840
rect 111380 694600 111470 694840
rect 111710 694600 111800 694840
rect 112040 694600 112150 694840
rect 112390 694600 112480 694840
rect 112720 694600 112810 694840
rect 113050 694600 113140 694840
rect 113380 694600 113490 694840
rect 113730 694600 113820 694840
rect 114060 694600 114150 694840
rect 114390 694600 114480 694840
rect 114720 694600 114830 694840
rect 115070 694600 115160 694840
rect 115400 694600 115490 694840
rect 115730 694600 115820 694840
rect 116060 694600 116170 694840
rect 116410 694600 116500 694840
rect 116740 694600 116830 694840
rect 117070 694600 117160 694840
rect 117400 694600 117510 694840
rect 117750 694600 117840 694840
rect 118080 694600 118170 694840
rect 118410 694600 118500 694840
rect 118740 694600 118850 694840
rect 119090 694600 119180 694840
rect 119420 694600 119510 694840
rect 119750 694600 119840 694840
rect 120080 694600 120190 694840
rect 120430 694600 120520 694840
rect 120760 694600 120850 694840
rect 121090 694600 121180 694840
rect 121420 694600 121530 694840
rect 121770 694600 121790 694840
rect 110790 694490 121790 694600
rect 110790 694250 110810 694490
rect 111050 694250 111140 694490
rect 111380 694250 111470 694490
rect 111710 694250 111800 694490
rect 112040 694250 112150 694490
rect 112390 694250 112480 694490
rect 112720 694250 112810 694490
rect 113050 694250 113140 694490
rect 113380 694250 113490 694490
rect 113730 694250 113820 694490
rect 114060 694250 114150 694490
rect 114390 694250 114480 694490
rect 114720 694250 114830 694490
rect 115070 694250 115160 694490
rect 115400 694250 115490 694490
rect 115730 694250 115820 694490
rect 116060 694250 116170 694490
rect 116410 694250 116500 694490
rect 116740 694250 116830 694490
rect 117070 694250 117160 694490
rect 117400 694250 117510 694490
rect 117750 694250 117840 694490
rect 118080 694250 118170 694490
rect 118410 694250 118500 694490
rect 118740 694250 118850 694490
rect 119090 694250 119180 694490
rect 119420 694250 119510 694490
rect 119750 694250 119840 694490
rect 120080 694250 120190 694490
rect 120430 694250 120520 694490
rect 120760 694250 120850 694490
rect 121090 694250 121180 694490
rect 121420 694250 121530 694490
rect 121770 694250 121790 694490
rect 110790 694160 121790 694250
rect 110790 693920 110810 694160
rect 111050 693920 111140 694160
rect 111380 693920 111470 694160
rect 111710 693920 111800 694160
rect 112040 693920 112150 694160
rect 112390 693920 112480 694160
rect 112720 693920 112810 694160
rect 113050 693920 113140 694160
rect 113380 693920 113490 694160
rect 113730 693920 113820 694160
rect 114060 693920 114150 694160
rect 114390 693920 114480 694160
rect 114720 693920 114830 694160
rect 115070 693920 115160 694160
rect 115400 693920 115490 694160
rect 115730 693920 115820 694160
rect 116060 693920 116170 694160
rect 116410 693920 116500 694160
rect 116740 693920 116830 694160
rect 117070 693920 117160 694160
rect 117400 693920 117510 694160
rect 117750 693920 117840 694160
rect 118080 693920 118170 694160
rect 118410 693920 118500 694160
rect 118740 693920 118850 694160
rect 119090 693920 119180 694160
rect 119420 693920 119510 694160
rect 119750 693920 119840 694160
rect 120080 693920 120190 694160
rect 120430 693920 120520 694160
rect 120760 693920 120850 694160
rect 121090 693920 121180 694160
rect 121420 693920 121530 694160
rect 121770 693920 121790 694160
rect 110790 693830 121790 693920
rect 110790 693590 110810 693830
rect 111050 693590 111140 693830
rect 111380 693590 111470 693830
rect 111710 693590 111800 693830
rect 112040 693590 112150 693830
rect 112390 693590 112480 693830
rect 112720 693590 112810 693830
rect 113050 693590 113140 693830
rect 113380 693590 113490 693830
rect 113730 693590 113820 693830
rect 114060 693590 114150 693830
rect 114390 693590 114480 693830
rect 114720 693590 114830 693830
rect 115070 693590 115160 693830
rect 115400 693590 115490 693830
rect 115730 693590 115820 693830
rect 116060 693590 116170 693830
rect 116410 693590 116500 693830
rect 116740 693590 116830 693830
rect 117070 693590 117160 693830
rect 117400 693590 117510 693830
rect 117750 693590 117840 693830
rect 118080 693590 118170 693830
rect 118410 693590 118500 693830
rect 118740 693590 118850 693830
rect 119090 693590 119180 693830
rect 119420 693590 119510 693830
rect 119750 693590 119840 693830
rect 120080 693590 120190 693830
rect 120430 693590 120520 693830
rect 120760 693590 120850 693830
rect 121090 693590 121180 693830
rect 121420 693590 121530 693830
rect 121770 693590 121790 693830
rect 110790 693500 121790 693590
rect 110790 693260 110810 693500
rect 111050 693260 111140 693500
rect 111380 693260 111470 693500
rect 111710 693260 111800 693500
rect 112040 693260 112150 693500
rect 112390 693260 112480 693500
rect 112720 693260 112810 693500
rect 113050 693260 113140 693500
rect 113380 693260 113490 693500
rect 113730 693260 113820 693500
rect 114060 693260 114150 693500
rect 114390 693260 114480 693500
rect 114720 693260 114830 693500
rect 115070 693260 115160 693500
rect 115400 693260 115490 693500
rect 115730 693260 115820 693500
rect 116060 693260 116170 693500
rect 116410 693260 116500 693500
rect 116740 693260 116830 693500
rect 117070 693260 117160 693500
rect 117400 693260 117510 693500
rect 117750 693260 117840 693500
rect 118080 693260 118170 693500
rect 118410 693260 118500 693500
rect 118740 693260 118850 693500
rect 119090 693260 119180 693500
rect 119420 693260 119510 693500
rect 119750 693260 119840 693500
rect 120080 693260 120190 693500
rect 120430 693260 120520 693500
rect 120760 693260 120850 693500
rect 121090 693260 121180 693500
rect 121420 693260 121530 693500
rect 121770 693260 121790 693500
rect 110790 693150 121790 693260
rect 110790 692910 110810 693150
rect 111050 692910 111140 693150
rect 111380 692910 111470 693150
rect 111710 692910 111800 693150
rect 112040 692910 112150 693150
rect 112390 692910 112480 693150
rect 112720 692910 112810 693150
rect 113050 692910 113140 693150
rect 113380 692910 113490 693150
rect 113730 692910 113820 693150
rect 114060 692910 114150 693150
rect 114390 692910 114480 693150
rect 114720 692910 114830 693150
rect 115070 692910 115160 693150
rect 115400 692910 115490 693150
rect 115730 692910 115820 693150
rect 116060 692910 116170 693150
rect 116410 692910 116500 693150
rect 116740 692910 116830 693150
rect 117070 692910 117160 693150
rect 117400 692910 117510 693150
rect 117750 692910 117840 693150
rect 118080 692910 118170 693150
rect 118410 692910 118500 693150
rect 118740 692910 118850 693150
rect 119090 692910 119180 693150
rect 119420 692910 119510 693150
rect 119750 692910 119840 693150
rect 120080 692910 120190 693150
rect 120430 692910 120520 693150
rect 120760 692910 120850 693150
rect 121090 692910 121180 693150
rect 121420 692910 121530 693150
rect 121770 692910 121790 693150
rect 110790 692820 121790 692910
rect 110790 692580 110810 692820
rect 111050 692580 111140 692820
rect 111380 692580 111470 692820
rect 111710 692580 111800 692820
rect 112040 692580 112150 692820
rect 112390 692580 112480 692820
rect 112720 692580 112810 692820
rect 113050 692580 113140 692820
rect 113380 692580 113490 692820
rect 113730 692580 113820 692820
rect 114060 692580 114150 692820
rect 114390 692580 114480 692820
rect 114720 692580 114830 692820
rect 115070 692580 115160 692820
rect 115400 692580 115490 692820
rect 115730 692580 115820 692820
rect 116060 692580 116170 692820
rect 116410 692580 116500 692820
rect 116740 692580 116830 692820
rect 117070 692580 117160 692820
rect 117400 692580 117510 692820
rect 117750 692580 117840 692820
rect 118080 692580 118170 692820
rect 118410 692580 118500 692820
rect 118740 692580 118850 692820
rect 119090 692580 119180 692820
rect 119420 692580 119510 692820
rect 119750 692580 119840 692820
rect 120080 692580 120190 692820
rect 120430 692580 120520 692820
rect 120760 692580 120850 692820
rect 121090 692580 121180 692820
rect 121420 692580 121530 692820
rect 121770 692580 121790 692820
rect 110790 692490 121790 692580
rect 110790 692250 110810 692490
rect 111050 692250 111140 692490
rect 111380 692250 111470 692490
rect 111710 692250 111800 692490
rect 112040 692250 112150 692490
rect 112390 692250 112480 692490
rect 112720 692250 112810 692490
rect 113050 692250 113140 692490
rect 113380 692250 113490 692490
rect 113730 692250 113820 692490
rect 114060 692250 114150 692490
rect 114390 692250 114480 692490
rect 114720 692250 114830 692490
rect 115070 692250 115160 692490
rect 115400 692250 115490 692490
rect 115730 692250 115820 692490
rect 116060 692250 116170 692490
rect 116410 692250 116500 692490
rect 116740 692250 116830 692490
rect 117070 692250 117160 692490
rect 117400 692250 117510 692490
rect 117750 692250 117840 692490
rect 118080 692250 118170 692490
rect 118410 692250 118500 692490
rect 118740 692250 118850 692490
rect 119090 692250 119180 692490
rect 119420 692250 119510 692490
rect 119750 692250 119840 692490
rect 120080 692250 120190 692490
rect 120430 692250 120520 692490
rect 120760 692250 120850 692490
rect 121090 692250 121180 692490
rect 121420 692250 121530 692490
rect 121770 692250 121790 692490
rect 110790 692160 121790 692250
rect 110790 691920 110810 692160
rect 111050 691920 111140 692160
rect 111380 691920 111470 692160
rect 111710 691920 111800 692160
rect 112040 691920 112150 692160
rect 112390 691920 112480 692160
rect 112720 691920 112810 692160
rect 113050 691920 113140 692160
rect 113380 691920 113490 692160
rect 113730 691920 113820 692160
rect 114060 691920 114150 692160
rect 114390 691920 114480 692160
rect 114720 691920 114830 692160
rect 115070 691920 115160 692160
rect 115400 691920 115490 692160
rect 115730 691920 115820 692160
rect 116060 691920 116170 692160
rect 116410 691920 116500 692160
rect 116740 691920 116830 692160
rect 117070 691920 117160 692160
rect 117400 691920 117510 692160
rect 117750 691920 117840 692160
rect 118080 691920 118170 692160
rect 118410 691920 118500 692160
rect 118740 691920 118850 692160
rect 119090 691920 119180 692160
rect 119420 691920 119510 692160
rect 119750 691920 119840 692160
rect 120080 691920 120190 692160
rect 120430 691920 120520 692160
rect 120760 691920 120850 692160
rect 121090 691920 121180 692160
rect 121420 691920 121530 692160
rect 121770 691920 121790 692160
rect 110790 691810 121790 691920
rect 110790 691570 110810 691810
rect 111050 691570 111140 691810
rect 111380 691570 111470 691810
rect 111710 691570 111800 691810
rect 112040 691570 112150 691810
rect 112390 691570 112480 691810
rect 112720 691570 112810 691810
rect 113050 691570 113140 691810
rect 113380 691570 113490 691810
rect 113730 691570 113820 691810
rect 114060 691570 114150 691810
rect 114390 691570 114480 691810
rect 114720 691570 114830 691810
rect 115070 691570 115160 691810
rect 115400 691570 115490 691810
rect 115730 691570 115820 691810
rect 116060 691570 116170 691810
rect 116410 691570 116500 691810
rect 116740 691570 116830 691810
rect 117070 691570 117160 691810
rect 117400 691570 117510 691810
rect 117750 691570 117840 691810
rect 118080 691570 118170 691810
rect 118410 691570 118500 691810
rect 118740 691570 118850 691810
rect 119090 691570 119180 691810
rect 119420 691570 119510 691810
rect 119750 691570 119840 691810
rect 120080 691570 120190 691810
rect 120430 691570 120520 691810
rect 120760 691570 120850 691810
rect 121090 691570 121180 691810
rect 121420 691570 121530 691810
rect 121770 691570 121790 691810
rect 110790 691480 121790 691570
rect 110790 691240 110810 691480
rect 111050 691240 111140 691480
rect 111380 691240 111470 691480
rect 111710 691240 111800 691480
rect 112040 691240 112150 691480
rect 112390 691240 112480 691480
rect 112720 691240 112810 691480
rect 113050 691240 113140 691480
rect 113380 691240 113490 691480
rect 113730 691240 113820 691480
rect 114060 691240 114150 691480
rect 114390 691240 114480 691480
rect 114720 691240 114830 691480
rect 115070 691240 115160 691480
rect 115400 691240 115490 691480
rect 115730 691240 115820 691480
rect 116060 691240 116170 691480
rect 116410 691240 116500 691480
rect 116740 691240 116830 691480
rect 117070 691240 117160 691480
rect 117400 691240 117510 691480
rect 117750 691240 117840 691480
rect 118080 691240 118170 691480
rect 118410 691240 118500 691480
rect 118740 691240 118850 691480
rect 119090 691240 119180 691480
rect 119420 691240 119510 691480
rect 119750 691240 119840 691480
rect 120080 691240 120190 691480
rect 120430 691240 120520 691480
rect 120760 691240 120850 691480
rect 121090 691240 121180 691480
rect 121420 691240 121530 691480
rect 121770 691240 121790 691480
rect 110790 691150 121790 691240
rect 110790 690910 110810 691150
rect 111050 690910 111140 691150
rect 111380 690910 111470 691150
rect 111710 690910 111800 691150
rect 112040 690910 112150 691150
rect 112390 690910 112480 691150
rect 112720 690910 112810 691150
rect 113050 690910 113140 691150
rect 113380 690910 113490 691150
rect 113730 690910 113820 691150
rect 114060 690910 114150 691150
rect 114390 690910 114480 691150
rect 114720 690910 114830 691150
rect 115070 690910 115160 691150
rect 115400 690910 115490 691150
rect 115730 690910 115820 691150
rect 116060 690910 116170 691150
rect 116410 690910 116500 691150
rect 116740 690910 116830 691150
rect 117070 690910 117160 691150
rect 117400 690910 117510 691150
rect 117750 690910 117840 691150
rect 118080 690910 118170 691150
rect 118410 690910 118500 691150
rect 118740 690910 118850 691150
rect 119090 690910 119180 691150
rect 119420 690910 119510 691150
rect 119750 690910 119840 691150
rect 120080 690910 120190 691150
rect 120430 690910 120520 691150
rect 120760 690910 120850 691150
rect 121090 690910 121180 691150
rect 121420 690910 121530 691150
rect 121770 690910 121790 691150
rect 110790 690820 121790 690910
rect 110790 690580 110810 690820
rect 111050 690580 111140 690820
rect 111380 690580 111470 690820
rect 111710 690580 111800 690820
rect 112040 690580 112150 690820
rect 112390 690580 112480 690820
rect 112720 690580 112810 690820
rect 113050 690580 113140 690820
rect 113380 690580 113490 690820
rect 113730 690580 113820 690820
rect 114060 690580 114150 690820
rect 114390 690580 114480 690820
rect 114720 690580 114830 690820
rect 115070 690580 115160 690820
rect 115400 690580 115490 690820
rect 115730 690580 115820 690820
rect 116060 690580 116170 690820
rect 116410 690580 116500 690820
rect 116740 690580 116830 690820
rect 117070 690580 117160 690820
rect 117400 690580 117510 690820
rect 117750 690580 117840 690820
rect 118080 690580 118170 690820
rect 118410 690580 118500 690820
rect 118740 690580 118850 690820
rect 119090 690580 119180 690820
rect 119420 690580 119510 690820
rect 119750 690580 119840 690820
rect 120080 690580 120190 690820
rect 120430 690580 120520 690820
rect 120760 690580 120850 690820
rect 121090 690580 121180 690820
rect 121420 690580 121530 690820
rect 121770 690580 121790 690820
rect 110790 690470 121790 690580
rect 110790 690230 110810 690470
rect 111050 690230 111140 690470
rect 111380 690230 111470 690470
rect 111710 690230 111800 690470
rect 112040 690230 112150 690470
rect 112390 690230 112480 690470
rect 112720 690230 112810 690470
rect 113050 690230 113140 690470
rect 113380 690230 113490 690470
rect 113730 690230 113820 690470
rect 114060 690230 114150 690470
rect 114390 690230 114480 690470
rect 114720 690230 114830 690470
rect 115070 690230 115160 690470
rect 115400 690230 115490 690470
rect 115730 690230 115820 690470
rect 116060 690230 116170 690470
rect 116410 690230 116500 690470
rect 116740 690230 116830 690470
rect 117070 690230 117160 690470
rect 117400 690230 117510 690470
rect 117750 690230 117840 690470
rect 118080 690230 118170 690470
rect 118410 690230 118500 690470
rect 118740 690230 118850 690470
rect 119090 690230 119180 690470
rect 119420 690230 119510 690470
rect 119750 690230 119840 690470
rect 120080 690230 120190 690470
rect 120430 690230 120520 690470
rect 120760 690230 120850 690470
rect 121090 690230 121180 690470
rect 121420 690230 121530 690470
rect 121770 690230 121790 690470
rect 110790 690140 121790 690230
rect 110790 689900 110810 690140
rect 111050 689900 111140 690140
rect 111380 689900 111470 690140
rect 111710 689900 111800 690140
rect 112040 689900 112150 690140
rect 112390 689900 112480 690140
rect 112720 689900 112810 690140
rect 113050 689900 113140 690140
rect 113380 689900 113490 690140
rect 113730 689900 113820 690140
rect 114060 689900 114150 690140
rect 114390 689900 114480 690140
rect 114720 689900 114830 690140
rect 115070 689900 115160 690140
rect 115400 689900 115490 690140
rect 115730 689900 115820 690140
rect 116060 689900 116170 690140
rect 116410 689900 116500 690140
rect 116740 689900 116830 690140
rect 117070 689900 117160 690140
rect 117400 689900 117510 690140
rect 117750 689900 117840 690140
rect 118080 689900 118170 690140
rect 118410 689900 118500 690140
rect 118740 689900 118850 690140
rect 119090 689900 119180 690140
rect 119420 689900 119510 690140
rect 119750 689900 119840 690140
rect 120080 689900 120190 690140
rect 120430 689900 120520 690140
rect 120760 689900 120850 690140
rect 121090 689900 121180 690140
rect 121420 689900 121530 690140
rect 121770 689900 121790 690140
rect 110790 689810 121790 689900
rect 110790 689570 110810 689810
rect 111050 689570 111140 689810
rect 111380 689570 111470 689810
rect 111710 689570 111800 689810
rect 112040 689570 112150 689810
rect 112390 689570 112480 689810
rect 112720 689570 112810 689810
rect 113050 689570 113140 689810
rect 113380 689570 113490 689810
rect 113730 689570 113820 689810
rect 114060 689570 114150 689810
rect 114390 689570 114480 689810
rect 114720 689570 114830 689810
rect 115070 689570 115160 689810
rect 115400 689570 115490 689810
rect 115730 689570 115820 689810
rect 116060 689570 116170 689810
rect 116410 689570 116500 689810
rect 116740 689570 116830 689810
rect 117070 689570 117160 689810
rect 117400 689570 117510 689810
rect 117750 689570 117840 689810
rect 118080 689570 118170 689810
rect 118410 689570 118500 689810
rect 118740 689570 118850 689810
rect 119090 689570 119180 689810
rect 119420 689570 119510 689810
rect 119750 689570 119840 689810
rect 120080 689570 120190 689810
rect 120430 689570 120520 689810
rect 120760 689570 120850 689810
rect 121090 689570 121180 689810
rect 121420 689570 121530 689810
rect 121770 689570 121790 689810
rect 110790 689480 121790 689570
rect 110790 689240 110810 689480
rect 111050 689240 111140 689480
rect 111380 689240 111470 689480
rect 111710 689240 111800 689480
rect 112040 689240 112150 689480
rect 112390 689240 112480 689480
rect 112720 689240 112810 689480
rect 113050 689240 113140 689480
rect 113380 689240 113490 689480
rect 113730 689240 113820 689480
rect 114060 689240 114150 689480
rect 114390 689240 114480 689480
rect 114720 689240 114830 689480
rect 115070 689240 115160 689480
rect 115400 689240 115490 689480
rect 115730 689240 115820 689480
rect 116060 689240 116170 689480
rect 116410 689240 116500 689480
rect 116740 689240 116830 689480
rect 117070 689240 117160 689480
rect 117400 689240 117510 689480
rect 117750 689240 117840 689480
rect 118080 689240 118170 689480
rect 118410 689240 118500 689480
rect 118740 689240 118850 689480
rect 119090 689240 119180 689480
rect 119420 689240 119510 689480
rect 119750 689240 119840 689480
rect 120080 689240 120190 689480
rect 120430 689240 120520 689480
rect 120760 689240 120850 689480
rect 121090 689240 121180 689480
rect 121420 689240 121530 689480
rect 121770 689240 121790 689480
rect 110790 689130 121790 689240
rect 110790 688890 110810 689130
rect 111050 688890 111140 689130
rect 111380 688890 111470 689130
rect 111710 688890 111800 689130
rect 112040 688890 112150 689130
rect 112390 688890 112480 689130
rect 112720 688890 112810 689130
rect 113050 688890 113140 689130
rect 113380 688890 113490 689130
rect 113730 688890 113820 689130
rect 114060 688890 114150 689130
rect 114390 688890 114480 689130
rect 114720 688890 114830 689130
rect 115070 688890 115160 689130
rect 115400 688890 115490 689130
rect 115730 688890 115820 689130
rect 116060 688890 116170 689130
rect 116410 688890 116500 689130
rect 116740 688890 116830 689130
rect 117070 688890 117160 689130
rect 117400 688890 117510 689130
rect 117750 688890 117840 689130
rect 118080 688890 118170 689130
rect 118410 688890 118500 689130
rect 118740 688890 118850 689130
rect 119090 688890 119180 689130
rect 119420 688890 119510 689130
rect 119750 688890 119840 689130
rect 120080 688890 120190 689130
rect 120430 688890 120520 689130
rect 120760 688890 120850 689130
rect 121090 688890 121180 689130
rect 121420 688890 121530 689130
rect 121770 688890 121790 689130
rect 110790 688800 121790 688890
rect 110790 688560 110810 688800
rect 111050 688560 111140 688800
rect 111380 688560 111470 688800
rect 111710 688560 111800 688800
rect 112040 688560 112150 688800
rect 112390 688560 112480 688800
rect 112720 688560 112810 688800
rect 113050 688560 113140 688800
rect 113380 688560 113490 688800
rect 113730 688560 113820 688800
rect 114060 688560 114150 688800
rect 114390 688560 114480 688800
rect 114720 688560 114830 688800
rect 115070 688560 115160 688800
rect 115400 688560 115490 688800
rect 115730 688560 115820 688800
rect 116060 688560 116170 688800
rect 116410 688560 116500 688800
rect 116740 688560 116830 688800
rect 117070 688560 117160 688800
rect 117400 688560 117510 688800
rect 117750 688560 117840 688800
rect 118080 688560 118170 688800
rect 118410 688560 118500 688800
rect 118740 688560 118850 688800
rect 119090 688560 119180 688800
rect 119420 688560 119510 688800
rect 119750 688560 119840 688800
rect 120080 688560 120190 688800
rect 120430 688560 120520 688800
rect 120760 688560 120850 688800
rect 121090 688560 121180 688800
rect 121420 688560 121530 688800
rect 121770 688560 121790 688800
rect 110790 688470 121790 688560
rect 110790 688230 110810 688470
rect 111050 688230 111140 688470
rect 111380 688230 111470 688470
rect 111710 688230 111800 688470
rect 112040 688230 112150 688470
rect 112390 688230 112480 688470
rect 112720 688230 112810 688470
rect 113050 688230 113140 688470
rect 113380 688230 113490 688470
rect 113730 688230 113820 688470
rect 114060 688230 114150 688470
rect 114390 688230 114480 688470
rect 114720 688230 114830 688470
rect 115070 688230 115160 688470
rect 115400 688230 115490 688470
rect 115730 688230 115820 688470
rect 116060 688230 116170 688470
rect 116410 688230 116500 688470
rect 116740 688230 116830 688470
rect 117070 688230 117160 688470
rect 117400 688230 117510 688470
rect 117750 688230 117840 688470
rect 118080 688230 118170 688470
rect 118410 688230 118500 688470
rect 118740 688230 118850 688470
rect 119090 688230 119180 688470
rect 119420 688230 119510 688470
rect 119750 688230 119840 688470
rect 120080 688230 120190 688470
rect 120430 688230 120520 688470
rect 120760 688230 120850 688470
rect 121090 688230 121180 688470
rect 121420 688230 121530 688470
rect 121770 688230 121790 688470
rect 110790 688140 121790 688230
rect 110790 687900 110810 688140
rect 111050 687900 111140 688140
rect 111380 687900 111470 688140
rect 111710 687900 111800 688140
rect 112040 687900 112150 688140
rect 112390 687900 112480 688140
rect 112720 687900 112810 688140
rect 113050 687900 113140 688140
rect 113380 687900 113490 688140
rect 113730 687900 113820 688140
rect 114060 687900 114150 688140
rect 114390 687900 114480 688140
rect 114720 687900 114830 688140
rect 115070 687900 115160 688140
rect 115400 687900 115490 688140
rect 115730 687900 115820 688140
rect 116060 687900 116170 688140
rect 116410 687900 116500 688140
rect 116740 687900 116830 688140
rect 117070 687900 117160 688140
rect 117400 687900 117510 688140
rect 117750 687900 117840 688140
rect 118080 687900 118170 688140
rect 118410 687900 118500 688140
rect 118740 687900 118850 688140
rect 119090 687900 119180 688140
rect 119420 687900 119510 688140
rect 119750 687900 119840 688140
rect 120080 687900 120190 688140
rect 120430 687900 120520 688140
rect 120760 687900 120850 688140
rect 121090 687900 121180 688140
rect 121420 687900 121530 688140
rect 121770 687900 121790 688140
rect 110790 687790 121790 687900
rect 110790 687550 110810 687790
rect 111050 687550 111140 687790
rect 111380 687550 111470 687790
rect 111710 687550 111800 687790
rect 112040 687550 112150 687790
rect 112390 687550 112480 687790
rect 112720 687550 112810 687790
rect 113050 687550 113140 687790
rect 113380 687550 113490 687790
rect 113730 687550 113820 687790
rect 114060 687550 114150 687790
rect 114390 687550 114480 687790
rect 114720 687550 114830 687790
rect 115070 687550 115160 687790
rect 115400 687550 115490 687790
rect 115730 687550 115820 687790
rect 116060 687550 116170 687790
rect 116410 687550 116500 687790
rect 116740 687550 116830 687790
rect 117070 687550 117160 687790
rect 117400 687550 117510 687790
rect 117750 687550 117840 687790
rect 118080 687550 118170 687790
rect 118410 687550 118500 687790
rect 118740 687550 118850 687790
rect 119090 687550 119180 687790
rect 119420 687550 119510 687790
rect 119750 687550 119840 687790
rect 120080 687550 120190 687790
rect 120430 687550 120520 687790
rect 120760 687550 120850 687790
rect 121090 687550 121180 687790
rect 121420 687550 121530 687790
rect 121770 687550 121790 687790
rect 110790 687460 121790 687550
rect 110790 687220 110810 687460
rect 111050 687220 111140 687460
rect 111380 687220 111470 687460
rect 111710 687220 111800 687460
rect 112040 687220 112150 687460
rect 112390 687220 112480 687460
rect 112720 687220 112810 687460
rect 113050 687220 113140 687460
rect 113380 687220 113490 687460
rect 113730 687220 113820 687460
rect 114060 687220 114150 687460
rect 114390 687220 114480 687460
rect 114720 687220 114830 687460
rect 115070 687220 115160 687460
rect 115400 687220 115490 687460
rect 115730 687220 115820 687460
rect 116060 687220 116170 687460
rect 116410 687220 116500 687460
rect 116740 687220 116830 687460
rect 117070 687220 117160 687460
rect 117400 687220 117510 687460
rect 117750 687220 117840 687460
rect 118080 687220 118170 687460
rect 118410 687220 118500 687460
rect 118740 687220 118850 687460
rect 119090 687220 119180 687460
rect 119420 687220 119510 687460
rect 119750 687220 119840 687460
rect 120080 687220 120190 687460
rect 120430 687220 120520 687460
rect 120760 687220 120850 687460
rect 121090 687220 121180 687460
rect 121420 687220 121530 687460
rect 121770 687220 121790 687460
rect 110790 687130 121790 687220
rect 110790 686890 110810 687130
rect 111050 686890 111140 687130
rect 111380 686890 111470 687130
rect 111710 686890 111800 687130
rect 112040 686890 112150 687130
rect 112390 686890 112480 687130
rect 112720 686890 112810 687130
rect 113050 686890 113140 687130
rect 113380 686890 113490 687130
rect 113730 686890 113820 687130
rect 114060 686890 114150 687130
rect 114390 686890 114480 687130
rect 114720 686890 114830 687130
rect 115070 686890 115160 687130
rect 115400 686890 115490 687130
rect 115730 686890 115820 687130
rect 116060 686890 116170 687130
rect 116410 686890 116500 687130
rect 116740 686890 116830 687130
rect 117070 686890 117160 687130
rect 117400 686890 117510 687130
rect 117750 686890 117840 687130
rect 118080 686890 118170 687130
rect 118410 686890 118500 687130
rect 118740 686890 118850 687130
rect 119090 686890 119180 687130
rect 119420 686890 119510 687130
rect 119750 686890 119840 687130
rect 120080 686890 120190 687130
rect 120430 686890 120520 687130
rect 120760 686890 120850 687130
rect 121090 686890 121180 687130
rect 121420 686890 121530 687130
rect 121770 686890 121790 687130
rect 110790 686800 121790 686890
rect 110790 686560 110810 686800
rect 111050 686560 111140 686800
rect 111380 686560 111470 686800
rect 111710 686560 111800 686800
rect 112040 686560 112150 686800
rect 112390 686560 112480 686800
rect 112720 686560 112810 686800
rect 113050 686560 113140 686800
rect 113380 686560 113490 686800
rect 113730 686560 113820 686800
rect 114060 686560 114150 686800
rect 114390 686560 114480 686800
rect 114720 686560 114830 686800
rect 115070 686560 115160 686800
rect 115400 686560 115490 686800
rect 115730 686560 115820 686800
rect 116060 686560 116170 686800
rect 116410 686560 116500 686800
rect 116740 686560 116830 686800
rect 117070 686560 117160 686800
rect 117400 686560 117510 686800
rect 117750 686560 117840 686800
rect 118080 686560 118170 686800
rect 118410 686560 118500 686800
rect 118740 686560 118850 686800
rect 119090 686560 119180 686800
rect 119420 686560 119510 686800
rect 119750 686560 119840 686800
rect 120080 686560 120190 686800
rect 120430 686560 120520 686800
rect 120760 686560 120850 686800
rect 121090 686560 121180 686800
rect 121420 686560 121530 686800
rect 121770 686560 121790 686800
rect 110790 686450 121790 686560
rect 110790 686210 110810 686450
rect 111050 686210 111140 686450
rect 111380 686210 111470 686450
rect 111710 686210 111800 686450
rect 112040 686210 112150 686450
rect 112390 686210 112480 686450
rect 112720 686210 112810 686450
rect 113050 686210 113140 686450
rect 113380 686210 113490 686450
rect 113730 686210 113820 686450
rect 114060 686210 114150 686450
rect 114390 686210 114480 686450
rect 114720 686210 114830 686450
rect 115070 686210 115160 686450
rect 115400 686210 115490 686450
rect 115730 686210 115820 686450
rect 116060 686210 116170 686450
rect 116410 686210 116500 686450
rect 116740 686210 116830 686450
rect 117070 686210 117160 686450
rect 117400 686210 117510 686450
rect 117750 686210 117840 686450
rect 118080 686210 118170 686450
rect 118410 686210 118500 686450
rect 118740 686210 118850 686450
rect 119090 686210 119180 686450
rect 119420 686210 119510 686450
rect 119750 686210 119840 686450
rect 120080 686210 120190 686450
rect 120430 686210 120520 686450
rect 120760 686210 120850 686450
rect 121090 686210 121180 686450
rect 121420 686210 121530 686450
rect 121770 686210 121790 686450
rect 110790 686120 121790 686210
rect 110790 685880 110810 686120
rect 111050 685880 111140 686120
rect 111380 685880 111470 686120
rect 111710 685880 111800 686120
rect 112040 685880 112150 686120
rect 112390 685880 112480 686120
rect 112720 685880 112810 686120
rect 113050 685880 113140 686120
rect 113380 685880 113490 686120
rect 113730 685880 113820 686120
rect 114060 685880 114150 686120
rect 114390 685880 114480 686120
rect 114720 685880 114830 686120
rect 115070 685880 115160 686120
rect 115400 685880 115490 686120
rect 115730 685880 115820 686120
rect 116060 685880 116170 686120
rect 116410 685880 116500 686120
rect 116740 685880 116830 686120
rect 117070 685880 117160 686120
rect 117400 685880 117510 686120
rect 117750 685880 117840 686120
rect 118080 685880 118170 686120
rect 118410 685880 118500 686120
rect 118740 685880 118850 686120
rect 119090 685880 119180 686120
rect 119420 685880 119510 686120
rect 119750 685880 119840 686120
rect 120080 685880 120190 686120
rect 120430 685880 120520 686120
rect 120760 685880 120850 686120
rect 121090 685880 121180 686120
rect 121420 685880 121530 686120
rect 121770 685880 121790 686120
rect 110790 685790 121790 685880
rect 110790 685550 110810 685790
rect 111050 685550 111140 685790
rect 111380 685550 111470 685790
rect 111710 685550 111800 685790
rect 112040 685550 112150 685790
rect 112390 685550 112480 685790
rect 112720 685550 112810 685790
rect 113050 685550 113140 685790
rect 113380 685550 113490 685790
rect 113730 685550 113820 685790
rect 114060 685550 114150 685790
rect 114390 685550 114480 685790
rect 114720 685550 114830 685790
rect 115070 685550 115160 685790
rect 115400 685550 115490 685790
rect 115730 685550 115820 685790
rect 116060 685550 116170 685790
rect 116410 685550 116500 685790
rect 116740 685550 116830 685790
rect 117070 685550 117160 685790
rect 117400 685550 117510 685790
rect 117750 685550 117840 685790
rect 118080 685550 118170 685790
rect 118410 685550 118500 685790
rect 118740 685550 118850 685790
rect 119090 685550 119180 685790
rect 119420 685550 119510 685790
rect 119750 685550 119840 685790
rect 120080 685550 120190 685790
rect 120430 685550 120520 685790
rect 120760 685550 120850 685790
rect 121090 685550 121180 685790
rect 121420 685550 121530 685790
rect 121770 685550 121790 685790
rect 110790 685460 121790 685550
rect 110790 685220 110810 685460
rect 111050 685220 111140 685460
rect 111380 685220 111470 685460
rect 111710 685220 111800 685460
rect 112040 685220 112150 685460
rect 112390 685220 112480 685460
rect 112720 685220 112810 685460
rect 113050 685220 113140 685460
rect 113380 685220 113490 685460
rect 113730 685220 113820 685460
rect 114060 685220 114150 685460
rect 114390 685220 114480 685460
rect 114720 685220 114830 685460
rect 115070 685220 115160 685460
rect 115400 685220 115490 685460
rect 115730 685220 115820 685460
rect 116060 685220 116170 685460
rect 116410 685220 116500 685460
rect 116740 685220 116830 685460
rect 117070 685220 117160 685460
rect 117400 685220 117510 685460
rect 117750 685220 117840 685460
rect 118080 685220 118170 685460
rect 118410 685220 118500 685460
rect 118740 685220 118850 685460
rect 119090 685220 119180 685460
rect 119420 685220 119510 685460
rect 119750 685220 119840 685460
rect 120080 685220 120190 685460
rect 120430 685220 120520 685460
rect 120760 685220 120850 685460
rect 121090 685220 121180 685460
rect 121420 685220 121530 685460
rect 121770 685220 121790 685460
rect 110790 685110 121790 685220
rect 110790 684870 110810 685110
rect 111050 684870 111140 685110
rect 111380 684870 111470 685110
rect 111710 684870 111800 685110
rect 112040 684870 112150 685110
rect 112390 684870 112480 685110
rect 112720 684870 112810 685110
rect 113050 684870 113140 685110
rect 113380 684870 113490 685110
rect 113730 684870 113820 685110
rect 114060 684870 114150 685110
rect 114390 684870 114480 685110
rect 114720 684870 114830 685110
rect 115070 684870 115160 685110
rect 115400 684870 115490 685110
rect 115730 684870 115820 685110
rect 116060 684870 116170 685110
rect 116410 684870 116500 685110
rect 116740 684870 116830 685110
rect 117070 684870 117160 685110
rect 117400 684870 117510 685110
rect 117750 684870 117840 685110
rect 118080 684870 118170 685110
rect 118410 684870 118500 685110
rect 118740 684870 118850 685110
rect 119090 684870 119180 685110
rect 119420 684870 119510 685110
rect 119750 684870 119840 685110
rect 120080 684870 120190 685110
rect 120430 684870 120520 685110
rect 120760 684870 120850 685110
rect 121090 684870 121180 685110
rect 121420 684870 121530 685110
rect 121770 684870 121790 685110
rect 110790 684780 121790 684870
rect 110790 684540 110810 684780
rect 111050 684540 111140 684780
rect 111380 684540 111470 684780
rect 111710 684540 111800 684780
rect 112040 684540 112150 684780
rect 112390 684540 112480 684780
rect 112720 684540 112810 684780
rect 113050 684540 113140 684780
rect 113380 684540 113490 684780
rect 113730 684540 113820 684780
rect 114060 684540 114150 684780
rect 114390 684540 114480 684780
rect 114720 684540 114830 684780
rect 115070 684540 115160 684780
rect 115400 684540 115490 684780
rect 115730 684540 115820 684780
rect 116060 684540 116170 684780
rect 116410 684540 116500 684780
rect 116740 684540 116830 684780
rect 117070 684540 117160 684780
rect 117400 684540 117510 684780
rect 117750 684540 117840 684780
rect 118080 684540 118170 684780
rect 118410 684540 118500 684780
rect 118740 684540 118850 684780
rect 119090 684540 119180 684780
rect 119420 684540 119510 684780
rect 119750 684540 119840 684780
rect 120080 684540 120190 684780
rect 120430 684540 120520 684780
rect 120760 684540 120850 684780
rect 121090 684540 121180 684780
rect 121420 684540 121530 684780
rect 121770 684540 121790 684780
rect 110790 684450 121790 684540
rect 110790 684210 110810 684450
rect 111050 684210 111140 684450
rect 111380 684210 111470 684450
rect 111710 684210 111800 684450
rect 112040 684210 112150 684450
rect 112390 684210 112480 684450
rect 112720 684210 112810 684450
rect 113050 684210 113140 684450
rect 113380 684210 113490 684450
rect 113730 684210 113820 684450
rect 114060 684210 114150 684450
rect 114390 684210 114480 684450
rect 114720 684210 114830 684450
rect 115070 684210 115160 684450
rect 115400 684210 115490 684450
rect 115730 684210 115820 684450
rect 116060 684210 116170 684450
rect 116410 684210 116500 684450
rect 116740 684210 116830 684450
rect 117070 684210 117160 684450
rect 117400 684210 117510 684450
rect 117750 684210 117840 684450
rect 118080 684210 118170 684450
rect 118410 684210 118500 684450
rect 118740 684210 118850 684450
rect 119090 684210 119180 684450
rect 119420 684210 119510 684450
rect 119750 684210 119840 684450
rect 120080 684210 120190 684450
rect 120430 684210 120520 684450
rect 120760 684210 120850 684450
rect 121090 684210 121180 684450
rect 121420 684210 121530 684450
rect 121770 684210 121790 684450
rect 110790 684120 121790 684210
rect 110790 683880 110810 684120
rect 111050 683880 111140 684120
rect 111380 683880 111470 684120
rect 111710 683880 111800 684120
rect 112040 683880 112150 684120
rect 112390 683880 112480 684120
rect 112720 683880 112810 684120
rect 113050 683880 113140 684120
rect 113380 683880 113490 684120
rect 113730 683880 113820 684120
rect 114060 683880 114150 684120
rect 114390 683880 114480 684120
rect 114720 683880 114830 684120
rect 115070 683880 115160 684120
rect 115400 683880 115490 684120
rect 115730 683880 115820 684120
rect 116060 683880 116170 684120
rect 116410 683880 116500 684120
rect 116740 683880 116830 684120
rect 117070 683880 117160 684120
rect 117400 683880 117510 684120
rect 117750 683880 117840 684120
rect 118080 683880 118170 684120
rect 118410 683880 118500 684120
rect 118740 683880 118850 684120
rect 119090 683880 119180 684120
rect 119420 683880 119510 684120
rect 119750 683880 119840 684120
rect 120080 683880 120190 684120
rect 120430 683880 120520 684120
rect 120760 683880 120850 684120
rect 121090 683880 121180 684120
rect 121420 683880 121530 684120
rect 121770 683880 121790 684120
rect 110790 683860 121790 683880
rect 122170 694840 133170 694860
rect 122170 694600 122190 694840
rect 122430 694600 122520 694840
rect 122760 694600 122850 694840
rect 123090 694600 123180 694840
rect 123420 694600 123530 694840
rect 123770 694600 123860 694840
rect 124100 694600 124190 694840
rect 124430 694600 124520 694840
rect 124760 694600 124870 694840
rect 125110 694600 125200 694840
rect 125440 694600 125530 694840
rect 125770 694600 125860 694840
rect 126100 694600 126210 694840
rect 126450 694600 126540 694840
rect 126780 694600 126870 694840
rect 127110 694600 127200 694840
rect 127440 694600 127550 694840
rect 127790 694600 127880 694840
rect 128120 694600 128210 694840
rect 128450 694600 128540 694840
rect 128780 694600 128890 694840
rect 129130 694600 129220 694840
rect 129460 694600 129550 694840
rect 129790 694600 129880 694840
rect 130120 694600 130230 694840
rect 130470 694600 130560 694840
rect 130800 694600 130890 694840
rect 131130 694600 131220 694840
rect 131460 694600 131570 694840
rect 131810 694600 131900 694840
rect 132140 694600 132230 694840
rect 132470 694600 132560 694840
rect 132800 694600 132910 694840
rect 133150 694600 133170 694840
rect 122170 694490 133170 694600
rect 122170 694250 122190 694490
rect 122430 694250 122520 694490
rect 122760 694250 122850 694490
rect 123090 694250 123180 694490
rect 123420 694250 123530 694490
rect 123770 694250 123860 694490
rect 124100 694250 124190 694490
rect 124430 694250 124520 694490
rect 124760 694250 124870 694490
rect 125110 694250 125200 694490
rect 125440 694250 125530 694490
rect 125770 694250 125860 694490
rect 126100 694250 126210 694490
rect 126450 694250 126540 694490
rect 126780 694250 126870 694490
rect 127110 694250 127200 694490
rect 127440 694250 127550 694490
rect 127790 694250 127880 694490
rect 128120 694250 128210 694490
rect 128450 694250 128540 694490
rect 128780 694250 128890 694490
rect 129130 694250 129220 694490
rect 129460 694250 129550 694490
rect 129790 694250 129880 694490
rect 130120 694250 130230 694490
rect 130470 694250 130560 694490
rect 130800 694250 130890 694490
rect 131130 694250 131220 694490
rect 131460 694250 131570 694490
rect 131810 694250 131900 694490
rect 132140 694250 132230 694490
rect 132470 694250 132560 694490
rect 132800 694250 132910 694490
rect 133150 694250 133170 694490
rect 122170 694160 133170 694250
rect 122170 693920 122190 694160
rect 122430 693920 122520 694160
rect 122760 693920 122850 694160
rect 123090 693920 123180 694160
rect 123420 693920 123530 694160
rect 123770 693920 123860 694160
rect 124100 693920 124190 694160
rect 124430 693920 124520 694160
rect 124760 693920 124870 694160
rect 125110 693920 125200 694160
rect 125440 693920 125530 694160
rect 125770 693920 125860 694160
rect 126100 693920 126210 694160
rect 126450 693920 126540 694160
rect 126780 693920 126870 694160
rect 127110 693920 127200 694160
rect 127440 693920 127550 694160
rect 127790 693920 127880 694160
rect 128120 693920 128210 694160
rect 128450 693920 128540 694160
rect 128780 693920 128890 694160
rect 129130 693920 129220 694160
rect 129460 693920 129550 694160
rect 129790 693920 129880 694160
rect 130120 693920 130230 694160
rect 130470 693920 130560 694160
rect 130800 693920 130890 694160
rect 131130 693920 131220 694160
rect 131460 693920 131570 694160
rect 131810 693920 131900 694160
rect 132140 693920 132230 694160
rect 132470 693920 132560 694160
rect 132800 693920 132910 694160
rect 133150 693920 133170 694160
rect 122170 693830 133170 693920
rect 122170 693590 122190 693830
rect 122430 693590 122520 693830
rect 122760 693590 122850 693830
rect 123090 693590 123180 693830
rect 123420 693590 123530 693830
rect 123770 693590 123860 693830
rect 124100 693590 124190 693830
rect 124430 693590 124520 693830
rect 124760 693590 124870 693830
rect 125110 693590 125200 693830
rect 125440 693590 125530 693830
rect 125770 693590 125860 693830
rect 126100 693590 126210 693830
rect 126450 693590 126540 693830
rect 126780 693590 126870 693830
rect 127110 693590 127200 693830
rect 127440 693590 127550 693830
rect 127790 693590 127880 693830
rect 128120 693590 128210 693830
rect 128450 693590 128540 693830
rect 128780 693590 128890 693830
rect 129130 693590 129220 693830
rect 129460 693590 129550 693830
rect 129790 693590 129880 693830
rect 130120 693590 130230 693830
rect 130470 693590 130560 693830
rect 130800 693590 130890 693830
rect 131130 693590 131220 693830
rect 131460 693590 131570 693830
rect 131810 693590 131900 693830
rect 132140 693590 132230 693830
rect 132470 693590 132560 693830
rect 132800 693590 132910 693830
rect 133150 693590 133170 693830
rect 122170 693500 133170 693590
rect 122170 693260 122190 693500
rect 122430 693260 122520 693500
rect 122760 693260 122850 693500
rect 123090 693260 123180 693500
rect 123420 693260 123530 693500
rect 123770 693260 123860 693500
rect 124100 693260 124190 693500
rect 124430 693260 124520 693500
rect 124760 693260 124870 693500
rect 125110 693260 125200 693500
rect 125440 693260 125530 693500
rect 125770 693260 125860 693500
rect 126100 693260 126210 693500
rect 126450 693260 126540 693500
rect 126780 693260 126870 693500
rect 127110 693260 127200 693500
rect 127440 693260 127550 693500
rect 127790 693260 127880 693500
rect 128120 693260 128210 693500
rect 128450 693260 128540 693500
rect 128780 693260 128890 693500
rect 129130 693260 129220 693500
rect 129460 693260 129550 693500
rect 129790 693260 129880 693500
rect 130120 693260 130230 693500
rect 130470 693260 130560 693500
rect 130800 693260 130890 693500
rect 131130 693260 131220 693500
rect 131460 693260 131570 693500
rect 131810 693260 131900 693500
rect 132140 693260 132230 693500
rect 132470 693260 132560 693500
rect 132800 693260 132910 693500
rect 133150 693260 133170 693500
rect 122170 693150 133170 693260
rect 122170 692910 122190 693150
rect 122430 692910 122520 693150
rect 122760 692910 122850 693150
rect 123090 692910 123180 693150
rect 123420 692910 123530 693150
rect 123770 692910 123860 693150
rect 124100 692910 124190 693150
rect 124430 692910 124520 693150
rect 124760 692910 124870 693150
rect 125110 692910 125200 693150
rect 125440 692910 125530 693150
rect 125770 692910 125860 693150
rect 126100 692910 126210 693150
rect 126450 692910 126540 693150
rect 126780 692910 126870 693150
rect 127110 692910 127200 693150
rect 127440 692910 127550 693150
rect 127790 692910 127880 693150
rect 128120 692910 128210 693150
rect 128450 692910 128540 693150
rect 128780 692910 128890 693150
rect 129130 692910 129220 693150
rect 129460 692910 129550 693150
rect 129790 692910 129880 693150
rect 130120 692910 130230 693150
rect 130470 692910 130560 693150
rect 130800 692910 130890 693150
rect 131130 692910 131220 693150
rect 131460 692910 131570 693150
rect 131810 692910 131900 693150
rect 132140 692910 132230 693150
rect 132470 692910 132560 693150
rect 132800 692910 132910 693150
rect 133150 692910 133170 693150
rect 122170 692820 133170 692910
rect 122170 692580 122190 692820
rect 122430 692580 122520 692820
rect 122760 692580 122850 692820
rect 123090 692580 123180 692820
rect 123420 692580 123530 692820
rect 123770 692580 123860 692820
rect 124100 692580 124190 692820
rect 124430 692580 124520 692820
rect 124760 692580 124870 692820
rect 125110 692580 125200 692820
rect 125440 692580 125530 692820
rect 125770 692580 125860 692820
rect 126100 692580 126210 692820
rect 126450 692580 126540 692820
rect 126780 692580 126870 692820
rect 127110 692580 127200 692820
rect 127440 692580 127550 692820
rect 127790 692580 127880 692820
rect 128120 692580 128210 692820
rect 128450 692580 128540 692820
rect 128780 692580 128890 692820
rect 129130 692580 129220 692820
rect 129460 692580 129550 692820
rect 129790 692580 129880 692820
rect 130120 692580 130230 692820
rect 130470 692580 130560 692820
rect 130800 692580 130890 692820
rect 131130 692580 131220 692820
rect 131460 692580 131570 692820
rect 131810 692580 131900 692820
rect 132140 692580 132230 692820
rect 132470 692580 132560 692820
rect 132800 692580 132910 692820
rect 133150 692580 133170 692820
rect 122170 692490 133170 692580
rect 122170 692250 122190 692490
rect 122430 692250 122520 692490
rect 122760 692250 122850 692490
rect 123090 692250 123180 692490
rect 123420 692250 123530 692490
rect 123770 692250 123860 692490
rect 124100 692250 124190 692490
rect 124430 692250 124520 692490
rect 124760 692250 124870 692490
rect 125110 692250 125200 692490
rect 125440 692250 125530 692490
rect 125770 692250 125860 692490
rect 126100 692250 126210 692490
rect 126450 692250 126540 692490
rect 126780 692250 126870 692490
rect 127110 692250 127200 692490
rect 127440 692250 127550 692490
rect 127790 692250 127880 692490
rect 128120 692250 128210 692490
rect 128450 692250 128540 692490
rect 128780 692250 128890 692490
rect 129130 692250 129220 692490
rect 129460 692250 129550 692490
rect 129790 692250 129880 692490
rect 130120 692250 130230 692490
rect 130470 692250 130560 692490
rect 130800 692250 130890 692490
rect 131130 692250 131220 692490
rect 131460 692250 131570 692490
rect 131810 692250 131900 692490
rect 132140 692250 132230 692490
rect 132470 692250 132560 692490
rect 132800 692250 132910 692490
rect 133150 692250 133170 692490
rect 122170 692160 133170 692250
rect 122170 691920 122190 692160
rect 122430 691920 122520 692160
rect 122760 691920 122850 692160
rect 123090 691920 123180 692160
rect 123420 691920 123530 692160
rect 123770 691920 123860 692160
rect 124100 691920 124190 692160
rect 124430 691920 124520 692160
rect 124760 691920 124870 692160
rect 125110 691920 125200 692160
rect 125440 691920 125530 692160
rect 125770 691920 125860 692160
rect 126100 691920 126210 692160
rect 126450 691920 126540 692160
rect 126780 691920 126870 692160
rect 127110 691920 127200 692160
rect 127440 691920 127550 692160
rect 127790 691920 127880 692160
rect 128120 691920 128210 692160
rect 128450 691920 128540 692160
rect 128780 691920 128890 692160
rect 129130 691920 129220 692160
rect 129460 691920 129550 692160
rect 129790 691920 129880 692160
rect 130120 691920 130230 692160
rect 130470 691920 130560 692160
rect 130800 691920 130890 692160
rect 131130 691920 131220 692160
rect 131460 691920 131570 692160
rect 131810 691920 131900 692160
rect 132140 691920 132230 692160
rect 132470 691920 132560 692160
rect 132800 691920 132910 692160
rect 133150 691920 133170 692160
rect 122170 691810 133170 691920
rect 122170 691570 122190 691810
rect 122430 691570 122520 691810
rect 122760 691570 122850 691810
rect 123090 691570 123180 691810
rect 123420 691570 123530 691810
rect 123770 691570 123860 691810
rect 124100 691570 124190 691810
rect 124430 691570 124520 691810
rect 124760 691570 124870 691810
rect 125110 691570 125200 691810
rect 125440 691570 125530 691810
rect 125770 691570 125860 691810
rect 126100 691570 126210 691810
rect 126450 691570 126540 691810
rect 126780 691570 126870 691810
rect 127110 691570 127200 691810
rect 127440 691570 127550 691810
rect 127790 691570 127880 691810
rect 128120 691570 128210 691810
rect 128450 691570 128540 691810
rect 128780 691570 128890 691810
rect 129130 691570 129220 691810
rect 129460 691570 129550 691810
rect 129790 691570 129880 691810
rect 130120 691570 130230 691810
rect 130470 691570 130560 691810
rect 130800 691570 130890 691810
rect 131130 691570 131220 691810
rect 131460 691570 131570 691810
rect 131810 691570 131900 691810
rect 132140 691570 132230 691810
rect 132470 691570 132560 691810
rect 132800 691570 132910 691810
rect 133150 691570 133170 691810
rect 122170 691480 133170 691570
rect 122170 691240 122190 691480
rect 122430 691240 122520 691480
rect 122760 691240 122850 691480
rect 123090 691240 123180 691480
rect 123420 691240 123530 691480
rect 123770 691240 123860 691480
rect 124100 691240 124190 691480
rect 124430 691240 124520 691480
rect 124760 691240 124870 691480
rect 125110 691240 125200 691480
rect 125440 691240 125530 691480
rect 125770 691240 125860 691480
rect 126100 691240 126210 691480
rect 126450 691240 126540 691480
rect 126780 691240 126870 691480
rect 127110 691240 127200 691480
rect 127440 691240 127550 691480
rect 127790 691240 127880 691480
rect 128120 691240 128210 691480
rect 128450 691240 128540 691480
rect 128780 691240 128890 691480
rect 129130 691240 129220 691480
rect 129460 691240 129550 691480
rect 129790 691240 129880 691480
rect 130120 691240 130230 691480
rect 130470 691240 130560 691480
rect 130800 691240 130890 691480
rect 131130 691240 131220 691480
rect 131460 691240 131570 691480
rect 131810 691240 131900 691480
rect 132140 691240 132230 691480
rect 132470 691240 132560 691480
rect 132800 691240 132910 691480
rect 133150 691240 133170 691480
rect 122170 691150 133170 691240
rect 122170 690910 122190 691150
rect 122430 690910 122520 691150
rect 122760 690910 122850 691150
rect 123090 690910 123180 691150
rect 123420 690910 123530 691150
rect 123770 690910 123860 691150
rect 124100 690910 124190 691150
rect 124430 690910 124520 691150
rect 124760 690910 124870 691150
rect 125110 690910 125200 691150
rect 125440 690910 125530 691150
rect 125770 690910 125860 691150
rect 126100 690910 126210 691150
rect 126450 690910 126540 691150
rect 126780 690910 126870 691150
rect 127110 690910 127200 691150
rect 127440 690910 127550 691150
rect 127790 690910 127880 691150
rect 128120 690910 128210 691150
rect 128450 690910 128540 691150
rect 128780 690910 128890 691150
rect 129130 690910 129220 691150
rect 129460 690910 129550 691150
rect 129790 690910 129880 691150
rect 130120 690910 130230 691150
rect 130470 690910 130560 691150
rect 130800 690910 130890 691150
rect 131130 690910 131220 691150
rect 131460 690910 131570 691150
rect 131810 690910 131900 691150
rect 132140 690910 132230 691150
rect 132470 690910 132560 691150
rect 132800 690910 132910 691150
rect 133150 690910 133170 691150
rect 122170 690820 133170 690910
rect 122170 690580 122190 690820
rect 122430 690580 122520 690820
rect 122760 690580 122850 690820
rect 123090 690580 123180 690820
rect 123420 690580 123530 690820
rect 123770 690580 123860 690820
rect 124100 690580 124190 690820
rect 124430 690580 124520 690820
rect 124760 690580 124870 690820
rect 125110 690580 125200 690820
rect 125440 690580 125530 690820
rect 125770 690580 125860 690820
rect 126100 690580 126210 690820
rect 126450 690580 126540 690820
rect 126780 690580 126870 690820
rect 127110 690580 127200 690820
rect 127440 690580 127550 690820
rect 127790 690580 127880 690820
rect 128120 690580 128210 690820
rect 128450 690580 128540 690820
rect 128780 690580 128890 690820
rect 129130 690580 129220 690820
rect 129460 690580 129550 690820
rect 129790 690580 129880 690820
rect 130120 690580 130230 690820
rect 130470 690580 130560 690820
rect 130800 690580 130890 690820
rect 131130 690580 131220 690820
rect 131460 690580 131570 690820
rect 131810 690580 131900 690820
rect 132140 690580 132230 690820
rect 132470 690580 132560 690820
rect 132800 690580 132910 690820
rect 133150 690580 133170 690820
rect 122170 690470 133170 690580
rect 122170 690230 122190 690470
rect 122430 690230 122520 690470
rect 122760 690230 122850 690470
rect 123090 690230 123180 690470
rect 123420 690230 123530 690470
rect 123770 690230 123860 690470
rect 124100 690230 124190 690470
rect 124430 690230 124520 690470
rect 124760 690230 124870 690470
rect 125110 690230 125200 690470
rect 125440 690230 125530 690470
rect 125770 690230 125860 690470
rect 126100 690230 126210 690470
rect 126450 690230 126540 690470
rect 126780 690230 126870 690470
rect 127110 690230 127200 690470
rect 127440 690230 127550 690470
rect 127790 690230 127880 690470
rect 128120 690230 128210 690470
rect 128450 690230 128540 690470
rect 128780 690230 128890 690470
rect 129130 690230 129220 690470
rect 129460 690230 129550 690470
rect 129790 690230 129880 690470
rect 130120 690230 130230 690470
rect 130470 690230 130560 690470
rect 130800 690230 130890 690470
rect 131130 690230 131220 690470
rect 131460 690230 131570 690470
rect 131810 690230 131900 690470
rect 132140 690230 132230 690470
rect 132470 690230 132560 690470
rect 132800 690230 132910 690470
rect 133150 690230 133170 690470
rect 122170 690140 133170 690230
rect 122170 689900 122190 690140
rect 122430 689900 122520 690140
rect 122760 689900 122850 690140
rect 123090 689900 123180 690140
rect 123420 689900 123530 690140
rect 123770 689900 123860 690140
rect 124100 689900 124190 690140
rect 124430 689900 124520 690140
rect 124760 689900 124870 690140
rect 125110 689900 125200 690140
rect 125440 689900 125530 690140
rect 125770 689900 125860 690140
rect 126100 689900 126210 690140
rect 126450 689900 126540 690140
rect 126780 689900 126870 690140
rect 127110 689900 127200 690140
rect 127440 689900 127550 690140
rect 127790 689900 127880 690140
rect 128120 689900 128210 690140
rect 128450 689900 128540 690140
rect 128780 689900 128890 690140
rect 129130 689900 129220 690140
rect 129460 689900 129550 690140
rect 129790 689900 129880 690140
rect 130120 689900 130230 690140
rect 130470 689900 130560 690140
rect 130800 689900 130890 690140
rect 131130 689900 131220 690140
rect 131460 689900 131570 690140
rect 131810 689900 131900 690140
rect 132140 689900 132230 690140
rect 132470 689900 132560 690140
rect 132800 689900 132910 690140
rect 133150 689900 133170 690140
rect 122170 689810 133170 689900
rect 122170 689570 122190 689810
rect 122430 689570 122520 689810
rect 122760 689570 122850 689810
rect 123090 689570 123180 689810
rect 123420 689570 123530 689810
rect 123770 689570 123860 689810
rect 124100 689570 124190 689810
rect 124430 689570 124520 689810
rect 124760 689570 124870 689810
rect 125110 689570 125200 689810
rect 125440 689570 125530 689810
rect 125770 689570 125860 689810
rect 126100 689570 126210 689810
rect 126450 689570 126540 689810
rect 126780 689570 126870 689810
rect 127110 689570 127200 689810
rect 127440 689570 127550 689810
rect 127790 689570 127880 689810
rect 128120 689570 128210 689810
rect 128450 689570 128540 689810
rect 128780 689570 128890 689810
rect 129130 689570 129220 689810
rect 129460 689570 129550 689810
rect 129790 689570 129880 689810
rect 130120 689570 130230 689810
rect 130470 689570 130560 689810
rect 130800 689570 130890 689810
rect 131130 689570 131220 689810
rect 131460 689570 131570 689810
rect 131810 689570 131900 689810
rect 132140 689570 132230 689810
rect 132470 689570 132560 689810
rect 132800 689570 132910 689810
rect 133150 689570 133170 689810
rect 122170 689480 133170 689570
rect 122170 689240 122190 689480
rect 122430 689240 122520 689480
rect 122760 689240 122850 689480
rect 123090 689240 123180 689480
rect 123420 689240 123530 689480
rect 123770 689240 123860 689480
rect 124100 689240 124190 689480
rect 124430 689240 124520 689480
rect 124760 689240 124870 689480
rect 125110 689240 125200 689480
rect 125440 689240 125530 689480
rect 125770 689240 125860 689480
rect 126100 689240 126210 689480
rect 126450 689240 126540 689480
rect 126780 689240 126870 689480
rect 127110 689240 127200 689480
rect 127440 689240 127550 689480
rect 127790 689240 127880 689480
rect 128120 689240 128210 689480
rect 128450 689240 128540 689480
rect 128780 689240 128890 689480
rect 129130 689240 129220 689480
rect 129460 689240 129550 689480
rect 129790 689240 129880 689480
rect 130120 689240 130230 689480
rect 130470 689240 130560 689480
rect 130800 689240 130890 689480
rect 131130 689240 131220 689480
rect 131460 689240 131570 689480
rect 131810 689240 131900 689480
rect 132140 689240 132230 689480
rect 132470 689240 132560 689480
rect 132800 689240 132910 689480
rect 133150 689240 133170 689480
rect 122170 689130 133170 689240
rect 122170 688890 122190 689130
rect 122430 688890 122520 689130
rect 122760 688890 122850 689130
rect 123090 688890 123180 689130
rect 123420 688890 123530 689130
rect 123770 688890 123860 689130
rect 124100 688890 124190 689130
rect 124430 688890 124520 689130
rect 124760 688890 124870 689130
rect 125110 688890 125200 689130
rect 125440 688890 125530 689130
rect 125770 688890 125860 689130
rect 126100 688890 126210 689130
rect 126450 688890 126540 689130
rect 126780 688890 126870 689130
rect 127110 688890 127200 689130
rect 127440 688890 127550 689130
rect 127790 688890 127880 689130
rect 128120 688890 128210 689130
rect 128450 688890 128540 689130
rect 128780 688890 128890 689130
rect 129130 688890 129220 689130
rect 129460 688890 129550 689130
rect 129790 688890 129880 689130
rect 130120 688890 130230 689130
rect 130470 688890 130560 689130
rect 130800 688890 130890 689130
rect 131130 688890 131220 689130
rect 131460 688890 131570 689130
rect 131810 688890 131900 689130
rect 132140 688890 132230 689130
rect 132470 688890 132560 689130
rect 132800 688890 132910 689130
rect 133150 688890 133170 689130
rect 122170 688800 133170 688890
rect 122170 688560 122190 688800
rect 122430 688560 122520 688800
rect 122760 688560 122850 688800
rect 123090 688560 123180 688800
rect 123420 688560 123530 688800
rect 123770 688560 123860 688800
rect 124100 688560 124190 688800
rect 124430 688560 124520 688800
rect 124760 688560 124870 688800
rect 125110 688560 125200 688800
rect 125440 688560 125530 688800
rect 125770 688560 125860 688800
rect 126100 688560 126210 688800
rect 126450 688560 126540 688800
rect 126780 688560 126870 688800
rect 127110 688560 127200 688800
rect 127440 688560 127550 688800
rect 127790 688560 127880 688800
rect 128120 688560 128210 688800
rect 128450 688560 128540 688800
rect 128780 688560 128890 688800
rect 129130 688560 129220 688800
rect 129460 688560 129550 688800
rect 129790 688560 129880 688800
rect 130120 688560 130230 688800
rect 130470 688560 130560 688800
rect 130800 688560 130890 688800
rect 131130 688560 131220 688800
rect 131460 688560 131570 688800
rect 131810 688560 131900 688800
rect 132140 688560 132230 688800
rect 132470 688560 132560 688800
rect 132800 688560 132910 688800
rect 133150 688560 133170 688800
rect 122170 688470 133170 688560
rect 122170 688230 122190 688470
rect 122430 688230 122520 688470
rect 122760 688230 122850 688470
rect 123090 688230 123180 688470
rect 123420 688230 123530 688470
rect 123770 688230 123860 688470
rect 124100 688230 124190 688470
rect 124430 688230 124520 688470
rect 124760 688230 124870 688470
rect 125110 688230 125200 688470
rect 125440 688230 125530 688470
rect 125770 688230 125860 688470
rect 126100 688230 126210 688470
rect 126450 688230 126540 688470
rect 126780 688230 126870 688470
rect 127110 688230 127200 688470
rect 127440 688230 127550 688470
rect 127790 688230 127880 688470
rect 128120 688230 128210 688470
rect 128450 688230 128540 688470
rect 128780 688230 128890 688470
rect 129130 688230 129220 688470
rect 129460 688230 129550 688470
rect 129790 688230 129880 688470
rect 130120 688230 130230 688470
rect 130470 688230 130560 688470
rect 130800 688230 130890 688470
rect 131130 688230 131220 688470
rect 131460 688230 131570 688470
rect 131810 688230 131900 688470
rect 132140 688230 132230 688470
rect 132470 688230 132560 688470
rect 132800 688230 132910 688470
rect 133150 688230 133170 688470
rect 122170 688140 133170 688230
rect 122170 687900 122190 688140
rect 122430 687900 122520 688140
rect 122760 687900 122850 688140
rect 123090 687900 123180 688140
rect 123420 687900 123530 688140
rect 123770 687900 123860 688140
rect 124100 687900 124190 688140
rect 124430 687900 124520 688140
rect 124760 687900 124870 688140
rect 125110 687900 125200 688140
rect 125440 687900 125530 688140
rect 125770 687900 125860 688140
rect 126100 687900 126210 688140
rect 126450 687900 126540 688140
rect 126780 687900 126870 688140
rect 127110 687900 127200 688140
rect 127440 687900 127550 688140
rect 127790 687900 127880 688140
rect 128120 687900 128210 688140
rect 128450 687900 128540 688140
rect 128780 687900 128890 688140
rect 129130 687900 129220 688140
rect 129460 687900 129550 688140
rect 129790 687900 129880 688140
rect 130120 687900 130230 688140
rect 130470 687900 130560 688140
rect 130800 687900 130890 688140
rect 131130 687900 131220 688140
rect 131460 687900 131570 688140
rect 131810 687900 131900 688140
rect 132140 687900 132230 688140
rect 132470 687900 132560 688140
rect 132800 687900 132910 688140
rect 133150 687900 133170 688140
rect 122170 687790 133170 687900
rect 122170 687550 122190 687790
rect 122430 687550 122520 687790
rect 122760 687550 122850 687790
rect 123090 687550 123180 687790
rect 123420 687550 123530 687790
rect 123770 687550 123860 687790
rect 124100 687550 124190 687790
rect 124430 687550 124520 687790
rect 124760 687550 124870 687790
rect 125110 687550 125200 687790
rect 125440 687550 125530 687790
rect 125770 687550 125860 687790
rect 126100 687550 126210 687790
rect 126450 687550 126540 687790
rect 126780 687550 126870 687790
rect 127110 687550 127200 687790
rect 127440 687550 127550 687790
rect 127790 687550 127880 687790
rect 128120 687550 128210 687790
rect 128450 687550 128540 687790
rect 128780 687550 128890 687790
rect 129130 687550 129220 687790
rect 129460 687550 129550 687790
rect 129790 687550 129880 687790
rect 130120 687550 130230 687790
rect 130470 687550 130560 687790
rect 130800 687550 130890 687790
rect 131130 687550 131220 687790
rect 131460 687550 131570 687790
rect 131810 687550 131900 687790
rect 132140 687550 132230 687790
rect 132470 687550 132560 687790
rect 132800 687550 132910 687790
rect 133150 687550 133170 687790
rect 122170 687460 133170 687550
rect 122170 687220 122190 687460
rect 122430 687220 122520 687460
rect 122760 687220 122850 687460
rect 123090 687220 123180 687460
rect 123420 687220 123530 687460
rect 123770 687220 123860 687460
rect 124100 687220 124190 687460
rect 124430 687220 124520 687460
rect 124760 687220 124870 687460
rect 125110 687220 125200 687460
rect 125440 687220 125530 687460
rect 125770 687220 125860 687460
rect 126100 687220 126210 687460
rect 126450 687220 126540 687460
rect 126780 687220 126870 687460
rect 127110 687220 127200 687460
rect 127440 687220 127550 687460
rect 127790 687220 127880 687460
rect 128120 687220 128210 687460
rect 128450 687220 128540 687460
rect 128780 687220 128890 687460
rect 129130 687220 129220 687460
rect 129460 687220 129550 687460
rect 129790 687220 129880 687460
rect 130120 687220 130230 687460
rect 130470 687220 130560 687460
rect 130800 687220 130890 687460
rect 131130 687220 131220 687460
rect 131460 687220 131570 687460
rect 131810 687220 131900 687460
rect 132140 687220 132230 687460
rect 132470 687220 132560 687460
rect 132800 687220 132910 687460
rect 133150 687220 133170 687460
rect 122170 687130 133170 687220
rect 122170 686890 122190 687130
rect 122430 686890 122520 687130
rect 122760 686890 122850 687130
rect 123090 686890 123180 687130
rect 123420 686890 123530 687130
rect 123770 686890 123860 687130
rect 124100 686890 124190 687130
rect 124430 686890 124520 687130
rect 124760 686890 124870 687130
rect 125110 686890 125200 687130
rect 125440 686890 125530 687130
rect 125770 686890 125860 687130
rect 126100 686890 126210 687130
rect 126450 686890 126540 687130
rect 126780 686890 126870 687130
rect 127110 686890 127200 687130
rect 127440 686890 127550 687130
rect 127790 686890 127880 687130
rect 128120 686890 128210 687130
rect 128450 686890 128540 687130
rect 128780 686890 128890 687130
rect 129130 686890 129220 687130
rect 129460 686890 129550 687130
rect 129790 686890 129880 687130
rect 130120 686890 130230 687130
rect 130470 686890 130560 687130
rect 130800 686890 130890 687130
rect 131130 686890 131220 687130
rect 131460 686890 131570 687130
rect 131810 686890 131900 687130
rect 132140 686890 132230 687130
rect 132470 686890 132560 687130
rect 132800 686890 132910 687130
rect 133150 686890 133170 687130
rect 122170 686800 133170 686890
rect 122170 686560 122190 686800
rect 122430 686560 122520 686800
rect 122760 686560 122850 686800
rect 123090 686560 123180 686800
rect 123420 686560 123530 686800
rect 123770 686560 123860 686800
rect 124100 686560 124190 686800
rect 124430 686560 124520 686800
rect 124760 686560 124870 686800
rect 125110 686560 125200 686800
rect 125440 686560 125530 686800
rect 125770 686560 125860 686800
rect 126100 686560 126210 686800
rect 126450 686560 126540 686800
rect 126780 686560 126870 686800
rect 127110 686560 127200 686800
rect 127440 686560 127550 686800
rect 127790 686560 127880 686800
rect 128120 686560 128210 686800
rect 128450 686560 128540 686800
rect 128780 686560 128890 686800
rect 129130 686560 129220 686800
rect 129460 686560 129550 686800
rect 129790 686560 129880 686800
rect 130120 686560 130230 686800
rect 130470 686560 130560 686800
rect 130800 686560 130890 686800
rect 131130 686560 131220 686800
rect 131460 686560 131570 686800
rect 131810 686560 131900 686800
rect 132140 686560 132230 686800
rect 132470 686560 132560 686800
rect 132800 686560 132910 686800
rect 133150 686560 133170 686800
rect 122170 686450 133170 686560
rect 122170 686210 122190 686450
rect 122430 686210 122520 686450
rect 122760 686210 122850 686450
rect 123090 686210 123180 686450
rect 123420 686210 123530 686450
rect 123770 686210 123860 686450
rect 124100 686210 124190 686450
rect 124430 686210 124520 686450
rect 124760 686210 124870 686450
rect 125110 686210 125200 686450
rect 125440 686210 125530 686450
rect 125770 686210 125860 686450
rect 126100 686210 126210 686450
rect 126450 686210 126540 686450
rect 126780 686210 126870 686450
rect 127110 686210 127200 686450
rect 127440 686210 127550 686450
rect 127790 686210 127880 686450
rect 128120 686210 128210 686450
rect 128450 686210 128540 686450
rect 128780 686210 128890 686450
rect 129130 686210 129220 686450
rect 129460 686210 129550 686450
rect 129790 686210 129880 686450
rect 130120 686210 130230 686450
rect 130470 686210 130560 686450
rect 130800 686210 130890 686450
rect 131130 686210 131220 686450
rect 131460 686210 131570 686450
rect 131810 686210 131900 686450
rect 132140 686210 132230 686450
rect 132470 686210 132560 686450
rect 132800 686210 132910 686450
rect 133150 686210 133170 686450
rect 122170 686120 133170 686210
rect 122170 685880 122190 686120
rect 122430 685880 122520 686120
rect 122760 685880 122850 686120
rect 123090 685880 123180 686120
rect 123420 685880 123530 686120
rect 123770 685880 123860 686120
rect 124100 685880 124190 686120
rect 124430 685880 124520 686120
rect 124760 685880 124870 686120
rect 125110 685880 125200 686120
rect 125440 685880 125530 686120
rect 125770 685880 125860 686120
rect 126100 685880 126210 686120
rect 126450 685880 126540 686120
rect 126780 685880 126870 686120
rect 127110 685880 127200 686120
rect 127440 685880 127550 686120
rect 127790 685880 127880 686120
rect 128120 685880 128210 686120
rect 128450 685880 128540 686120
rect 128780 685880 128890 686120
rect 129130 685880 129220 686120
rect 129460 685880 129550 686120
rect 129790 685880 129880 686120
rect 130120 685880 130230 686120
rect 130470 685880 130560 686120
rect 130800 685880 130890 686120
rect 131130 685880 131220 686120
rect 131460 685880 131570 686120
rect 131810 685880 131900 686120
rect 132140 685880 132230 686120
rect 132470 685880 132560 686120
rect 132800 685880 132910 686120
rect 133150 685880 133170 686120
rect 122170 685790 133170 685880
rect 122170 685550 122190 685790
rect 122430 685550 122520 685790
rect 122760 685550 122850 685790
rect 123090 685550 123180 685790
rect 123420 685550 123530 685790
rect 123770 685550 123860 685790
rect 124100 685550 124190 685790
rect 124430 685550 124520 685790
rect 124760 685550 124870 685790
rect 125110 685550 125200 685790
rect 125440 685550 125530 685790
rect 125770 685550 125860 685790
rect 126100 685550 126210 685790
rect 126450 685550 126540 685790
rect 126780 685550 126870 685790
rect 127110 685550 127200 685790
rect 127440 685550 127550 685790
rect 127790 685550 127880 685790
rect 128120 685550 128210 685790
rect 128450 685550 128540 685790
rect 128780 685550 128890 685790
rect 129130 685550 129220 685790
rect 129460 685550 129550 685790
rect 129790 685550 129880 685790
rect 130120 685550 130230 685790
rect 130470 685550 130560 685790
rect 130800 685550 130890 685790
rect 131130 685550 131220 685790
rect 131460 685550 131570 685790
rect 131810 685550 131900 685790
rect 132140 685550 132230 685790
rect 132470 685550 132560 685790
rect 132800 685550 132910 685790
rect 133150 685550 133170 685790
rect 122170 685460 133170 685550
rect 122170 685220 122190 685460
rect 122430 685220 122520 685460
rect 122760 685220 122850 685460
rect 123090 685220 123180 685460
rect 123420 685220 123530 685460
rect 123770 685220 123860 685460
rect 124100 685220 124190 685460
rect 124430 685220 124520 685460
rect 124760 685220 124870 685460
rect 125110 685220 125200 685460
rect 125440 685220 125530 685460
rect 125770 685220 125860 685460
rect 126100 685220 126210 685460
rect 126450 685220 126540 685460
rect 126780 685220 126870 685460
rect 127110 685220 127200 685460
rect 127440 685220 127550 685460
rect 127790 685220 127880 685460
rect 128120 685220 128210 685460
rect 128450 685220 128540 685460
rect 128780 685220 128890 685460
rect 129130 685220 129220 685460
rect 129460 685220 129550 685460
rect 129790 685220 129880 685460
rect 130120 685220 130230 685460
rect 130470 685220 130560 685460
rect 130800 685220 130890 685460
rect 131130 685220 131220 685460
rect 131460 685220 131570 685460
rect 131810 685220 131900 685460
rect 132140 685220 132230 685460
rect 132470 685220 132560 685460
rect 132800 685220 132910 685460
rect 133150 685220 133170 685460
rect 122170 685110 133170 685220
rect 122170 684870 122190 685110
rect 122430 684870 122520 685110
rect 122760 684870 122850 685110
rect 123090 684870 123180 685110
rect 123420 684870 123530 685110
rect 123770 684870 123860 685110
rect 124100 684870 124190 685110
rect 124430 684870 124520 685110
rect 124760 684870 124870 685110
rect 125110 684870 125200 685110
rect 125440 684870 125530 685110
rect 125770 684870 125860 685110
rect 126100 684870 126210 685110
rect 126450 684870 126540 685110
rect 126780 684870 126870 685110
rect 127110 684870 127200 685110
rect 127440 684870 127550 685110
rect 127790 684870 127880 685110
rect 128120 684870 128210 685110
rect 128450 684870 128540 685110
rect 128780 684870 128890 685110
rect 129130 684870 129220 685110
rect 129460 684870 129550 685110
rect 129790 684870 129880 685110
rect 130120 684870 130230 685110
rect 130470 684870 130560 685110
rect 130800 684870 130890 685110
rect 131130 684870 131220 685110
rect 131460 684870 131570 685110
rect 131810 684870 131900 685110
rect 132140 684870 132230 685110
rect 132470 684870 132560 685110
rect 132800 684870 132910 685110
rect 133150 684870 133170 685110
rect 122170 684780 133170 684870
rect 122170 684540 122190 684780
rect 122430 684540 122520 684780
rect 122760 684540 122850 684780
rect 123090 684540 123180 684780
rect 123420 684540 123530 684780
rect 123770 684540 123860 684780
rect 124100 684540 124190 684780
rect 124430 684540 124520 684780
rect 124760 684540 124870 684780
rect 125110 684540 125200 684780
rect 125440 684540 125530 684780
rect 125770 684540 125860 684780
rect 126100 684540 126210 684780
rect 126450 684540 126540 684780
rect 126780 684540 126870 684780
rect 127110 684540 127200 684780
rect 127440 684540 127550 684780
rect 127790 684540 127880 684780
rect 128120 684540 128210 684780
rect 128450 684540 128540 684780
rect 128780 684540 128890 684780
rect 129130 684540 129220 684780
rect 129460 684540 129550 684780
rect 129790 684540 129880 684780
rect 130120 684540 130230 684780
rect 130470 684540 130560 684780
rect 130800 684540 130890 684780
rect 131130 684540 131220 684780
rect 131460 684540 131570 684780
rect 131810 684540 131900 684780
rect 132140 684540 132230 684780
rect 132470 684540 132560 684780
rect 132800 684540 132910 684780
rect 133150 684540 133170 684780
rect 122170 684450 133170 684540
rect 122170 684210 122190 684450
rect 122430 684210 122520 684450
rect 122760 684210 122850 684450
rect 123090 684210 123180 684450
rect 123420 684210 123530 684450
rect 123770 684210 123860 684450
rect 124100 684210 124190 684450
rect 124430 684210 124520 684450
rect 124760 684210 124870 684450
rect 125110 684210 125200 684450
rect 125440 684210 125530 684450
rect 125770 684210 125860 684450
rect 126100 684210 126210 684450
rect 126450 684210 126540 684450
rect 126780 684210 126870 684450
rect 127110 684210 127200 684450
rect 127440 684210 127550 684450
rect 127790 684210 127880 684450
rect 128120 684210 128210 684450
rect 128450 684210 128540 684450
rect 128780 684210 128890 684450
rect 129130 684210 129220 684450
rect 129460 684210 129550 684450
rect 129790 684210 129880 684450
rect 130120 684210 130230 684450
rect 130470 684210 130560 684450
rect 130800 684210 130890 684450
rect 131130 684210 131220 684450
rect 131460 684210 131570 684450
rect 131810 684210 131900 684450
rect 132140 684210 132230 684450
rect 132470 684210 132560 684450
rect 132800 684210 132910 684450
rect 133150 684210 133170 684450
rect 122170 684120 133170 684210
rect 122170 683880 122190 684120
rect 122430 683880 122520 684120
rect 122760 683880 122850 684120
rect 123090 683880 123180 684120
rect 123420 683880 123530 684120
rect 123770 683880 123860 684120
rect 124100 683880 124190 684120
rect 124430 683880 124520 684120
rect 124760 683880 124870 684120
rect 125110 683880 125200 684120
rect 125440 683880 125530 684120
rect 125770 683880 125860 684120
rect 126100 683880 126210 684120
rect 126450 683880 126540 684120
rect 126780 683880 126870 684120
rect 127110 683880 127200 684120
rect 127440 683880 127550 684120
rect 127790 683880 127880 684120
rect 128120 683880 128210 684120
rect 128450 683880 128540 684120
rect 128780 683880 128890 684120
rect 129130 683880 129220 684120
rect 129460 683880 129550 684120
rect 129790 683880 129880 684120
rect 130120 683880 130230 684120
rect 130470 683880 130560 684120
rect 130800 683880 130890 684120
rect 131130 683880 131220 684120
rect 131460 683880 131570 684120
rect 131810 683880 131900 684120
rect 132140 683880 132230 684120
rect 132470 683880 132560 684120
rect 132800 683880 132910 684120
rect 133150 683880 133170 684120
rect 122170 683860 133170 683880
rect 133550 694840 144550 694860
rect 133550 694600 133570 694840
rect 133810 694600 133900 694840
rect 134140 694600 134230 694840
rect 134470 694600 134560 694840
rect 134800 694600 134910 694840
rect 135150 694600 135240 694840
rect 135480 694600 135570 694840
rect 135810 694600 135900 694840
rect 136140 694600 136250 694840
rect 136490 694600 136580 694840
rect 136820 694600 136910 694840
rect 137150 694600 137240 694840
rect 137480 694600 137590 694840
rect 137830 694600 137920 694840
rect 138160 694600 138250 694840
rect 138490 694600 138580 694840
rect 138820 694600 138930 694840
rect 139170 694600 139260 694840
rect 139500 694600 139590 694840
rect 139830 694600 139920 694840
rect 140160 694600 140270 694840
rect 140510 694600 140600 694840
rect 140840 694600 140930 694840
rect 141170 694600 141260 694840
rect 141500 694600 141610 694840
rect 141850 694600 141940 694840
rect 142180 694600 142270 694840
rect 142510 694600 142600 694840
rect 142840 694600 142950 694840
rect 143190 694600 143280 694840
rect 143520 694600 143610 694840
rect 143850 694600 143940 694840
rect 144180 694600 144290 694840
rect 144530 694600 144550 694840
rect 133550 694490 144550 694600
rect 133550 694250 133570 694490
rect 133810 694250 133900 694490
rect 134140 694250 134230 694490
rect 134470 694250 134560 694490
rect 134800 694250 134910 694490
rect 135150 694250 135240 694490
rect 135480 694250 135570 694490
rect 135810 694250 135900 694490
rect 136140 694250 136250 694490
rect 136490 694250 136580 694490
rect 136820 694250 136910 694490
rect 137150 694250 137240 694490
rect 137480 694250 137590 694490
rect 137830 694250 137920 694490
rect 138160 694250 138250 694490
rect 138490 694250 138580 694490
rect 138820 694250 138930 694490
rect 139170 694250 139260 694490
rect 139500 694250 139590 694490
rect 139830 694250 139920 694490
rect 140160 694250 140270 694490
rect 140510 694250 140600 694490
rect 140840 694250 140930 694490
rect 141170 694250 141260 694490
rect 141500 694250 141610 694490
rect 141850 694250 141940 694490
rect 142180 694250 142270 694490
rect 142510 694250 142600 694490
rect 142840 694250 142950 694490
rect 143190 694250 143280 694490
rect 143520 694250 143610 694490
rect 143850 694250 143940 694490
rect 144180 694250 144290 694490
rect 144530 694250 144550 694490
rect 133550 694160 144550 694250
rect 133550 693920 133570 694160
rect 133810 693920 133900 694160
rect 134140 693920 134230 694160
rect 134470 693920 134560 694160
rect 134800 693920 134910 694160
rect 135150 693920 135240 694160
rect 135480 693920 135570 694160
rect 135810 693920 135900 694160
rect 136140 693920 136250 694160
rect 136490 693920 136580 694160
rect 136820 693920 136910 694160
rect 137150 693920 137240 694160
rect 137480 693920 137590 694160
rect 137830 693920 137920 694160
rect 138160 693920 138250 694160
rect 138490 693920 138580 694160
rect 138820 693920 138930 694160
rect 139170 693920 139260 694160
rect 139500 693920 139590 694160
rect 139830 693920 139920 694160
rect 140160 693920 140270 694160
rect 140510 693920 140600 694160
rect 140840 693920 140930 694160
rect 141170 693920 141260 694160
rect 141500 693920 141610 694160
rect 141850 693920 141940 694160
rect 142180 693920 142270 694160
rect 142510 693920 142600 694160
rect 142840 693920 142950 694160
rect 143190 693920 143280 694160
rect 143520 693920 143610 694160
rect 143850 693920 143940 694160
rect 144180 693920 144290 694160
rect 144530 693920 144550 694160
rect 133550 693830 144550 693920
rect 133550 693590 133570 693830
rect 133810 693590 133900 693830
rect 134140 693590 134230 693830
rect 134470 693590 134560 693830
rect 134800 693590 134910 693830
rect 135150 693590 135240 693830
rect 135480 693590 135570 693830
rect 135810 693590 135900 693830
rect 136140 693590 136250 693830
rect 136490 693590 136580 693830
rect 136820 693590 136910 693830
rect 137150 693590 137240 693830
rect 137480 693590 137590 693830
rect 137830 693590 137920 693830
rect 138160 693590 138250 693830
rect 138490 693590 138580 693830
rect 138820 693590 138930 693830
rect 139170 693590 139260 693830
rect 139500 693590 139590 693830
rect 139830 693590 139920 693830
rect 140160 693590 140270 693830
rect 140510 693590 140600 693830
rect 140840 693590 140930 693830
rect 141170 693590 141260 693830
rect 141500 693590 141610 693830
rect 141850 693590 141940 693830
rect 142180 693590 142270 693830
rect 142510 693590 142600 693830
rect 142840 693590 142950 693830
rect 143190 693590 143280 693830
rect 143520 693590 143610 693830
rect 143850 693590 143940 693830
rect 144180 693590 144290 693830
rect 144530 693590 144550 693830
rect 133550 693500 144550 693590
rect 133550 693260 133570 693500
rect 133810 693260 133900 693500
rect 134140 693260 134230 693500
rect 134470 693260 134560 693500
rect 134800 693260 134910 693500
rect 135150 693260 135240 693500
rect 135480 693260 135570 693500
rect 135810 693260 135900 693500
rect 136140 693260 136250 693500
rect 136490 693260 136580 693500
rect 136820 693260 136910 693500
rect 137150 693260 137240 693500
rect 137480 693260 137590 693500
rect 137830 693260 137920 693500
rect 138160 693260 138250 693500
rect 138490 693260 138580 693500
rect 138820 693260 138930 693500
rect 139170 693260 139260 693500
rect 139500 693260 139590 693500
rect 139830 693260 139920 693500
rect 140160 693260 140270 693500
rect 140510 693260 140600 693500
rect 140840 693260 140930 693500
rect 141170 693260 141260 693500
rect 141500 693260 141610 693500
rect 141850 693260 141940 693500
rect 142180 693260 142270 693500
rect 142510 693260 142600 693500
rect 142840 693260 142950 693500
rect 143190 693260 143280 693500
rect 143520 693260 143610 693500
rect 143850 693260 143940 693500
rect 144180 693260 144290 693500
rect 144530 693260 144550 693500
rect 133550 693150 144550 693260
rect 133550 692910 133570 693150
rect 133810 692910 133900 693150
rect 134140 692910 134230 693150
rect 134470 692910 134560 693150
rect 134800 692910 134910 693150
rect 135150 692910 135240 693150
rect 135480 692910 135570 693150
rect 135810 692910 135900 693150
rect 136140 692910 136250 693150
rect 136490 692910 136580 693150
rect 136820 692910 136910 693150
rect 137150 692910 137240 693150
rect 137480 692910 137590 693150
rect 137830 692910 137920 693150
rect 138160 692910 138250 693150
rect 138490 692910 138580 693150
rect 138820 692910 138930 693150
rect 139170 692910 139260 693150
rect 139500 692910 139590 693150
rect 139830 692910 139920 693150
rect 140160 692910 140270 693150
rect 140510 692910 140600 693150
rect 140840 692910 140930 693150
rect 141170 692910 141260 693150
rect 141500 692910 141610 693150
rect 141850 692910 141940 693150
rect 142180 692910 142270 693150
rect 142510 692910 142600 693150
rect 142840 692910 142950 693150
rect 143190 692910 143280 693150
rect 143520 692910 143610 693150
rect 143850 692910 143940 693150
rect 144180 692910 144290 693150
rect 144530 692910 144550 693150
rect 133550 692820 144550 692910
rect 133550 692580 133570 692820
rect 133810 692580 133900 692820
rect 134140 692580 134230 692820
rect 134470 692580 134560 692820
rect 134800 692580 134910 692820
rect 135150 692580 135240 692820
rect 135480 692580 135570 692820
rect 135810 692580 135900 692820
rect 136140 692580 136250 692820
rect 136490 692580 136580 692820
rect 136820 692580 136910 692820
rect 137150 692580 137240 692820
rect 137480 692580 137590 692820
rect 137830 692580 137920 692820
rect 138160 692580 138250 692820
rect 138490 692580 138580 692820
rect 138820 692580 138930 692820
rect 139170 692580 139260 692820
rect 139500 692580 139590 692820
rect 139830 692580 139920 692820
rect 140160 692580 140270 692820
rect 140510 692580 140600 692820
rect 140840 692580 140930 692820
rect 141170 692580 141260 692820
rect 141500 692580 141610 692820
rect 141850 692580 141940 692820
rect 142180 692580 142270 692820
rect 142510 692580 142600 692820
rect 142840 692580 142950 692820
rect 143190 692580 143280 692820
rect 143520 692580 143610 692820
rect 143850 692580 143940 692820
rect 144180 692580 144290 692820
rect 144530 692580 144550 692820
rect 133550 692490 144550 692580
rect 133550 692250 133570 692490
rect 133810 692250 133900 692490
rect 134140 692250 134230 692490
rect 134470 692250 134560 692490
rect 134800 692250 134910 692490
rect 135150 692250 135240 692490
rect 135480 692250 135570 692490
rect 135810 692250 135900 692490
rect 136140 692250 136250 692490
rect 136490 692250 136580 692490
rect 136820 692250 136910 692490
rect 137150 692250 137240 692490
rect 137480 692250 137590 692490
rect 137830 692250 137920 692490
rect 138160 692250 138250 692490
rect 138490 692250 138580 692490
rect 138820 692250 138930 692490
rect 139170 692250 139260 692490
rect 139500 692250 139590 692490
rect 139830 692250 139920 692490
rect 140160 692250 140270 692490
rect 140510 692250 140600 692490
rect 140840 692250 140930 692490
rect 141170 692250 141260 692490
rect 141500 692250 141610 692490
rect 141850 692250 141940 692490
rect 142180 692250 142270 692490
rect 142510 692250 142600 692490
rect 142840 692250 142950 692490
rect 143190 692250 143280 692490
rect 143520 692250 143610 692490
rect 143850 692250 143940 692490
rect 144180 692250 144290 692490
rect 144530 692250 144550 692490
rect 133550 692160 144550 692250
rect 133550 691920 133570 692160
rect 133810 691920 133900 692160
rect 134140 691920 134230 692160
rect 134470 691920 134560 692160
rect 134800 691920 134910 692160
rect 135150 691920 135240 692160
rect 135480 691920 135570 692160
rect 135810 691920 135900 692160
rect 136140 691920 136250 692160
rect 136490 691920 136580 692160
rect 136820 691920 136910 692160
rect 137150 691920 137240 692160
rect 137480 691920 137590 692160
rect 137830 691920 137920 692160
rect 138160 691920 138250 692160
rect 138490 691920 138580 692160
rect 138820 691920 138930 692160
rect 139170 691920 139260 692160
rect 139500 691920 139590 692160
rect 139830 691920 139920 692160
rect 140160 691920 140270 692160
rect 140510 691920 140600 692160
rect 140840 691920 140930 692160
rect 141170 691920 141260 692160
rect 141500 691920 141610 692160
rect 141850 691920 141940 692160
rect 142180 691920 142270 692160
rect 142510 691920 142600 692160
rect 142840 691920 142950 692160
rect 143190 691920 143280 692160
rect 143520 691920 143610 692160
rect 143850 691920 143940 692160
rect 144180 691920 144290 692160
rect 144530 691920 144550 692160
rect 133550 691810 144550 691920
rect 133550 691570 133570 691810
rect 133810 691570 133900 691810
rect 134140 691570 134230 691810
rect 134470 691570 134560 691810
rect 134800 691570 134910 691810
rect 135150 691570 135240 691810
rect 135480 691570 135570 691810
rect 135810 691570 135900 691810
rect 136140 691570 136250 691810
rect 136490 691570 136580 691810
rect 136820 691570 136910 691810
rect 137150 691570 137240 691810
rect 137480 691570 137590 691810
rect 137830 691570 137920 691810
rect 138160 691570 138250 691810
rect 138490 691570 138580 691810
rect 138820 691570 138930 691810
rect 139170 691570 139260 691810
rect 139500 691570 139590 691810
rect 139830 691570 139920 691810
rect 140160 691570 140270 691810
rect 140510 691570 140600 691810
rect 140840 691570 140930 691810
rect 141170 691570 141260 691810
rect 141500 691570 141610 691810
rect 141850 691570 141940 691810
rect 142180 691570 142270 691810
rect 142510 691570 142600 691810
rect 142840 691570 142950 691810
rect 143190 691570 143280 691810
rect 143520 691570 143610 691810
rect 143850 691570 143940 691810
rect 144180 691570 144290 691810
rect 144530 691570 144550 691810
rect 133550 691480 144550 691570
rect 133550 691240 133570 691480
rect 133810 691240 133900 691480
rect 134140 691240 134230 691480
rect 134470 691240 134560 691480
rect 134800 691240 134910 691480
rect 135150 691240 135240 691480
rect 135480 691240 135570 691480
rect 135810 691240 135900 691480
rect 136140 691240 136250 691480
rect 136490 691240 136580 691480
rect 136820 691240 136910 691480
rect 137150 691240 137240 691480
rect 137480 691240 137590 691480
rect 137830 691240 137920 691480
rect 138160 691240 138250 691480
rect 138490 691240 138580 691480
rect 138820 691240 138930 691480
rect 139170 691240 139260 691480
rect 139500 691240 139590 691480
rect 139830 691240 139920 691480
rect 140160 691240 140270 691480
rect 140510 691240 140600 691480
rect 140840 691240 140930 691480
rect 141170 691240 141260 691480
rect 141500 691240 141610 691480
rect 141850 691240 141940 691480
rect 142180 691240 142270 691480
rect 142510 691240 142600 691480
rect 142840 691240 142950 691480
rect 143190 691240 143280 691480
rect 143520 691240 143610 691480
rect 143850 691240 143940 691480
rect 144180 691240 144290 691480
rect 144530 691240 144550 691480
rect 133550 691150 144550 691240
rect 133550 690910 133570 691150
rect 133810 690910 133900 691150
rect 134140 690910 134230 691150
rect 134470 690910 134560 691150
rect 134800 690910 134910 691150
rect 135150 690910 135240 691150
rect 135480 690910 135570 691150
rect 135810 690910 135900 691150
rect 136140 690910 136250 691150
rect 136490 690910 136580 691150
rect 136820 690910 136910 691150
rect 137150 690910 137240 691150
rect 137480 690910 137590 691150
rect 137830 690910 137920 691150
rect 138160 690910 138250 691150
rect 138490 690910 138580 691150
rect 138820 690910 138930 691150
rect 139170 690910 139260 691150
rect 139500 690910 139590 691150
rect 139830 690910 139920 691150
rect 140160 690910 140270 691150
rect 140510 690910 140600 691150
rect 140840 690910 140930 691150
rect 141170 690910 141260 691150
rect 141500 690910 141610 691150
rect 141850 690910 141940 691150
rect 142180 690910 142270 691150
rect 142510 690910 142600 691150
rect 142840 690910 142950 691150
rect 143190 690910 143280 691150
rect 143520 690910 143610 691150
rect 143850 690910 143940 691150
rect 144180 690910 144290 691150
rect 144530 690910 144550 691150
rect 133550 690820 144550 690910
rect 133550 690580 133570 690820
rect 133810 690580 133900 690820
rect 134140 690580 134230 690820
rect 134470 690580 134560 690820
rect 134800 690580 134910 690820
rect 135150 690580 135240 690820
rect 135480 690580 135570 690820
rect 135810 690580 135900 690820
rect 136140 690580 136250 690820
rect 136490 690580 136580 690820
rect 136820 690580 136910 690820
rect 137150 690580 137240 690820
rect 137480 690580 137590 690820
rect 137830 690580 137920 690820
rect 138160 690580 138250 690820
rect 138490 690580 138580 690820
rect 138820 690580 138930 690820
rect 139170 690580 139260 690820
rect 139500 690580 139590 690820
rect 139830 690580 139920 690820
rect 140160 690580 140270 690820
rect 140510 690580 140600 690820
rect 140840 690580 140930 690820
rect 141170 690580 141260 690820
rect 141500 690580 141610 690820
rect 141850 690580 141940 690820
rect 142180 690580 142270 690820
rect 142510 690580 142600 690820
rect 142840 690580 142950 690820
rect 143190 690580 143280 690820
rect 143520 690580 143610 690820
rect 143850 690580 143940 690820
rect 144180 690580 144290 690820
rect 144530 690580 144550 690820
rect 133550 690470 144550 690580
rect 133550 690230 133570 690470
rect 133810 690230 133900 690470
rect 134140 690230 134230 690470
rect 134470 690230 134560 690470
rect 134800 690230 134910 690470
rect 135150 690230 135240 690470
rect 135480 690230 135570 690470
rect 135810 690230 135900 690470
rect 136140 690230 136250 690470
rect 136490 690230 136580 690470
rect 136820 690230 136910 690470
rect 137150 690230 137240 690470
rect 137480 690230 137590 690470
rect 137830 690230 137920 690470
rect 138160 690230 138250 690470
rect 138490 690230 138580 690470
rect 138820 690230 138930 690470
rect 139170 690230 139260 690470
rect 139500 690230 139590 690470
rect 139830 690230 139920 690470
rect 140160 690230 140270 690470
rect 140510 690230 140600 690470
rect 140840 690230 140930 690470
rect 141170 690230 141260 690470
rect 141500 690230 141610 690470
rect 141850 690230 141940 690470
rect 142180 690230 142270 690470
rect 142510 690230 142600 690470
rect 142840 690230 142950 690470
rect 143190 690230 143280 690470
rect 143520 690230 143610 690470
rect 143850 690230 143940 690470
rect 144180 690230 144290 690470
rect 144530 690230 144550 690470
rect 133550 690140 144550 690230
rect 133550 689900 133570 690140
rect 133810 689900 133900 690140
rect 134140 689900 134230 690140
rect 134470 689900 134560 690140
rect 134800 689900 134910 690140
rect 135150 689900 135240 690140
rect 135480 689900 135570 690140
rect 135810 689900 135900 690140
rect 136140 689900 136250 690140
rect 136490 689900 136580 690140
rect 136820 689900 136910 690140
rect 137150 689900 137240 690140
rect 137480 689900 137590 690140
rect 137830 689900 137920 690140
rect 138160 689900 138250 690140
rect 138490 689900 138580 690140
rect 138820 689900 138930 690140
rect 139170 689900 139260 690140
rect 139500 689900 139590 690140
rect 139830 689900 139920 690140
rect 140160 689900 140270 690140
rect 140510 689900 140600 690140
rect 140840 689900 140930 690140
rect 141170 689900 141260 690140
rect 141500 689900 141610 690140
rect 141850 689900 141940 690140
rect 142180 689900 142270 690140
rect 142510 689900 142600 690140
rect 142840 689900 142950 690140
rect 143190 689900 143280 690140
rect 143520 689900 143610 690140
rect 143850 689900 143940 690140
rect 144180 689900 144290 690140
rect 144530 689900 144550 690140
rect 133550 689810 144550 689900
rect 133550 689570 133570 689810
rect 133810 689570 133900 689810
rect 134140 689570 134230 689810
rect 134470 689570 134560 689810
rect 134800 689570 134910 689810
rect 135150 689570 135240 689810
rect 135480 689570 135570 689810
rect 135810 689570 135900 689810
rect 136140 689570 136250 689810
rect 136490 689570 136580 689810
rect 136820 689570 136910 689810
rect 137150 689570 137240 689810
rect 137480 689570 137590 689810
rect 137830 689570 137920 689810
rect 138160 689570 138250 689810
rect 138490 689570 138580 689810
rect 138820 689570 138930 689810
rect 139170 689570 139260 689810
rect 139500 689570 139590 689810
rect 139830 689570 139920 689810
rect 140160 689570 140270 689810
rect 140510 689570 140600 689810
rect 140840 689570 140930 689810
rect 141170 689570 141260 689810
rect 141500 689570 141610 689810
rect 141850 689570 141940 689810
rect 142180 689570 142270 689810
rect 142510 689570 142600 689810
rect 142840 689570 142950 689810
rect 143190 689570 143280 689810
rect 143520 689570 143610 689810
rect 143850 689570 143940 689810
rect 144180 689570 144290 689810
rect 144530 689570 144550 689810
rect 133550 689480 144550 689570
rect 133550 689240 133570 689480
rect 133810 689240 133900 689480
rect 134140 689240 134230 689480
rect 134470 689240 134560 689480
rect 134800 689240 134910 689480
rect 135150 689240 135240 689480
rect 135480 689240 135570 689480
rect 135810 689240 135900 689480
rect 136140 689240 136250 689480
rect 136490 689240 136580 689480
rect 136820 689240 136910 689480
rect 137150 689240 137240 689480
rect 137480 689240 137590 689480
rect 137830 689240 137920 689480
rect 138160 689240 138250 689480
rect 138490 689240 138580 689480
rect 138820 689240 138930 689480
rect 139170 689240 139260 689480
rect 139500 689240 139590 689480
rect 139830 689240 139920 689480
rect 140160 689240 140270 689480
rect 140510 689240 140600 689480
rect 140840 689240 140930 689480
rect 141170 689240 141260 689480
rect 141500 689240 141610 689480
rect 141850 689240 141940 689480
rect 142180 689240 142270 689480
rect 142510 689240 142600 689480
rect 142840 689240 142950 689480
rect 143190 689240 143280 689480
rect 143520 689240 143610 689480
rect 143850 689240 143940 689480
rect 144180 689240 144290 689480
rect 144530 689240 144550 689480
rect 133550 689130 144550 689240
rect 133550 688890 133570 689130
rect 133810 688890 133900 689130
rect 134140 688890 134230 689130
rect 134470 688890 134560 689130
rect 134800 688890 134910 689130
rect 135150 688890 135240 689130
rect 135480 688890 135570 689130
rect 135810 688890 135900 689130
rect 136140 688890 136250 689130
rect 136490 688890 136580 689130
rect 136820 688890 136910 689130
rect 137150 688890 137240 689130
rect 137480 688890 137590 689130
rect 137830 688890 137920 689130
rect 138160 688890 138250 689130
rect 138490 688890 138580 689130
rect 138820 688890 138930 689130
rect 139170 688890 139260 689130
rect 139500 688890 139590 689130
rect 139830 688890 139920 689130
rect 140160 688890 140270 689130
rect 140510 688890 140600 689130
rect 140840 688890 140930 689130
rect 141170 688890 141260 689130
rect 141500 688890 141610 689130
rect 141850 688890 141940 689130
rect 142180 688890 142270 689130
rect 142510 688890 142600 689130
rect 142840 688890 142950 689130
rect 143190 688890 143280 689130
rect 143520 688890 143610 689130
rect 143850 688890 143940 689130
rect 144180 688890 144290 689130
rect 144530 688890 144550 689130
rect 133550 688800 144550 688890
rect 133550 688560 133570 688800
rect 133810 688560 133900 688800
rect 134140 688560 134230 688800
rect 134470 688560 134560 688800
rect 134800 688560 134910 688800
rect 135150 688560 135240 688800
rect 135480 688560 135570 688800
rect 135810 688560 135900 688800
rect 136140 688560 136250 688800
rect 136490 688560 136580 688800
rect 136820 688560 136910 688800
rect 137150 688560 137240 688800
rect 137480 688560 137590 688800
rect 137830 688560 137920 688800
rect 138160 688560 138250 688800
rect 138490 688560 138580 688800
rect 138820 688560 138930 688800
rect 139170 688560 139260 688800
rect 139500 688560 139590 688800
rect 139830 688560 139920 688800
rect 140160 688560 140270 688800
rect 140510 688560 140600 688800
rect 140840 688560 140930 688800
rect 141170 688560 141260 688800
rect 141500 688560 141610 688800
rect 141850 688560 141940 688800
rect 142180 688560 142270 688800
rect 142510 688560 142600 688800
rect 142840 688560 142950 688800
rect 143190 688560 143280 688800
rect 143520 688560 143610 688800
rect 143850 688560 143940 688800
rect 144180 688560 144290 688800
rect 144530 688560 144550 688800
rect 133550 688470 144550 688560
rect 133550 688230 133570 688470
rect 133810 688230 133900 688470
rect 134140 688230 134230 688470
rect 134470 688230 134560 688470
rect 134800 688230 134910 688470
rect 135150 688230 135240 688470
rect 135480 688230 135570 688470
rect 135810 688230 135900 688470
rect 136140 688230 136250 688470
rect 136490 688230 136580 688470
rect 136820 688230 136910 688470
rect 137150 688230 137240 688470
rect 137480 688230 137590 688470
rect 137830 688230 137920 688470
rect 138160 688230 138250 688470
rect 138490 688230 138580 688470
rect 138820 688230 138930 688470
rect 139170 688230 139260 688470
rect 139500 688230 139590 688470
rect 139830 688230 139920 688470
rect 140160 688230 140270 688470
rect 140510 688230 140600 688470
rect 140840 688230 140930 688470
rect 141170 688230 141260 688470
rect 141500 688230 141610 688470
rect 141850 688230 141940 688470
rect 142180 688230 142270 688470
rect 142510 688230 142600 688470
rect 142840 688230 142950 688470
rect 143190 688230 143280 688470
rect 143520 688230 143610 688470
rect 143850 688230 143940 688470
rect 144180 688230 144290 688470
rect 144530 688230 144550 688470
rect 133550 688140 144550 688230
rect 133550 687900 133570 688140
rect 133810 687900 133900 688140
rect 134140 687900 134230 688140
rect 134470 687900 134560 688140
rect 134800 687900 134910 688140
rect 135150 687900 135240 688140
rect 135480 687900 135570 688140
rect 135810 687900 135900 688140
rect 136140 687900 136250 688140
rect 136490 687900 136580 688140
rect 136820 687900 136910 688140
rect 137150 687900 137240 688140
rect 137480 687900 137590 688140
rect 137830 687900 137920 688140
rect 138160 687900 138250 688140
rect 138490 687900 138580 688140
rect 138820 687900 138930 688140
rect 139170 687900 139260 688140
rect 139500 687900 139590 688140
rect 139830 687900 139920 688140
rect 140160 687900 140270 688140
rect 140510 687900 140600 688140
rect 140840 687900 140930 688140
rect 141170 687900 141260 688140
rect 141500 687900 141610 688140
rect 141850 687900 141940 688140
rect 142180 687900 142270 688140
rect 142510 687900 142600 688140
rect 142840 687900 142950 688140
rect 143190 687900 143280 688140
rect 143520 687900 143610 688140
rect 143850 687900 143940 688140
rect 144180 687900 144290 688140
rect 144530 687900 144550 688140
rect 133550 687790 144550 687900
rect 133550 687550 133570 687790
rect 133810 687550 133900 687790
rect 134140 687550 134230 687790
rect 134470 687550 134560 687790
rect 134800 687550 134910 687790
rect 135150 687550 135240 687790
rect 135480 687550 135570 687790
rect 135810 687550 135900 687790
rect 136140 687550 136250 687790
rect 136490 687550 136580 687790
rect 136820 687550 136910 687790
rect 137150 687550 137240 687790
rect 137480 687550 137590 687790
rect 137830 687550 137920 687790
rect 138160 687550 138250 687790
rect 138490 687550 138580 687790
rect 138820 687550 138930 687790
rect 139170 687550 139260 687790
rect 139500 687550 139590 687790
rect 139830 687550 139920 687790
rect 140160 687550 140270 687790
rect 140510 687550 140600 687790
rect 140840 687550 140930 687790
rect 141170 687550 141260 687790
rect 141500 687550 141610 687790
rect 141850 687550 141940 687790
rect 142180 687550 142270 687790
rect 142510 687550 142600 687790
rect 142840 687550 142950 687790
rect 143190 687550 143280 687790
rect 143520 687550 143610 687790
rect 143850 687550 143940 687790
rect 144180 687550 144290 687790
rect 144530 687550 144550 687790
rect 133550 687460 144550 687550
rect 133550 687220 133570 687460
rect 133810 687220 133900 687460
rect 134140 687220 134230 687460
rect 134470 687220 134560 687460
rect 134800 687220 134910 687460
rect 135150 687220 135240 687460
rect 135480 687220 135570 687460
rect 135810 687220 135900 687460
rect 136140 687220 136250 687460
rect 136490 687220 136580 687460
rect 136820 687220 136910 687460
rect 137150 687220 137240 687460
rect 137480 687220 137590 687460
rect 137830 687220 137920 687460
rect 138160 687220 138250 687460
rect 138490 687220 138580 687460
rect 138820 687220 138930 687460
rect 139170 687220 139260 687460
rect 139500 687220 139590 687460
rect 139830 687220 139920 687460
rect 140160 687220 140270 687460
rect 140510 687220 140600 687460
rect 140840 687220 140930 687460
rect 141170 687220 141260 687460
rect 141500 687220 141610 687460
rect 141850 687220 141940 687460
rect 142180 687220 142270 687460
rect 142510 687220 142600 687460
rect 142840 687220 142950 687460
rect 143190 687220 143280 687460
rect 143520 687220 143610 687460
rect 143850 687220 143940 687460
rect 144180 687220 144290 687460
rect 144530 687220 144550 687460
rect 133550 687130 144550 687220
rect 133550 686890 133570 687130
rect 133810 686890 133900 687130
rect 134140 686890 134230 687130
rect 134470 686890 134560 687130
rect 134800 686890 134910 687130
rect 135150 686890 135240 687130
rect 135480 686890 135570 687130
rect 135810 686890 135900 687130
rect 136140 686890 136250 687130
rect 136490 686890 136580 687130
rect 136820 686890 136910 687130
rect 137150 686890 137240 687130
rect 137480 686890 137590 687130
rect 137830 686890 137920 687130
rect 138160 686890 138250 687130
rect 138490 686890 138580 687130
rect 138820 686890 138930 687130
rect 139170 686890 139260 687130
rect 139500 686890 139590 687130
rect 139830 686890 139920 687130
rect 140160 686890 140270 687130
rect 140510 686890 140600 687130
rect 140840 686890 140930 687130
rect 141170 686890 141260 687130
rect 141500 686890 141610 687130
rect 141850 686890 141940 687130
rect 142180 686890 142270 687130
rect 142510 686890 142600 687130
rect 142840 686890 142950 687130
rect 143190 686890 143280 687130
rect 143520 686890 143610 687130
rect 143850 686890 143940 687130
rect 144180 686890 144290 687130
rect 144530 686890 144550 687130
rect 133550 686800 144550 686890
rect 133550 686560 133570 686800
rect 133810 686560 133900 686800
rect 134140 686560 134230 686800
rect 134470 686560 134560 686800
rect 134800 686560 134910 686800
rect 135150 686560 135240 686800
rect 135480 686560 135570 686800
rect 135810 686560 135900 686800
rect 136140 686560 136250 686800
rect 136490 686560 136580 686800
rect 136820 686560 136910 686800
rect 137150 686560 137240 686800
rect 137480 686560 137590 686800
rect 137830 686560 137920 686800
rect 138160 686560 138250 686800
rect 138490 686560 138580 686800
rect 138820 686560 138930 686800
rect 139170 686560 139260 686800
rect 139500 686560 139590 686800
rect 139830 686560 139920 686800
rect 140160 686560 140270 686800
rect 140510 686560 140600 686800
rect 140840 686560 140930 686800
rect 141170 686560 141260 686800
rect 141500 686560 141610 686800
rect 141850 686560 141940 686800
rect 142180 686560 142270 686800
rect 142510 686560 142600 686800
rect 142840 686560 142950 686800
rect 143190 686560 143280 686800
rect 143520 686560 143610 686800
rect 143850 686560 143940 686800
rect 144180 686560 144290 686800
rect 144530 686560 144550 686800
rect 133550 686450 144550 686560
rect 133550 686210 133570 686450
rect 133810 686210 133900 686450
rect 134140 686210 134230 686450
rect 134470 686210 134560 686450
rect 134800 686210 134910 686450
rect 135150 686210 135240 686450
rect 135480 686210 135570 686450
rect 135810 686210 135900 686450
rect 136140 686210 136250 686450
rect 136490 686210 136580 686450
rect 136820 686210 136910 686450
rect 137150 686210 137240 686450
rect 137480 686210 137590 686450
rect 137830 686210 137920 686450
rect 138160 686210 138250 686450
rect 138490 686210 138580 686450
rect 138820 686210 138930 686450
rect 139170 686210 139260 686450
rect 139500 686210 139590 686450
rect 139830 686210 139920 686450
rect 140160 686210 140270 686450
rect 140510 686210 140600 686450
rect 140840 686210 140930 686450
rect 141170 686210 141260 686450
rect 141500 686210 141610 686450
rect 141850 686210 141940 686450
rect 142180 686210 142270 686450
rect 142510 686210 142600 686450
rect 142840 686210 142950 686450
rect 143190 686210 143280 686450
rect 143520 686210 143610 686450
rect 143850 686210 143940 686450
rect 144180 686210 144290 686450
rect 144530 686210 144550 686450
rect 133550 686120 144550 686210
rect 133550 685880 133570 686120
rect 133810 685880 133900 686120
rect 134140 685880 134230 686120
rect 134470 685880 134560 686120
rect 134800 685880 134910 686120
rect 135150 685880 135240 686120
rect 135480 685880 135570 686120
rect 135810 685880 135900 686120
rect 136140 685880 136250 686120
rect 136490 685880 136580 686120
rect 136820 685880 136910 686120
rect 137150 685880 137240 686120
rect 137480 685880 137590 686120
rect 137830 685880 137920 686120
rect 138160 685880 138250 686120
rect 138490 685880 138580 686120
rect 138820 685880 138930 686120
rect 139170 685880 139260 686120
rect 139500 685880 139590 686120
rect 139830 685880 139920 686120
rect 140160 685880 140270 686120
rect 140510 685880 140600 686120
rect 140840 685880 140930 686120
rect 141170 685880 141260 686120
rect 141500 685880 141610 686120
rect 141850 685880 141940 686120
rect 142180 685880 142270 686120
rect 142510 685880 142600 686120
rect 142840 685880 142950 686120
rect 143190 685880 143280 686120
rect 143520 685880 143610 686120
rect 143850 685880 143940 686120
rect 144180 685880 144290 686120
rect 144530 685880 144550 686120
rect 133550 685790 144550 685880
rect 133550 685550 133570 685790
rect 133810 685550 133900 685790
rect 134140 685550 134230 685790
rect 134470 685550 134560 685790
rect 134800 685550 134910 685790
rect 135150 685550 135240 685790
rect 135480 685550 135570 685790
rect 135810 685550 135900 685790
rect 136140 685550 136250 685790
rect 136490 685550 136580 685790
rect 136820 685550 136910 685790
rect 137150 685550 137240 685790
rect 137480 685550 137590 685790
rect 137830 685550 137920 685790
rect 138160 685550 138250 685790
rect 138490 685550 138580 685790
rect 138820 685550 138930 685790
rect 139170 685550 139260 685790
rect 139500 685550 139590 685790
rect 139830 685550 139920 685790
rect 140160 685550 140270 685790
rect 140510 685550 140600 685790
rect 140840 685550 140930 685790
rect 141170 685550 141260 685790
rect 141500 685550 141610 685790
rect 141850 685550 141940 685790
rect 142180 685550 142270 685790
rect 142510 685550 142600 685790
rect 142840 685550 142950 685790
rect 143190 685550 143280 685790
rect 143520 685550 143610 685790
rect 143850 685550 143940 685790
rect 144180 685550 144290 685790
rect 144530 685550 144550 685790
rect 133550 685460 144550 685550
rect 133550 685220 133570 685460
rect 133810 685220 133900 685460
rect 134140 685220 134230 685460
rect 134470 685220 134560 685460
rect 134800 685220 134910 685460
rect 135150 685220 135240 685460
rect 135480 685220 135570 685460
rect 135810 685220 135900 685460
rect 136140 685220 136250 685460
rect 136490 685220 136580 685460
rect 136820 685220 136910 685460
rect 137150 685220 137240 685460
rect 137480 685220 137590 685460
rect 137830 685220 137920 685460
rect 138160 685220 138250 685460
rect 138490 685220 138580 685460
rect 138820 685220 138930 685460
rect 139170 685220 139260 685460
rect 139500 685220 139590 685460
rect 139830 685220 139920 685460
rect 140160 685220 140270 685460
rect 140510 685220 140600 685460
rect 140840 685220 140930 685460
rect 141170 685220 141260 685460
rect 141500 685220 141610 685460
rect 141850 685220 141940 685460
rect 142180 685220 142270 685460
rect 142510 685220 142600 685460
rect 142840 685220 142950 685460
rect 143190 685220 143280 685460
rect 143520 685220 143610 685460
rect 143850 685220 143940 685460
rect 144180 685220 144290 685460
rect 144530 685220 144550 685460
rect 133550 685110 144550 685220
rect 133550 684870 133570 685110
rect 133810 684870 133900 685110
rect 134140 684870 134230 685110
rect 134470 684870 134560 685110
rect 134800 684870 134910 685110
rect 135150 684870 135240 685110
rect 135480 684870 135570 685110
rect 135810 684870 135900 685110
rect 136140 684870 136250 685110
rect 136490 684870 136580 685110
rect 136820 684870 136910 685110
rect 137150 684870 137240 685110
rect 137480 684870 137590 685110
rect 137830 684870 137920 685110
rect 138160 684870 138250 685110
rect 138490 684870 138580 685110
rect 138820 684870 138930 685110
rect 139170 684870 139260 685110
rect 139500 684870 139590 685110
rect 139830 684870 139920 685110
rect 140160 684870 140270 685110
rect 140510 684870 140600 685110
rect 140840 684870 140930 685110
rect 141170 684870 141260 685110
rect 141500 684870 141610 685110
rect 141850 684870 141940 685110
rect 142180 684870 142270 685110
rect 142510 684870 142600 685110
rect 142840 684870 142950 685110
rect 143190 684870 143280 685110
rect 143520 684870 143610 685110
rect 143850 684870 143940 685110
rect 144180 684870 144290 685110
rect 144530 684870 144550 685110
rect 133550 684780 144550 684870
rect 133550 684540 133570 684780
rect 133810 684540 133900 684780
rect 134140 684540 134230 684780
rect 134470 684540 134560 684780
rect 134800 684540 134910 684780
rect 135150 684540 135240 684780
rect 135480 684540 135570 684780
rect 135810 684540 135900 684780
rect 136140 684540 136250 684780
rect 136490 684540 136580 684780
rect 136820 684540 136910 684780
rect 137150 684540 137240 684780
rect 137480 684540 137590 684780
rect 137830 684540 137920 684780
rect 138160 684540 138250 684780
rect 138490 684540 138580 684780
rect 138820 684540 138930 684780
rect 139170 684540 139260 684780
rect 139500 684540 139590 684780
rect 139830 684540 139920 684780
rect 140160 684540 140270 684780
rect 140510 684540 140600 684780
rect 140840 684540 140930 684780
rect 141170 684540 141260 684780
rect 141500 684540 141610 684780
rect 141850 684540 141940 684780
rect 142180 684540 142270 684780
rect 142510 684540 142600 684780
rect 142840 684540 142950 684780
rect 143190 684540 143280 684780
rect 143520 684540 143610 684780
rect 143850 684540 143940 684780
rect 144180 684540 144290 684780
rect 144530 684540 144550 684780
rect 133550 684450 144550 684540
rect 133550 684210 133570 684450
rect 133810 684210 133900 684450
rect 134140 684210 134230 684450
rect 134470 684210 134560 684450
rect 134800 684210 134910 684450
rect 135150 684210 135240 684450
rect 135480 684210 135570 684450
rect 135810 684210 135900 684450
rect 136140 684210 136250 684450
rect 136490 684210 136580 684450
rect 136820 684210 136910 684450
rect 137150 684210 137240 684450
rect 137480 684210 137590 684450
rect 137830 684210 137920 684450
rect 138160 684210 138250 684450
rect 138490 684210 138580 684450
rect 138820 684210 138930 684450
rect 139170 684210 139260 684450
rect 139500 684210 139590 684450
rect 139830 684210 139920 684450
rect 140160 684210 140270 684450
rect 140510 684210 140600 684450
rect 140840 684210 140930 684450
rect 141170 684210 141260 684450
rect 141500 684210 141610 684450
rect 141850 684210 141940 684450
rect 142180 684210 142270 684450
rect 142510 684210 142600 684450
rect 142840 684210 142950 684450
rect 143190 684210 143280 684450
rect 143520 684210 143610 684450
rect 143850 684210 143940 684450
rect 144180 684210 144290 684450
rect 144530 684210 144550 684450
rect 133550 684120 144550 684210
rect 133550 683880 133570 684120
rect 133810 683880 133900 684120
rect 134140 683880 134230 684120
rect 134470 683880 134560 684120
rect 134800 683880 134910 684120
rect 135150 683880 135240 684120
rect 135480 683880 135570 684120
rect 135810 683880 135900 684120
rect 136140 683880 136250 684120
rect 136490 683880 136580 684120
rect 136820 683880 136910 684120
rect 137150 683880 137240 684120
rect 137480 683880 137590 684120
rect 137830 683880 137920 684120
rect 138160 683880 138250 684120
rect 138490 683880 138580 684120
rect 138820 683880 138930 684120
rect 139170 683880 139260 684120
rect 139500 683880 139590 684120
rect 139830 683880 139920 684120
rect 140160 683880 140270 684120
rect 140510 683880 140600 684120
rect 140840 683880 140930 684120
rect 141170 683880 141260 684120
rect 141500 683880 141610 684120
rect 141850 683880 141940 684120
rect 142180 683880 142270 684120
rect 142510 683880 142600 684120
rect 142840 683880 142950 684120
rect 143190 683880 143280 684120
rect 143520 683880 143610 684120
rect 143850 683880 143940 684120
rect 144180 683880 144290 684120
rect 144530 683880 144550 684120
rect 133550 683860 144550 683880
rect 144930 694840 155930 694860
rect 144930 694600 144950 694840
rect 145190 694600 145280 694840
rect 145520 694600 145610 694840
rect 145850 694600 145940 694840
rect 146180 694600 146290 694840
rect 146530 694600 146620 694840
rect 146860 694600 146950 694840
rect 147190 694600 147280 694840
rect 147520 694600 147630 694840
rect 147870 694600 147960 694840
rect 148200 694600 148290 694840
rect 148530 694600 148620 694840
rect 148860 694600 148970 694840
rect 149210 694600 149300 694840
rect 149540 694600 149630 694840
rect 149870 694600 149960 694840
rect 150200 694600 150310 694840
rect 150550 694600 150640 694840
rect 150880 694600 150970 694840
rect 151210 694600 151300 694840
rect 151540 694600 151650 694840
rect 151890 694600 151980 694840
rect 152220 694600 152310 694840
rect 152550 694600 152640 694840
rect 152880 694600 152990 694840
rect 153230 694600 153320 694840
rect 153560 694600 153650 694840
rect 153890 694600 153980 694840
rect 154220 694600 154330 694840
rect 154570 694600 154660 694840
rect 154900 694600 154990 694840
rect 155230 694600 155320 694840
rect 155560 694600 155670 694840
rect 155910 694600 155930 694840
rect 144930 694490 155930 694600
rect 144930 694250 144950 694490
rect 145190 694250 145280 694490
rect 145520 694250 145610 694490
rect 145850 694250 145940 694490
rect 146180 694250 146290 694490
rect 146530 694250 146620 694490
rect 146860 694250 146950 694490
rect 147190 694250 147280 694490
rect 147520 694250 147630 694490
rect 147870 694250 147960 694490
rect 148200 694250 148290 694490
rect 148530 694250 148620 694490
rect 148860 694250 148970 694490
rect 149210 694250 149300 694490
rect 149540 694250 149630 694490
rect 149870 694250 149960 694490
rect 150200 694250 150310 694490
rect 150550 694250 150640 694490
rect 150880 694250 150970 694490
rect 151210 694250 151300 694490
rect 151540 694250 151650 694490
rect 151890 694250 151980 694490
rect 152220 694250 152310 694490
rect 152550 694250 152640 694490
rect 152880 694250 152990 694490
rect 153230 694250 153320 694490
rect 153560 694250 153650 694490
rect 153890 694250 153980 694490
rect 154220 694250 154330 694490
rect 154570 694250 154660 694490
rect 154900 694250 154990 694490
rect 155230 694250 155320 694490
rect 155560 694250 155670 694490
rect 155910 694250 155930 694490
rect 144930 694160 155930 694250
rect 144930 693920 144950 694160
rect 145190 693920 145280 694160
rect 145520 693920 145610 694160
rect 145850 693920 145940 694160
rect 146180 693920 146290 694160
rect 146530 693920 146620 694160
rect 146860 693920 146950 694160
rect 147190 693920 147280 694160
rect 147520 693920 147630 694160
rect 147870 693920 147960 694160
rect 148200 693920 148290 694160
rect 148530 693920 148620 694160
rect 148860 693920 148970 694160
rect 149210 693920 149300 694160
rect 149540 693920 149630 694160
rect 149870 693920 149960 694160
rect 150200 693920 150310 694160
rect 150550 693920 150640 694160
rect 150880 693920 150970 694160
rect 151210 693920 151300 694160
rect 151540 693920 151650 694160
rect 151890 693920 151980 694160
rect 152220 693920 152310 694160
rect 152550 693920 152640 694160
rect 152880 693920 152990 694160
rect 153230 693920 153320 694160
rect 153560 693920 153650 694160
rect 153890 693920 153980 694160
rect 154220 693920 154330 694160
rect 154570 693920 154660 694160
rect 154900 693920 154990 694160
rect 155230 693920 155320 694160
rect 155560 693920 155670 694160
rect 155910 693920 155930 694160
rect 144930 693830 155930 693920
rect 144930 693590 144950 693830
rect 145190 693590 145280 693830
rect 145520 693590 145610 693830
rect 145850 693590 145940 693830
rect 146180 693590 146290 693830
rect 146530 693590 146620 693830
rect 146860 693590 146950 693830
rect 147190 693590 147280 693830
rect 147520 693590 147630 693830
rect 147870 693590 147960 693830
rect 148200 693590 148290 693830
rect 148530 693590 148620 693830
rect 148860 693590 148970 693830
rect 149210 693590 149300 693830
rect 149540 693590 149630 693830
rect 149870 693590 149960 693830
rect 150200 693590 150310 693830
rect 150550 693590 150640 693830
rect 150880 693590 150970 693830
rect 151210 693590 151300 693830
rect 151540 693590 151650 693830
rect 151890 693590 151980 693830
rect 152220 693590 152310 693830
rect 152550 693590 152640 693830
rect 152880 693590 152990 693830
rect 153230 693590 153320 693830
rect 153560 693590 153650 693830
rect 153890 693590 153980 693830
rect 154220 693590 154330 693830
rect 154570 693590 154660 693830
rect 154900 693590 154990 693830
rect 155230 693590 155320 693830
rect 155560 693590 155670 693830
rect 155910 693590 155930 693830
rect 144930 693500 155930 693590
rect 144930 693260 144950 693500
rect 145190 693260 145280 693500
rect 145520 693260 145610 693500
rect 145850 693260 145940 693500
rect 146180 693260 146290 693500
rect 146530 693260 146620 693500
rect 146860 693260 146950 693500
rect 147190 693260 147280 693500
rect 147520 693260 147630 693500
rect 147870 693260 147960 693500
rect 148200 693260 148290 693500
rect 148530 693260 148620 693500
rect 148860 693260 148970 693500
rect 149210 693260 149300 693500
rect 149540 693260 149630 693500
rect 149870 693260 149960 693500
rect 150200 693260 150310 693500
rect 150550 693260 150640 693500
rect 150880 693260 150970 693500
rect 151210 693260 151300 693500
rect 151540 693260 151650 693500
rect 151890 693260 151980 693500
rect 152220 693260 152310 693500
rect 152550 693260 152640 693500
rect 152880 693260 152990 693500
rect 153230 693260 153320 693500
rect 153560 693260 153650 693500
rect 153890 693260 153980 693500
rect 154220 693260 154330 693500
rect 154570 693260 154660 693500
rect 154900 693260 154990 693500
rect 155230 693260 155320 693500
rect 155560 693260 155670 693500
rect 155910 693260 155930 693500
rect 144930 693150 155930 693260
rect 144930 692910 144950 693150
rect 145190 692910 145280 693150
rect 145520 692910 145610 693150
rect 145850 692910 145940 693150
rect 146180 692910 146290 693150
rect 146530 692910 146620 693150
rect 146860 692910 146950 693150
rect 147190 692910 147280 693150
rect 147520 692910 147630 693150
rect 147870 692910 147960 693150
rect 148200 692910 148290 693150
rect 148530 692910 148620 693150
rect 148860 692910 148970 693150
rect 149210 692910 149300 693150
rect 149540 692910 149630 693150
rect 149870 692910 149960 693150
rect 150200 692910 150310 693150
rect 150550 692910 150640 693150
rect 150880 692910 150970 693150
rect 151210 692910 151300 693150
rect 151540 692910 151650 693150
rect 151890 692910 151980 693150
rect 152220 692910 152310 693150
rect 152550 692910 152640 693150
rect 152880 692910 152990 693150
rect 153230 692910 153320 693150
rect 153560 692910 153650 693150
rect 153890 692910 153980 693150
rect 154220 692910 154330 693150
rect 154570 692910 154660 693150
rect 154900 692910 154990 693150
rect 155230 692910 155320 693150
rect 155560 692910 155670 693150
rect 155910 692910 155930 693150
rect 144930 692820 155930 692910
rect 144930 692580 144950 692820
rect 145190 692580 145280 692820
rect 145520 692580 145610 692820
rect 145850 692580 145940 692820
rect 146180 692580 146290 692820
rect 146530 692580 146620 692820
rect 146860 692580 146950 692820
rect 147190 692580 147280 692820
rect 147520 692580 147630 692820
rect 147870 692580 147960 692820
rect 148200 692580 148290 692820
rect 148530 692580 148620 692820
rect 148860 692580 148970 692820
rect 149210 692580 149300 692820
rect 149540 692580 149630 692820
rect 149870 692580 149960 692820
rect 150200 692580 150310 692820
rect 150550 692580 150640 692820
rect 150880 692580 150970 692820
rect 151210 692580 151300 692820
rect 151540 692580 151650 692820
rect 151890 692580 151980 692820
rect 152220 692580 152310 692820
rect 152550 692580 152640 692820
rect 152880 692580 152990 692820
rect 153230 692580 153320 692820
rect 153560 692580 153650 692820
rect 153890 692580 153980 692820
rect 154220 692580 154330 692820
rect 154570 692580 154660 692820
rect 154900 692580 154990 692820
rect 155230 692580 155320 692820
rect 155560 692580 155670 692820
rect 155910 692580 155930 692820
rect 144930 692490 155930 692580
rect 144930 692250 144950 692490
rect 145190 692250 145280 692490
rect 145520 692250 145610 692490
rect 145850 692250 145940 692490
rect 146180 692250 146290 692490
rect 146530 692250 146620 692490
rect 146860 692250 146950 692490
rect 147190 692250 147280 692490
rect 147520 692250 147630 692490
rect 147870 692250 147960 692490
rect 148200 692250 148290 692490
rect 148530 692250 148620 692490
rect 148860 692250 148970 692490
rect 149210 692250 149300 692490
rect 149540 692250 149630 692490
rect 149870 692250 149960 692490
rect 150200 692250 150310 692490
rect 150550 692250 150640 692490
rect 150880 692250 150970 692490
rect 151210 692250 151300 692490
rect 151540 692250 151650 692490
rect 151890 692250 151980 692490
rect 152220 692250 152310 692490
rect 152550 692250 152640 692490
rect 152880 692250 152990 692490
rect 153230 692250 153320 692490
rect 153560 692250 153650 692490
rect 153890 692250 153980 692490
rect 154220 692250 154330 692490
rect 154570 692250 154660 692490
rect 154900 692250 154990 692490
rect 155230 692250 155320 692490
rect 155560 692250 155670 692490
rect 155910 692250 155930 692490
rect 144930 692160 155930 692250
rect 144930 691920 144950 692160
rect 145190 691920 145280 692160
rect 145520 691920 145610 692160
rect 145850 691920 145940 692160
rect 146180 691920 146290 692160
rect 146530 691920 146620 692160
rect 146860 691920 146950 692160
rect 147190 691920 147280 692160
rect 147520 691920 147630 692160
rect 147870 691920 147960 692160
rect 148200 691920 148290 692160
rect 148530 691920 148620 692160
rect 148860 691920 148970 692160
rect 149210 691920 149300 692160
rect 149540 691920 149630 692160
rect 149870 691920 149960 692160
rect 150200 691920 150310 692160
rect 150550 691920 150640 692160
rect 150880 691920 150970 692160
rect 151210 691920 151300 692160
rect 151540 691920 151650 692160
rect 151890 691920 151980 692160
rect 152220 691920 152310 692160
rect 152550 691920 152640 692160
rect 152880 691920 152990 692160
rect 153230 691920 153320 692160
rect 153560 691920 153650 692160
rect 153890 691920 153980 692160
rect 154220 691920 154330 692160
rect 154570 691920 154660 692160
rect 154900 691920 154990 692160
rect 155230 691920 155320 692160
rect 155560 691920 155670 692160
rect 155910 691920 155930 692160
rect 144930 691810 155930 691920
rect 144930 691570 144950 691810
rect 145190 691570 145280 691810
rect 145520 691570 145610 691810
rect 145850 691570 145940 691810
rect 146180 691570 146290 691810
rect 146530 691570 146620 691810
rect 146860 691570 146950 691810
rect 147190 691570 147280 691810
rect 147520 691570 147630 691810
rect 147870 691570 147960 691810
rect 148200 691570 148290 691810
rect 148530 691570 148620 691810
rect 148860 691570 148970 691810
rect 149210 691570 149300 691810
rect 149540 691570 149630 691810
rect 149870 691570 149960 691810
rect 150200 691570 150310 691810
rect 150550 691570 150640 691810
rect 150880 691570 150970 691810
rect 151210 691570 151300 691810
rect 151540 691570 151650 691810
rect 151890 691570 151980 691810
rect 152220 691570 152310 691810
rect 152550 691570 152640 691810
rect 152880 691570 152990 691810
rect 153230 691570 153320 691810
rect 153560 691570 153650 691810
rect 153890 691570 153980 691810
rect 154220 691570 154330 691810
rect 154570 691570 154660 691810
rect 154900 691570 154990 691810
rect 155230 691570 155320 691810
rect 155560 691570 155670 691810
rect 155910 691570 155930 691810
rect 144930 691480 155930 691570
rect 144930 691240 144950 691480
rect 145190 691240 145280 691480
rect 145520 691240 145610 691480
rect 145850 691240 145940 691480
rect 146180 691240 146290 691480
rect 146530 691240 146620 691480
rect 146860 691240 146950 691480
rect 147190 691240 147280 691480
rect 147520 691240 147630 691480
rect 147870 691240 147960 691480
rect 148200 691240 148290 691480
rect 148530 691240 148620 691480
rect 148860 691240 148970 691480
rect 149210 691240 149300 691480
rect 149540 691240 149630 691480
rect 149870 691240 149960 691480
rect 150200 691240 150310 691480
rect 150550 691240 150640 691480
rect 150880 691240 150970 691480
rect 151210 691240 151300 691480
rect 151540 691240 151650 691480
rect 151890 691240 151980 691480
rect 152220 691240 152310 691480
rect 152550 691240 152640 691480
rect 152880 691240 152990 691480
rect 153230 691240 153320 691480
rect 153560 691240 153650 691480
rect 153890 691240 153980 691480
rect 154220 691240 154330 691480
rect 154570 691240 154660 691480
rect 154900 691240 154990 691480
rect 155230 691240 155320 691480
rect 155560 691240 155670 691480
rect 155910 691240 155930 691480
rect 144930 691150 155930 691240
rect 144930 690910 144950 691150
rect 145190 690910 145280 691150
rect 145520 690910 145610 691150
rect 145850 690910 145940 691150
rect 146180 690910 146290 691150
rect 146530 690910 146620 691150
rect 146860 690910 146950 691150
rect 147190 690910 147280 691150
rect 147520 690910 147630 691150
rect 147870 690910 147960 691150
rect 148200 690910 148290 691150
rect 148530 690910 148620 691150
rect 148860 690910 148970 691150
rect 149210 690910 149300 691150
rect 149540 690910 149630 691150
rect 149870 690910 149960 691150
rect 150200 690910 150310 691150
rect 150550 690910 150640 691150
rect 150880 690910 150970 691150
rect 151210 690910 151300 691150
rect 151540 690910 151650 691150
rect 151890 690910 151980 691150
rect 152220 690910 152310 691150
rect 152550 690910 152640 691150
rect 152880 690910 152990 691150
rect 153230 690910 153320 691150
rect 153560 690910 153650 691150
rect 153890 690910 153980 691150
rect 154220 690910 154330 691150
rect 154570 690910 154660 691150
rect 154900 690910 154990 691150
rect 155230 690910 155320 691150
rect 155560 690910 155670 691150
rect 155910 690910 155930 691150
rect 144930 690820 155930 690910
rect 144930 690580 144950 690820
rect 145190 690580 145280 690820
rect 145520 690580 145610 690820
rect 145850 690580 145940 690820
rect 146180 690580 146290 690820
rect 146530 690580 146620 690820
rect 146860 690580 146950 690820
rect 147190 690580 147280 690820
rect 147520 690580 147630 690820
rect 147870 690580 147960 690820
rect 148200 690580 148290 690820
rect 148530 690580 148620 690820
rect 148860 690580 148970 690820
rect 149210 690580 149300 690820
rect 149540 690580 149630 690820
rect 149870 690580 149960 690820
rect 150200 690580 150310 690820
rect 150550 690580 150640 690820
rect 150880 690580 150970 690820
rect 151210 690580 151300 690820
rect 151540 690580 151650 690820
rect 151890 690580 151980 690820
rect 152220 690580 152310 690820
rect 152550 690580 152640 690820
rect 152880 690580 152990 690820
rect 153230 690580 153320 690820
rect 153560 690580 153650 690820
rect 153890 690580 153980 690820
rect 154220 690580 154330 690820
rect 154570 690580 154660 690820
rect 154900 690580 154990 690820
rect 155230 690580 155320 690820
rect 155560 690580 155670 690820
rect 155910 690580 155930 690820
rect 144930 690470 155930 690580
rect 144930 690230 144950 690470
rect 145190 690230 145280 690470
rect 145520 690230 145610 690470
rect 145850 690230 145940 690470
rect 146180 690230 146290 690470
rect 146530 690230 146620 690470
rect 146860 690230 146950 690470
rect 147190 690230 147280 690470
rect 147520 690230 147630 690470
rect 147870 690230 147960 690470
rect 148200 690230 148290 690470
rect 148530 690230 148620 690470
rect 148860 690230 148970 690470
rect 149210 690230 149300 690470
rect 149540 690230 149630 690470
rect 149870 690230 149960 690470
rect 150200 690230 150310 690470
rect 150550 690230 150640 690470
rect 150880 690230 150970 690470
rect 151210 690230 151300 690470
rect 151540 690230 151650 690470
rect 151890 690230 151980 690470
rect 152220 690230 152310 690470
rect 152550 690230 152640 690470
rect 152880 690230 152990 690470
rect 153230 690230 153320 690470
rect 153560 690230 153650 690470
rect 153890 690230 153980 690470
rect 154220 690230 154330 690470
rect 154570 690230 154660 690470
rect 154900 690230 154990 690470
rect 155230 690230 155320 690470
rect 155560 690230 155670 690470
rect 155910 690230 155930 690470
rect 144930 690140 155930 690230
rect 144930 689900 144950 690140
rect 145190 689900 145280 690140
rect 145520 689900 145610 690140
rect 145850 689900 145940 690140
rect 146180 689900 146290 690140
rect 146530 689900 146620 690140
rect 146860 689900 146950 690140
rect 147190 689900 147280 690140
rect 147520 689900 147630 690140
rect 147870 689900 147960 690140
rect 148200 689900 148290 690140
rect 148530 689900 148620 690140
rect 148860 689900 148970 690140
rect 149210 689900 149300 690140
rect 149540 689900 149630 690140
rect 149870 689900 149960 690140
rect 150200 689900 150310 690140
rect 150550 689900 150640 690140
rect 150880 689900 150970 690140
rect 151210 689900 151300 690140
rect 151540 689900 151650 690140
rect 151890 689900 151980 690140
rect 152220 689900 152310 690140
rect 152550 689900 152640 690140
rect 152880 689900 152990 690140
rect 153230 689900 153320 690140
rect 153560 689900 153650 690140
rect 153890 689900 153980 690140
rect 154220 689900 154330 690140
rect 154570 689900 154660 690140
rect 154900 689900 154990 690140
rect 155230 689900 155320 690140
rect 155560 689900 155670 690140
rect 155910 689900 155930 690140
rect 144930 689810 155930 689900
rect 144930 689570 144950 689810
rect 145190 689570 145280 689810
rect 145520 689570 145610 689810
rect 145850 689570 145940 689810
rect 146180 689570 146290 689810
rect 146530 689570 146620 689810
rect 146860 689570 146950 689810
rect 147190 689570 147280 689810
rect 147520 689570 147630 689810
rect 147870 689570 147960 689810
rect 148200 689570 148290 689810
rect 148530 689570 148620 689810
rect 148860 689570 148970 689810
rect 149210 689570 149300 689810
rect 149540 689570 149630 689810
rect 149870 689570 149960 689810
rect 150200 689570 150310 689810
rect 150550 689570 150640 689810
rect 150880 689570 150970 689810
rect 151210 689570 151300 689810
rect 151540 689570 151650 689810
rect 151890 689570 151980 689810
rect 152220 689570 152310 689810
rect 152550 689570 152640 689810
rect 152880 689570 152990 689810
rect 153230 689570 153320 689810
rect 153560 689570 153650 689810
rect 153890 689570 153980 689810
rect 154220 689570 154330 689810
rect 154570 689570 154660 689810
rect 154900 689570 154990 689810
rect 155230 689570 155320 689810
rect 155560 689570 155670 689810
rect 155910 689570 155930 689810
rect 144930 689480 155930 689570
rect 144930 689240 144950 689480
rect 145190 689240 145280 689480
rect 145520 689240 145610 689480
rect 145850 689240 145940 689480
rect 146180 689240 146290 689480
rect 146530 689240 146620 689480
rect 146860 689240 146950 689480
rect 147190 689240 147280 689480
rect 147520 689240 147630 689480
rect 147870 689240 147960 689480
rect 148200 689240 148290 689480
rect 148530 689240 148620 689480
rect 148860 689240 148970 689480
rect 149210 689240 149300 689480
rect 149540 689240 149630 689480
rect 149870 689240 149960 689480
rect 150200 689240 150310 689480
rect 150550 689240 150640 689480
rect 150880 689240 150970 689480
rect 151210 689240 151300 689480
rect 151540 689240 151650 689480
rect 151890 689240 151980 689480
rect 152220 689240 152310 689480
rect 152550 689240 152640 689480
rect 152880 689240 152990 689480
rect 153230 689240 153320 689480
rect 153560 689240 153650 689480
rect 153890 689240 153980 689480
rect 154220 689240 154330 689480
rect 154570 689240 154660 689480
rect 154900 689240 154990 689480
rect 155230 689240 155320 689480
rect 155560 689240 155670 689480
rect 155910 689240 155930 689480
rect 144930 689130 155930 689240
rect 144930 688890 144950 689130
rect 145190 688890 145280 689130
rect 145520 688890 145610 689130
rect 145850 688890 145940 689130
rect 146180 688890 146290 689130
rect 146530 688890 146620 689130
rect 146860 688890 146950 689130
rect 147190 688890 147280 689130
rect 147520 688890 147630 689130
rect 147870 688890 147960 689130
rect 148200 688890 148290 689130
rect 148530 688890 148620 689130
rect 148860 688890 148970 689130
rect 149210 688890 149300 689130
rect 149540 688890 149630 689130
rect 149870 688890 149960 689130
rect 150200 688890 150310 689130
rect 150550 688890 150640 689130
rect 150880 688890 150970 689130
rect 151210 688890 151300 689130
rect 151540 688890 151650 689130
rect 151890 688890 151980 689130
rect 152220 688890 152310 689130
rect 152550 688890 152640 689130
rect 152880 688890 152990 689130
rect 153230 688890 153320 689130
rect 153560 688890 153650 689130
rect 153890 688890 153980 689130
rect 154220 688890 154330 689130
rect 154570 688890 154660 689130
rect 154900 688890 154990 689130
rect 155230 688890 155320 689130
rect 155560 688890 155670 689130
rect 155910 688890 155930 689130
rect 144930 688800 155930 688890
rect 144930 688560 144950 688800
rect 145190 688560 145280 688800
rect 145520 688560 145610 688800
rect 145850 688560 145940 688800
rect 146180 688560 146290 688800
rect 146530 688560 146620 688800
rect 146860 688560 146950 688800
rect 147190 688560 147280 688800
rect 147520 688560 147630 688800
rect 147870 688560 147960 688800
rect 148200 688560 148290 688800
rect 148530 688560 148620 688800
rect 148860 688560 148970 688800
rect 149210 688560 149300 688800
rect 149540 688560 149630 688800
rect 149870 688560 149960 688800
rect 150200 688560 150310 688800
rect 150550 688560 150640 688800
rect 150880 688560 150970 688800
rect 151210 688560 151300 688800
rect 151540 688560 151650 688800
rect 151890 688560 151980 688800
rect 152220 688560 152310 688800
rect 152550 688560 152640 688800
rect 152880 688560 152990 688800
rect 153230 688560 153320 688800
rect 153560 688560 153650 688800
rect 153890 688560 153980 688800
rect 154220 688560 154330 688800
rect 154570 688560 154660 688800
rect 154900 688560 154990 688800
rect 155230 688560 155320 688800
rect 155560 688560 155670 688800
rect 155910 688560 155930 688800
rect 144930 688470 155930 688560
rect 144930 688230 144950 688470
rect 145190 688230 145280 688470
rect 145520 688230 145610 688470
rect 145850 688230 145940 688470
rect 146180 688230 146290 688470
rect 146530 688230 146620 688470
rect 146860 688230 146950 688470
rect 147190 688230 147280 688470
rect 147520 688230 147630 688470
rect 147870 688230 147960 688470
rect 148200 688230 148290 688470
rect 148530 688230 148620 688470
rect 148860 688230 148970 688470
rect 149210 688230 149300 688470
rect 149540 688230 149630 688470
rect 149870 688230 149960 688470
rect 150200 688230 150310 688470
rect 150550 688230 150640 688470
rect 150880 688230 150970 688470
rect 151210 688230 151300 688470
rect 151540 688230 151650 688470
rect 151890 688230 151980 688470
rect 152220 688230 152310 688470
rect 152550 688230 152640 688470
rect 152880 688230 152990 688470
rect 153230 688230 153320 688470
rect 153560 688230 153650 688470
rect 153890 688230 153980 688470
rect 154220 688230 154330 688470
rect 154570 688230 154660 688470
rect 154900 688230 154990 688470
rect 155230 688230 155320 688470
rect 155560 688230 155670 688470
rect 155910 688230 155930 688470
rect 144930 688140 155930 688230
rect 144930 687900 144950 688140
rect 145190 687900 145280 688140
rect 145520 687900 145610 688140
rect 145850 687900 145940 688140
rect 146180 687900 146290 688140
rect 146530 687900 146620 688140
rect 146860 687900 146950 688140
rect 147190 687900 147280 688140
rect 147520 687900 147630 688140
rect 147870 687900 147960 688140
rect 148200 687900 148290 688140
rect 148530 687900 148620 688140
rect 148860 687900 148970 688140
rect 149210 687900 149300 688140
rect 149540 687900 149630 688140
rect 149870 687900 149960 688140
rect 150200 687900 150310 688140
rect 150550 687900 150640 688140
rect 150880 687900 150970 688140
rect 151210 687900 151300 688140
rect 151540 687900 151650 688140
rect 151890 687900 151980 688140
rect 152220 687900 152310 688140
rect 152550 687900 152640 688140
rect 152880 687900 152990 688140
rect 153230 687900 153320 688140
rect 153560 687900 153650 688140
rect 153890 687900 153980 688140
rect 154220 687900 154330 688140
rect 154570 687900 154660 688140
rect 154900 687900 154990 688140
rect 155230 687900 155320 688140
rect 155560 687900 155670 688140
rect 155910 687900 155930 688140
rect 144930 687790 155930 687900
rect 144930 687550 144950 687790
rect 145190 687550 145280 687790
rect 145520 687550 145610 687790
rect 145850 687550 145940 687790
rect 146180 687550 146290 687790
rect 146530 687550 146620 687790
rect 146860 687550 146950 687790
rect 147190 687550 147280 687790
rect 147520 687550 147630 687790
rect 147870 687550 147960 687790
rect 148200 687550 148290 687790
rect 148530 687550 148620 687790
rect 148860 687550 148970 687790
rect 149210 687550 149300 687790
rect 149540 687550 149630 687790
rect 149870 687550 149960 687790
rect 150200 687550 150310 687790
rect 150550 687550 150640 687790
rect 150880 687550 150970 687790
rect 151210 687550 151300 687790
rect 151540 687550 151650 687790
rect 151890 687550 151980 687790
rect 152220 687550 152310 687790
rect 152550 687550 152640 687790
rect 152880 687550 152990 687790
rect 153230 687550 153320 687790
rect 153560 687550 153650 687790
rect 153890 687550 153980 687790
rect 154220 687550 154330 687790
rect 154570 687550 154660 687790
rect 154900 687550 154990 687790
rect 155230 687550 155320 687790
rect 155560 687550 155670 687790
rect 155910 687550 155930 687790
rect 144930 687460 155930 687550
rect 144930 687220 144950 687460
rect 145190 687220 145280 687460
rect 145520 687220 145610 687460
rect 145850 687220 145940 687460
rect 146180 687220 146290 687460
rect 146530 687220 146620 687460
rect 146860 687220 146950 687460
rect 147190 687220 147280 687460
rect 147520 687220 147630 687460
rect 147870 687220 147960 687460
rect 148200 687220 148290 687460
rect 148530 687220 148620 687460
rect 148860 687220 148970 687460
rect 149210 687220 149300 687460
rect 149540 687220 149630 687460
rect 149870 687220 149960 687460
rect 150200 687220 150310 687460
rect 150550 687220 150640 687460
rect 150880 687220 150970 687460
rect 151210 687220 151300 687460
rect 151540 687220 151650 687460
rect 151890 687220 151980 687460
rect 152220 687220 152310 687460
rect 152550 687220 152640 687460
rect 152880 687220 152990 687460
rect 153230 687220 153320 687460
rect 153560 687220 153650 687460
rect 153890 687220 153980 687460
rect 154220 687220 154330 687460
rect 154570 687220 154660 687460
rect 154900 687220 154990 687460
rect 155230 687220 155320 687460
rect 155560 687220 155670 687460
rect 155910 687220 155930 687460
rect 144930 687130 155930 687220
rect 144930 686890 144950 687130
rect 145190 686890 145280 687130
rect 145520 686890 145610 687130
rect 145850 686890 145940 687130
rect 146180 686890 146290 687130
rect 146530 686890 146620 687130
rect 146860 686890 146950 687130
rect 147190 686890 147280 687130
rect 147520 686890 147630 687130
rect 147870 686890 147960 687130
rect 148200 686890 148290 687130
rect 148530 686890 148620 687130
rect 148860 686890 148970 687130
rect 149210 686890 149300 687130
rect 149540 686890 149630 687130
rect 149870 686890 149960 687130
rect 150200 686890 150310 687130
rect 150550 686890 150640 687130
rect 150880 686890 150970 687130
rect 151210 686890 151300 687130
rect 151540 686890 151650 687130
rect 151890 686890 151980 687130
rect 152220 686890 152310 687130
rect 152550 686890 152640 687130
rect 152880 686890 152990 687130
rect 153230 686890 153320 687130
rect 153560 686890 153650 687130
rect 153890 686890 153980 687130
rect 154220 686890 154330 687130
rect 154570 686890 154660 687130
rect 154900 686890 154990 687130
rect 155230 686890 155320 687130
rect 155560 686890 155670 687130
rect 155910 686890 155930 687130
rect 144930 686800 155930 686890
rect 144930 686560 144950 686800
rect 145190 686560 145280 686800
rect 145520 686560 145610 686800
rect 145850 686560 145940 686800
rect 146180 686560 146290 686800
rect 146530 686560 146620 686800
rect 146860 686560 146950 686800
rect 147190 686560 147280 686800
rect 147520 686560 147630 686800
rect 147870 686560 147960 686800
rect 148200 686560 148290 686800
rect 148530 686560 148620 686800
rect 148860 686560 148970 686800
rect 149210 686560 149300 686800
rect 149540 686560 149630 686800
rect 149870 686560 149960 686800
rect 150200 686560 150310 686800
rect 150550 686560 150640 686800
rect 150880 686560 150970 686800
rect 151210 686560 151300 686800
rect 151540 686560 151650 686800
rect 151890 686560 151980 686800
rect 152220 686560 152310 686800
rect 152550 686560 152640 686800
rect 152880 686560 152990 686800
rect 153230 686560 153320 686800
rect 153560 686560 153650 686800
rect 153890 686560 153980 686800
rect 154220 686560 154330 686800
rect 154570 686560 154660 686800
rect 154900 686560 154990 686800
rect 155230 686560 155320 686800
rect 155560 686560 155670 686800
rect 155910 686560 155930 686800
rect 144930 686450 155930 686560
rect 144930 686210 144950 686450
rect 145190 686210 145280 686450
rect 145520 686210 145610 686450
rect 145850 686210 145940 686450
rect 146180 686210 146290 686450
rect 146530 686210 146620 686450
rect 146860 686210 146950 686450
rect 147190 686210 147280 686450
rect 147520 686210 147630 686450
rect 147870 686210 147960 686450
rect 148200 686210 148290 686450
rect 148530 686210 148620 686450
rect 148860 686210 148970 686450
rect 149210 686210 149300 686450
rect 149540 686210 149630 686450
rect 149870 686210 149960 686450
rect 150200 686210 150310 686450
rect 150550 686210 150640 686450
rect 150880 686210 150970 686450
rect 151210 686210 151300 686450
rect 151540 686210 151650 686450
rect 151890 686210 151980 686450
rect 152220 686210 152310 686450
rect 152550 686210 152640 686450
rect 152880 686210 152990 686450
rect 153230 686210 153320 686450
rect 153560 686210 153650 686450
rect 153890 686210 153980 686450
rect 154220 686210 154330 686450
rect 154570 686210 154660 686450
rect 154900 686210 154990 686450
rect 155230 686210 155320 686450
rect 155560 686210 155670 686450
rect 155910 686210 155930 686450
rect 144930 686120 155930 686210
rect 144930 685880 144950 686120
rect 145190 685880 145280 686120
rect 145520 685880 145610 686120
rect 145850 685880 145940 686120
rect 146180 685880 146290 686120
rect 146530 685880 146620 686120
rect 146860 685880 146950 686120
rect 147190 685880 147280 686120
rect 147520 685880 147630 686120
rect 147870 685880 147960 686120
rect 148200 685880 148290 686120
rect 148530 685880 148620 686120
rect 148860 685880 148970 686120
rect 149210 685880 149300 686120
rect 149540 685880 149630 686120
rect 149870 685880 149960 686120
rect 150200 685880 150310 686120
rect 150550 685880 150640 686120
rect 150880 685880 150970 686120
rect 151210 685880 151300 686120
rect 151540 685880 151650 686120
rect 151890 685880 151980 686120
rect 152220 685880 152310 686120
rect 152550 685880 152640 686120
rect 152880 685880 152990 686120
rect 153230 685880 153320 686120
rect 153560 685880 153650 686120
rect 153890 685880 153980 686120
rect 154220 685880 154330 686120
rect 154570 685880 154660 686120
rect 154900 685880 154990 686120
rect 155230 685880 155320 686120
rect 155560 685880 155670 686120
rect 155910 685880 155930 686120
rect 144930 685790 155930 685880
rect 144930 685550 144950 685790
rect 145190 685550 145280 685790
rect 145520 685550 145610 685790
rect 145850 685550 145940 685790
rect 146180 685550 146290 685790
rect 146530 685550 146620 685790
rect 146860 685550 146950 685790
rect 147190 685550 147280 685790
rect 147520 685550 147630 685790
rect 147870 685550 147960 685790
rect 148200 685550 148290 685790
rect 148530 685550 148620 685790
rect 148860 685550 148970 685790
rect 149210 685550 149300 685790
rect 149540 685550 149630 685790
rect 149870 685550 149960 685790
rect 150200 685550 150310 685790
rect 150550 685550 150640 685790
rect 150880 685550 150970 685790
rect 151210 685550 151300 685790
rect 151540 685550 151650 685790
rect 151890 685550 151980 685790
rect 152220 685550 152310 685790
rect 152550 685550 152640 685790
rect 152880 685550 152990 685790
rect 153230 685550 153320 685790
rect 153560 685550 153650 685790
rect 153890 685550 153980 685790
rect 154220 685550 154330 685790
rect 154570 685550 154660 685790
rect 154900 685550 154990 685790
rect 155230 685550 155320 685790
rect 155560 685550 155670 685790
rect 155910 685550 155930 685790
rect 144930 685460 155930 685550
rect 144930 685220 144950 685460
rect 145190 685220 145280 685460
rect 145520 685220 145610 685460
rect 145850 685220 145940 685460
rect 146180 685220 146290 685460
rect 146530 685220 146620 685460
rect 146860 685220 146950 685460
rect 147190 685220 147280 685460
rect 147520 685220 147630 685460
rect 147870 685220 147960 685460
rect 148200 685220 148290 685460
rect 148530 685220 148620 685460
rect 148860 685220 148970 685460
rect 149210 685220 149300 685460
rect 149540 685220 149630 685460
rect 149870 685220 149960 685460
rect 150200 685220 150310 685460
rect 150550 685220 150640 685460
rect 150880 685220 150970 685460
rect 151210 685220 151300 685460
rect 151540 685220 151650 685460
rect 151890 685220 151980 685460
rect 152220 685220 152310 685460
rect 152550 685220 152640 685460
rect 152880 685220 152990 685460
rect 153230 685220 153320 685460
rect 153560 685220 153650 685460
rect 153890 685220 153980 685460
rect 154220 685220 154330 685460
rect 154570 685220 154660 685460
rect 154900 685220 154990 685460
rect 155230 685220 155320 685460
rect 155560 685220 155670 685460
rect 155910 685220 155930 685460
rect 144930 685110 155930 685220
rect 144930 684870 144950 685110
rect 145190 684870 145280 685110
rect 145520 684870 145610 685110
rect 145850 684870 145940 685110
rect 146180 684870 146290 685110
rect 146530 684870 146620 685110
rect 146860 684870 146950 685110
rect 147190 684870 147280 685110
rect 147520 684870 147630 685110
rect 147870 684870 147960 685110
rect 148200 684870 148290 685110
rect 148530 684870 148620 685110
rect 148860 684870 148970 685110
rect 149210 684870 149300 685110
rect 149540 684870 149630 685110
rect 149870 684870 149960 685110
rect 150200 684870 150310 685110
rect 150550 684870 150640 685110
rect 150880 684870 150970 685110
rect 151210 684870 151300 685110
rect 151540 684870 151650 685110
rect 151890 684870 151980 685110
rect 152220 684870 152310 685110
rect 152550 684870 152640 685110
rect 152880 684870 152990 685110
rect 153230 684870 153320 685110
rect 153560 684870 153650 685110
rect 153890 684870 153980 685110
rect 154220 684870 154330 685110
rect 154570 684870 154660 685110
rect 154900 684870 154990 685110
rect 155230 684870 155320 685110
rect 155560 684870 155670 685110
rect 155910 684870 155930 685110
rect 144930 684780 155930 684870
rect 144930 684540 144950 684780
rect 145190 684540 145280 684780
rect 145520 684540 145610 684780
rect 145850 684540 145940 684780
rect 146180 684540 146290 684780
rect 146530 684540 146620 684780
rect 146860 684540 146950 684780
rect 147190 684540 147280 684780
rect 147520 684540 147630 684780
rect 147870 684540 147960 684780
rect 148200 684540 148290 684780
rect 148530 684540 148620 684780
rect 148860 684540 148970 684780
rect 149210 684540 149300 684780
rect 149540 684540 149630 684780
rect 149870 684540 149960 684780
rect 150200 684540 150310 684780
rect 150550 684540 150640 684780
rect 150880 684540 150970 684780
rect 151210 684540 151300 684780
rect 151540 684540 151650 684780
rect 151890 684540 151980 684780
rect 152220 684540 152310 684780
rect 152550 684540 152640 684780
rect 152880 684540 152990 684780
rect 153230 684540 153320 684780
rect 153560 684540 153650 684780
rect 153890 684540 153980 684780
rect 154220 684540 154330 684780
rect 154570 684540 154660 684780
rect 154900 684540 154990 684780
rect 155230 684540 155320 684780
rect 155560 684540 155670 684780
rect 155910 684540 155930 684780
rect 144930 684450 155930 684540
rect 144930 684210 144950 684450
rect 145190 684210 145280 684450
rect 145520 684210 145610 684450
rect 145850 684210 145940 684450
rect 146180 684210 146290 684450
rect 146530 684210 146620 684450
rect 146860 684210 146950 684450
rect 147190 684210 147280 684450
rect 147520 684210 147630 684450
rect 147870 684210 147960 684450
rect 148200 684210 148290 684450
rect 148530 684210 148620 684450
rect 148860 684210 148970 684450
rect 149210 684210 149300 684450
rect 149540 684210 149630 684450
rect 149870 684210 149960 684450
rect 150200 684210 150310 684450
rect 150550 684210 150640 684450
rect 150880 684210 150970 684450
rect 151210 684210 151300 684450
rect 151540 684210 151650 684450
rect 151890 684210 151980 684450
rect 152220 684210 152310 684450
rect 152550 684210 152640 684450
rect 152880 684210 152990 684450
rect 153230 684210 153320 684450
rect 153560 684210 153650 684450
rect 153890 684210 153980 684450
rect 154220 684210 154330 684450
rect 154570 684210 154660 684450
rect 154900 684210 154990 684450
rect 155230 684210 155320 684450
rect 155560 684210 155670 684450
rect 155910 684210 155930 684450
rect 144930 684120 155930 684210
rect 144930 683880 144950 684120
rect 145190 683880 145280 684120
rect 145520 683880 145610 684120
rect 145850 683880 145940 684120
rect 146180 683880 146290 684120
rect 146530 683880 146620 684120
rect 146860 683880 146950 684120
rect 147190 683880 147280 684120
rect 147520 683880 147630 684120
rect 147870 683880 147960 684120
rect 148200 683880 148290 684120
rect 148530 683880 148620 684120
rect 148860 683880 148970 684120
rect 149210 683880 149300 684120
rect 149540 683880 149630 684120
rect 149870 683880 149960 684120
rect 150200 683880 150310 684120
rect 150550 683880 150640 684120
rect 150880 683880 150970 684120
rect 151210 683880 151300 684120
rect 151540 683880 151650 684120
rect 151890 683880 151980 684120
rect 152220 683880 152310 684120
rect 152550 683880 152640 684120
rect 152880 683880 152990 684120
rect 153230 683880 153320 684120
rect 153560 683880 153650 684120
rect 153890 683880 153980 684120
rect 154220 683880 154330 684120
rect 154570 683880 154660 684120
rect 154900 683880 154990 684120
rect 155230 683880 155320 684120
rect 155560 683880 155670 684120
rect 155910 683880 155930 684120
rect 144930 683860 155930 683880
rect 110790 683280 121790 683300
rect 110790 683040 110810 683280
rect 111050 683040 111160 683280
rect 111400 683040 111490 683280
rect 111730 683040 111820 683280
rect 112060 683040 112150 683280
rect 112390 683040 112500 683280
rect 112740 683040 112830 683280
rect 113070 683040 113160 683280
rect 113400 683040 113490 683280
rect 113730 683040 113840 683280
rect 114080 683040 114170 683280
rect 114410 683040 114500 683280
rect 114740 683040 114830 683280
rect 115070 683040 115180 683280
rect 115420 683040 115510 683280
rect 115750 683040 115840 683280
rect 116080 683040 116170 683280
rect 116410 683040 116520 683280
rect 116760 683040 116850 683280
rect 117090 683040 117180 683280
rect 117420 683040 117510 683280
rect 117750 683040 117860 683280
rect 118100 683040 118190 683280
rect 118430 683040 118520 683280
rect 118760 683040 118850 683280
rect 119090 683040 119200 683280
rect 119440 683040 119530 683280
rect 119770 683040 119860 683280
rect 120100 683040 120190 683280
rect 120430 683040 120540 683280
rect 120780 683040 120870 683280
rect 121110 683040 121200 683280
rect 121440 683040 121530 683280
rect 121770 683040 121790 683280
rect 110790 682950 121790 683040
rect 110790 682710 110810 682950
rect 111050 682710 111160 682950
rect 111400 682710 111490 682950
rect 111730 682710 111820 682950
rect 112060 682710 112150 682950
rect 112390 682710 112500 682950
rect 112740 682710 112830 682950
rect 113070 682710 113160 682950
rect 113400 682710 113490 682950
rect 113730 682710 113840 682950
rect 114080 682710 114170 682950
rect 114410 682710 114500 682950
rect 114740 682710 114830 682950
rect 115070 682710 115180 682950
rect 115420 682710 115510 682950
rect 115750 682710 115840 682950
rect 116080 682710 116170 682950
rect 116410 682710 116520 682950
rect 116760 682710 116850 682950
rect 117090 682710 117180 682950
rect 117420 682710 117510 682950
rect 117750 682710 117860 682950
rect 118100 682710 118190 682950
rect 118430 682710 118520 682950
rect 118760 682710 118850 682950
rect 119090 682710 119200 682950
rect 119440 682710 119530 682950
rect 119770 682710 119860 682950
rect 120100 682710 120190 682950
rect 120430 682710 120540 682950
rect 120780 682710 120870 682950
rect 121110 682710 121200 682950
rect 121440 682710 121530 682950
rect 121770 682710 121790 682950
rect 110790 682620 121790 682710
rect 110790 682380 110810 682620
rect 111050 682380 111160 682620
rect 111400 682380 111490 682620
rect 111730 682380 111820 682620
rect 112060 682380 112150 682620
rect 112390 682380 112500 682620
rect 112740 682380 112830 682620
rect 113070 682380 113160 682620
rect 113400 682380 113490 682620
rect 113730 682380 113840 682620
rect 114080 682380 114170 682620
rect 114410 682380 114500 682620
rect 114740 682380 114830 682620
rect 115070 682380 115180 682620
rect 115420 682380 115510 682620
rect 115750 682380 115840 682620
rect 116080 682380 116170 682620
rect 116410 682380 116520 682620
rect 116760 682380 116850 682620
rect 117090 682380 117180 682620
rect 117420 682380 117510 682620
rect 117750 682380 117860 682620
rect 118100 682380 118190 682620
rect 118430 682380 118520 682620
rect 118760 682380 118850 682620
rect 119090 682380 119200 682620
rect 119440 682380 119530 682620
rect 119770 682380 119860 682620
rect 120100 682380 120190 682620
rect 120430 682380 120540 682620
rect 120780 682380 120870 682620
rect 121110 682380 121200 682620
rect 121440 682380 121530 682620
rect 121770 682380 121790 682620
rect 110790 682290 121790 682380
rect 110790 682050 110810 682290
rect 111050 682050 111160 682290
rect 111400 682050 111490 682290
rect 111730 682050 111820 682290
rect 112060 682050 112150 682290
rect 112390 682050 112500 682290
rect 112740 682050 112830 682290
rect 113070 682050 113160 682290
rect 113400 682050 113490 682290
rect 113730 682050 113840 682290
rect 114080 682050 114170 682290
rect 114410 682050 114500 682290
rect 114740 682050 114830 682290
rect 115070 682050 115180 682290
rect 115420 682050 115510 682290
rect 115750 682050 115840 682290
rect 116080 682050 116170 682290
rect 116410 682050 116520 682290
rect 116760 682050 116850 682290
rect 117090 682050 117180 682290
rect 117420 682050 117510 682290
rect 117750 682050 117860 682290
rect 118100 682050 118190 682290
rect 118430 682050 118520 682290
rect 118760 682050 118850 682290
rect 119090 682050 119200 682290
rect 119440 682050 119530 682290
rect 119770 682050 119860 682290
rect 120100 682050 120190 682290
rect 120430 682050 120540 682290
rect 120780 682050 120870 682290
rect 121110 682050 121200 682290
rect 121440 682050 121530 682290
rect 121770 682050 121790 682290
rect 110790 681940 121790 682050
rect 110790 681700 110810 681940
rect 111050 681700 111160 681940
rect 111400 681700 111490 681940
rect 111730 681700 111820 681940
rect 112060 681700 112150 681940
rect 112390 681700 112500 681940
rect 112740 681700 112830 681940
rect 113070 681700 113160 681940
rect 113400 681700 113490 681940
rect 113730 681700 113840 681940
rect 114080 681700 114170 681940
rect 114410 681700 114500 681940
rect 114740 681700 114830 681940
rect 115070 681700 115180 681940
rect 115420 681700 115510 681940
rect 115750 681700 115840 681940
rect 116080 681700 116170 681940
rect 116410 681700 116520 681940
rect 116760 681700 116850 681940
rect 117090 681700 117180 681940
rect 117420 681700 117510 681940
rect 117750 681700 117860 681940
rect 118100 681700 118190 681940
rect 118430 681700 118520 681940
rect 118760 681700 118850 681940
rect 119090 681700 119200 681940
rect 119440 681700 119530 681940
rect 119770 681700 119860 681940
rect 120100 681700 120190 681940
rect 120430 681700 120540 681940
rect 120780 681700 120870 681940
rect 121110 681700 121200 681940
rect 121440 681700 121530 681940
rect 121770 681700 121790 681940
rect 110790 681610 121790 681700
rect 110790 681370 110810 681610
rect 111050 681370 111160 681610
rect 111400 681370 111490 681610
rect 111730 681370 111820 681610
rect 112060 681370 112150 681610
rect 112390 681370 112500 681610
rect 112740 681370 112830 681610
rect 113070 681370 113160 681610
rect 113400 681370 113490 681610
rect 113730 681370 113840 681610
rect 114080 681370 114170 681610
rect 114410 681370 114500 681610
rect 114740 681370 114830 681610
rect 115070 681370 115180 681610
rect 115420 681370 115510 681610
rect 115750 681370 115840 681610
rect 116080 681370 116170 681610
rect 116410 681370 116520 681610
rect 116760 681370 116850 681610
rect 117090 681370 117180 681610
rect 117420 681370 117510 681610
rect 117750 681370 117860 681610
rect 118100 681370 118190 681610
rect 118430 681370 118520 681610
rect 118760 681370 118850 681610
rect 119090 681370 119200 681610
rect 119440 681370 119530 681610
rect 119770 681370 119860 681610
rect 120100 681370 120190 681610
rect 120430 681370 120540 681610
rect 120780 681370 120870 681610
rect 121110 681370 121200 681610
rect 121440 681370 121530 681610
rect 121770 681370 121790 681610
rect 110790 681280 121790 681370
rect 110790 681040 110810 681280
rect 111050 681040 111160 681280
rect 111400 681040 111490 681280
rect 111730 681040 111820 681280
rect 112060 681040 112150 681280
rect 112390 681040 112500 681280
rect 112740 681040 112830 681280
rect 113070 681040 113160 681280
rect 113400 681040 113490 681280
rect 113730 681040 113840 681280
rect 114080 681040 114170 681280
rect 114410 681040 114500 681280
rect 114740 681040 114830 681280
rect 115070 681040 115180 681280
rect 115420 681040 115510 681280
rect 115750 681040 115840 681280
rect 116080 681040 116170 681280
rect 116410 681040 116520 681280
rect 116760 681040 116850 681280
rect 117090 681040 117180 681280
rect 117420 681040 117510 681280
rect 117750 681040 117860 681280
rect 118100 681040 118190 681280
rect 118430 681040 118520 681280
rect 118760 681040 118850 681280
rect 119090 681040 119200 681280
rect 119440 681040 119530 681280
rect 119770 681040 119860 681280
rect 120100 681040 120190 681280
rect 120430 681040 120540 681280
rect 120780 681040 120870 681280
rect 121110 681040 121200 681280
rect 121440 681040 121530 681280
rect 121770 681040 121790 681280
rect 110790 680950 121790 681040
rect 110790 680710 110810 680950
rect 111050 680710 111160 680950
rect 111400 680710 111490 680950
rect 111730 680710 111820 680950
rect 112060 680710 112150 680950
rect 112390 680710 112500 680950
rect 112740 680710 112830 680950
rect 113070 680710 113160 680950
rect 113400 680710 113490 680950
rect 113730 680710 113840 680950
rect 114080 680710 114170 680950
rect 114410 680710 114500 680950
rect 114740 680710 114830 680950
rect 115070 680710 115180 680950
rect 115420 680710 115510 680950
rect 115750 680710 115840 680950
rect 116080 680710 116170 680950
rect 116410 680710 116520 680950
rect 116760 680710 116850 680950
rect 117090 680710 117180 680950
rect 117420 680710 117510 680950
rect 117750 680710 117860 680950
rect 118100 680710 118190 680950
rect 118430 680710 118520 680950
rect 118760 680710 118850 680950
rect 119090 680710 119200 680950
rect 119440 680710 119530 680950
rect 119770 680710 119860 680950
rect 120100 680710 120190 680950
rect 120430 680710 120540 680950
rect 120780 680710 120870 680950
rect 121110 680710 121200 680950
rect 121440 680710 121530 680950
rect 121770 680710 121790 680950
rect 110790 680600 121790 680710
rect 110790 680360 110810 680600
rect 111050 680360 111160 680600
rect 111400 680360 111490 680600
rect 111730 680360 111820 680600
rect 112060 680360 112150 680600
rect 112390 680360 112500 680600
rect 112740 680360 112830 680600
rect 113070 680360 113160 680600
rect 113400 680360 113490 680600
rect 113730 680360 113840 680600
rect 114080 680360 114170 680600
rect 114410 680360 114500 680600
rect 114740 680360 114830 680600
rect 115070 680360 115180 680600
rect 115420 680360 115510 680600
rect 115750 680360 115840 680600
rect 116080 680360 116170 680600
rect 116410 680360 116520 680600
rect 116760 680360 116850 680600
rect 117090 680360 117180 680600
rect 117420 680360 117510 680600
rect 117750 680360 117860 680600
rect 118100 680360 118190 680600
rect 118430 680360 118520 680600
rect 118760 680360 118850 680600
rect 119090 680360 119200 680600
rect 119440 680360 119530 680600
rect 119770 680360 119860 680600
rect 120100 680360 120190 680600
rect 120430 680360 120540 680600
rect 120780 680360 120870 680600
rect 121110 680360 121200 680600
rect 121440 680360 121530 680600
rect 121770 680360 121790 680600
rect 110790 680270 121790 680360
rect 110790 680030 110810 680270
rect 111050 680030 111160 680270
rect 111400 680030 111490 680270
rect 111730 680030 111820 680270
rect 112060 680030 112150 680270
rect 112390 680030 112500 680270
rect 112740 680030 112830 680270
rect 113070 680030 113160 680270
rect 113400 680030 113490 680270
rect 113730 680030 113840 680270
rect 114080 680030 114170 680270
rect 114410 680030 114500 680270
rect 114740 680030 114830 680270
rect 115070 680030 115180 680270
rect 115420 680030 115510 680270
rect 115750 680030 115840 680270
rect 116080 680030 116170 680270
rect 116410 680030 116520 680270
rect 116760 680030 116850 680270
rect 117090 680030 117180 680270
rect 117420 680030 117510 680270
rect 117750 680030 117860 680270
rect 118100 680030 118190 680270
rect 118430 680030 118520 680270
rect 118760 680030 118850 680270
rect 119090 680030 119200 680270
rect 119440 680030 119530 680270
rect 119770 680030 119860 680270
rect 120100 680030 120190 680270
rect 120430 680030 120540 680270
rect 120780 680030 120870 680270
rect 121110 680030 121200 680270
rect 121440 680030 121530 680270
rect 121770 680030 121790 680270
rect 110790 679940 121790 680030
rect 110790 679700 110810 679940
rect 111050 679700 111160 679940
rect 111400 679700 111490 679940
rect 111730 679700 111820 679940
rect 112060 679700 112150 679940
rect 112390 679700 112500 679940
rect 112740 679700 112830 679940
rect 113070 679700 113160 679940
rect 113400 679700 113490 679940
rect 113730 679700 113840 679940
rect 114080 679700 114170 679940
rect 114410 679700 114500 679940
rect 114740 679700 114830 679940
rect 115070 679700 115180 679940
rect 115420 679700 115510 679940
rect 115750 679700 115840 679940
rect 116080 679700 116170 679940
rect 116410 679700 116520 679940
rect 116760 679700 116850 679940
rect 117090 679700 117180 679940
rect 117420 679700 117510 679940
rect 117750 679700 117860 679940
rect 118100 679700 118190 679940
rect 118430 679700 118520 679940
rect 118760 679700 118850 679940
rect 119090 679700 119200 679940
rect 119440 679700 119530 679940
rect 119770 679700 119860 679940
rect 120100 679700 120190 679940
rect 120430 679700 120540 679940
rect 120780 679700 120870 679940
rect 121110 679700 121200 679940
rect 121440 679700 121530 679940
rect 121770 679700 121790 679940
rect 110790 679610 121790 679700
rect 110790 679370 110810 679610
rect 111050 679370 111160 679610
rect 111400 679370 111490 679610
rect 111730 679370 111820 679610
rect 112060 679370 112150 679610
rect 112390 679370 112500 679610
rect 112740 679370 112830 679610
rect 113070 679370 113160 679610
rect 113400 679370 113490 679610
rect 113730 679370 113840 679610
rect 114080 679370 114170 679610
rect 114410 679370 114500 679610
rect 114740 679370 114830 679610
rect 115070 679370 115180 679610
rect 115420 679370 115510 679610
rect 115750 679370 115840 679610
rect 116080 679370 116170 679610
rect 116410 679370 116520 679610
rect 116760 679370 116850 679610
rect 117090 679370 117180 679610
rect 117420 679370 117510 679610
rect 117750 679370 117860 679610
rect 118100 679370 118190 679610
rect 118430 679370 118520 679610
rect 118760 679370 118850 679610
rect 119090 679370 119200 679610
rect 119440 679370 119530 679610
rect 119770 679370 119860 679610
rect 120100 679370 120190 679610
rect 120430 679370 120540 679610
rect 120780 679370 120870 679610
rect 121110 679370 121200 679610
rect 121440 679370 121530 679610
rect 121770 679370 121790 679610
rect 110790 679260 121790 679370
rect 110790 679020 110810 679260
rect 111050 679020 111160 679260
rect 111400 679020 111490 679260
rect 111730 679020 111820 679260
rect 112060 679020 112150 679260
rect 112390 679020 112500 679260
rect 112740 679020 112830 679260
rect 113070 679020 113160 679260
rect 113400 679020 113490 679260
rect 113730 679020 113840 679260
rect 114080 679020 114170 679260
rect 114410 679020 114500 679260
rect 114740 679020 114830 679260
rect 115070 679020 115180 679260
rect 115420 679020 115510 679260
rect 115750 679020 115840 679260
rect 116080 679020 116170 679260
rect 116410 679020 116520 679260
rect 116760 679020 116850 679260
rect 117090 679020 117180 679260
rect 117420 679020 117510 679260
rect 117750 679020 117860 679260
rect 118100 679020 118190 679260
rect 118430 679020 118520 679260
rect 118760 679020 118850 679260
rect 119090 679020 119200 679260
rect 119440 679020 119530 679260
rect 119770 679020 119860 679260
rect 120100 679020 120190 679260
rect 120430 679020 120540 679260
rect 120780 679020 120870 679260
rect 121110 679020 121200 679260
rect 121440 679020 121530 679260
rect 121770 679020 121790 679260
rect 110790 678930 121790 679020
rect 110790 678690 110810 678930
rect 111050 678690 111160 678930
rect 111400 678690 111490 678930
rect 111730 678690 111820 678930
rect 112060 678690 112150 678930
rect 112390 678690 112500 678930
rect 112740 678690 112830 678930
rect 113070 678690 113160 678930
rect 113400 678690 113490 678930
rect 113730 678690 113840 678930
rect 114080 678690 114170 678930
rect 114410 678690 114500 678930
rect 114740 678690 114830 678930
rect 115070 678690 115180 678930
rect 115420 678690 115510 678930
rect 115750 678690 115840 678930
rect 116080 678690 116170 678930
rect 116410 678690 116520 678930
rect 116760 678690 116850 678930
rect 117090 678690 117180 678930
rect 117420 678690 117510 678930
rect 117750 678690 117860 678930
rect 118100 678690 118190 678930
rect 118430 678690 118520 678930
rect 118760 678690 118850 678930
rect 119090 678690 119200 678930
rect 119440 678690 119530 678930
rect 119770 678690 119860 678930
rect 120100 678690 120190 678930
rect 120430 678690 120540 678930
rect 120780 678690 120870 678930
rect 121110 678690 121200 678930
rect 121440 678690 121530 678930
rect 121770 678690 121790 678930
rect 110790 678600 121790 678690
rect 110790 678360 110810 678600
rect 111050 678360 111160 678600
rect 111400 678360 111490 678600
rect 111730 678360 111820 678600
rect 112060 678360 112150 678600
rect 112390 678360 112500 678600
rect 112740 678360 112830 678600
rect 113070 678360 113160 678600
rect 113400 678360 113490 678600
rect 113730 678360 113840 678600
rect 114080 678360 114170 678600
rect 114410 678360 114500 678600
rect 114740 678360 114830 678600
rect 115070 678360 115180 678600
rect 115420 678360 115510 678600
rect 115750 678360 115840 678600
rect 116080 678360 116170 678600
rect 116410 678360 116520 678600
rect 116760 678360 116850 678600
rect 117090 678360 117180 678600
rect 117420 678360 117510 678600
rect 117750 678360 117860 678600
rect 118100 678360 118190 678600
rect 118430 678360 118520 678600
rect 118760 678360 118850 678600
rect 119090 678360 119200 678600
rect 119440 678360 119530 678600
rect 119770 678360 119860 678600
rect 120100 678360 120190 678600
rect 120430 678360 120540 678600
rect 120780 678360 120870 678600
rect 121110 678360 121200 678600
rect 121440 678360 121530 678600
rect 121770 678360 121790 678600
rect 110790 678270 121790 678360
rect 110790 678030 110810 678270
rect 111050 678030 111160 678270
rect 111400 678030 111490 678270
rect 111730 678030 111820 678270
rect 112060 678030 112150 678270
rect 112390 678030 112500 678270
rect 112740 678030 112830 678270
rect 113070 678030 113160 678270
rect 113400 678030 113490 678270
rect 113730 678030 113840 678270
rect 114080 678030 114170 678270
rect 114410 678030 114500 678270
rect 114740 678030 114830 678270
rect 115070 678030 115180 678270
rect 115420 678030 115510 678270
rect 115750 678030 115840 678270
rect 116080 678030 116170 678270
rect 116410 678030 116520 678270
rect 116760 678030 116850 678270
rect 117090 678030 117180 678270
rect 117420 678030 117510 678270
rect 117750 678030 117860 678270
rect 118100 678030 118190 678270
rect 118430 678030 118520 678270
rect 118760 678030 118850 678270
rect 119090 678030 119200 678270
rect 119440 678030 119530 678270
rect 119770 678030 119860 678270
rect 120100 678030 120190 678270
rect 120430 678030 120540 678270
rect 120780 678030 120870 678270
rect 121110 678030 121200 678270
rect 121440 678030 121530 678270
rect 121770 678030 121790 678270
rect 110790 677920 121790 678030
rect 110790 677680 110810 677920
rect 111050 677680 111160 677920
rect 111400 677680 111490 677920
rect 111730 677680 111820 677920
rect 112060 677680 112150 677920
rect 112390 677680 112500 677920
rect 112740 677680 112830 677920
rect 113070 677680 113160 677920
rect 113400 677680 113490 677920
rect 113730 677680 113840 677920
rect 114080 677680 114170 677920
rect 114410 677680 114500 677920
rect 114740 677680 114830 677920
rect 115070 677680 115180 677920
rect 115420 677680 115510 677920
rect 115750 677680 115840 677920
rect 116080 677680 116170 677920
rect 116410 677680 116520 677920
rect 116760 677680 116850 677920
rect 117090 677680 117180 677920
rect 117420 677680 117510 677920
rect 117750 677680 117860 677920
rect 118100 677680 118190 677920
rect 118430 677680 118520 677920
rect 118760 677680 118850 677920
rect 119090 677680 119200 677920
rect 119440 677680 119530 677920
rect 119770 677680 119860 677920
rect 120100 677680 120190 677920
rect 120430 677680 120540 677920
rect 120780 677680 120870 677920
rect 121110 677680 121200 677920
rect 121440 677680 121530 677920
rect 121770 677680 121790 677920
rect 110790 677590 121790 677680
rect 110790 677350 110810 677590
rect 111050 677350 111160 677590
rect 111400 677350 111490 677590
rect 111730 677350 111820 677590
rect 112060 677350 112150 677590
rect 112390 677350 112500 677590
rect 112740 677350 112830 677590
rect 113070 677350 113160 677590
rect 113400 677350 113490 677590
rect 113730 677350 113840 677590
rect 114080 677350 114170 677590
rect 114410 677350 114500 677590
rect 114740 677350 114830 677590
rect 115070 677350 115180 677590
rect 115420 677350 115510 677590
rect 115750 677350 115840 677590
rect 116080 677350 116170 677590
rect 116410 677350 116520 677590
rect 116760 677350 116850 677590
rect 117090 677350 117180 677590
rect 117420 677350 117510 677590
rect 117750 677350 117860 677590
rect 118100 677350 118190 677590
rect 118430 677350 118520 677590
rect 118760 677350 118850 677590
rect 119090 677350 119200 677590
rect 119440 677350 119530 677590
rect 119770 677350 119860 677590
rect 120100 677350 120190 677590
rect 120430 677350 120540 677590
rect 120780 677350 120870 677590
rect 121110 677350 121200 677590
rect 121440 677350 121530 677590
rect 121770 677350 121790 677590
rect 110790 677260 121790 677350
rect 110790 677020 110810 677260
rect 111050 677020 111160 677260
rect 111400 677020 111490 677260
rect 111730 677020 111820 677260
rect 112060 677020 112150 677260
rect 112390 677020 112500 677260
rect 112740 677020 112830 677260
rect 113070 677020 113160 677260
rect 113400 677020 113490 677260
rect 113730 677020 113840 677260
rect 114080 677020 114170 677260
rect 114410 677020 114500 677260
rect 114740 677020 114830 677260
rect 115070 677020 115180 677260
rect 115420 677020 115510 677260
rect 115750 677020 115840 677260
rect 116080 677020 116170 677260
rect 116410 677020 116520 677260
rect 116760 677020 116850 677260
rect 117090 677020 117180 677260
rect 117420 677020 117510 677260
rect 117750 677020 117860 677260
rect 118100 677020 118190 677260
rect 118430 677020 118520 677260
rect 118760 677020 118850 677260
rect 119090 677020 119200 677260
rect 119440 677020 119530 677260
rect 119770 677020 119860 677260
rect 120100 677020 120190 677260
rect 120430 677020 120540 677260
rect 120780 677020 120870 677260
rect 121110 677020 121200 677260
rect 121440 677020 121530 677260
rect 121770 677020 121790 677260
rect 110790 676930 121790 677020
rect 110790 676690 110810 676930
rect 111050 676690 111160 676930
rect 111400 676690 111490 676930
rect 111730 676690 111820 676930
rect 112060 676690 112150 676930
rect 112390 676690 112500 676930
rect 112740 676690 112830 676930
rect 113070 676690 113160 676930
rect 113400 676690 113490 676930
rect 113730 676690 113840 676930
rect 114080 676690 114170 676930
rect 114410 676690 114500 676930
rect 114740 676690 114830 676930
rect 115070 676690 115180 676930
rect 115420 676690 115510 676930
rect 115750 676690 115840 676930
rect 116080 676690 116170 676930
rect 116410 676690 116520 676930
rect 116760 676690 116850 676930
rect 117090 676690 117180 676930
rect 117420 676690 117510 676930
rect 117750 676690 117860 676930
rect 118100 676690 118190 676930
rect 118430 676690 118520 676930
rect 118760 676690 118850 676930
rect 119090 676690 119200 676930
rect 119440 676690 119530 676930
rect 119770 676690 119860 676930
rect 120100 676690 120190 676930
rect 120430 676690 120540 676930
rect 120780 676690 120870 676930
rect 121110 676690 121200 676930
rect 121440 676690 121530 676930
rect 121770 676690 121790 676930
rect 110790 676580 121790 676690
rect 110790 676340 110810 676580
rect 111050 676340 111160 676580
rect 111400 676340 111490 676580
rect 111730 676340 111820 676580
rect 112060 676340 112150 676580
rect 112390 676340 112500 676580
rect 112740 676340 112830 676580
rect 113070 676340 113160 676580
rect 113400 676340 113490 676580
rect 113730 676340 113840 676580
rect 114080 676340 114170 676580
rect 114410 676340 114500 676580
rect 114740 676340 114830 676580
rect 115070 676340 115180 676580
rect 115420 676340 115510 676580
rect 115750 676340 115840 676580
rect 116080 676340 116170 676580
rect 116410 676340 116520 676580
rect 116760 676340 116850 676580
rect 117090 676340 117180 676580
rect 117420 676340 117510 676580
rect 117750 676340 117860 676580
rect 118100 676340 118190 676580
rect 118430 676340 118520 676580
rect 118760 676340 118850 676580
rect 119090 676340 119200 676580
rect 119440 676340 119530 676580
rect 119770 676340 119860 676580
rect 120100 676340 120190 676580
rect 120430 676340 120540 676580
rect 120780 676340 120870 676580
rect 121110 676340 121200 676580
rect 121440 676340 121530 676580
rect 121770 676340 121790 676580
rect 110790 676250 121790 676340
rect 110790 676010 110810 676250
rect 111050 676010 111160 676250
rect 111400 676010 111490 676250
rect 111730 676010 111820 676250
rect 112060 676010 112150 676250
rect 112390 676010 112500 676250
rect 112740 676010 112830 676250
rect 113070 676010 113160 676250
rect 113400 676010 113490 676250
rect 113730 676010 113840 676250
rect 114080 676010 114170 676250
rect 114410 676010 114500 676250
rect 114740 676010 114830 676250
rect 115070 676010 115180 676250
rect 115420 676010 115510 676250
rect 115750 676010 115840 676250
rect 116080 676010 116170 676250
rect 116410 676010 116520 676250
rect 116760 676010 116850 676250
rect 117090 676010 117180 676250
rect 117420 676010 117510 676250
rect 117750 676010 117860 676250
rect 118100 676010 118190 676250
rect 118430 676010 118520 676250
rect 118760 676010 118850 676250
rect 119090 676010 119200 676250
rect 119440 676010 119530 676250
rect 119770 676010 119860 676250
rect 120100 676010 120190 676250
rect 120430 676010 120540 676250
rect 120780 676010 120870 676250
rect 121110 676010 121200 676250
rect 121440 676010 121530 676250
rect 121770 676010 121790 676250
rect 110790 675920 121790 676010
rect 110790 675680 110810 675920
rect 111050 675680 111160 675920
rect 111400 675680 111490 675920
rect 111730 675680 111820 675920
rect 112060 675680 112150 675920
rect 112390 675680 112500 675920
rect 112740 675680 112830 675920
rect 113070 675680 113160 675920
rect 113400 675680 113490 675920
rect 113730 675680 113840 675920
rect 114080 675680 114170 675920
rect 114410 675680 114500 675920
rect 114740 675680 114830 675920
rect 115070 675680 115180 675920
rect 115420 675680 115510 675920
rect 115750 675680 115840 675920
rect 116080 675680 116170 675920
rect 116410 675680 116520 675920
rect 116760 675680 116850 675920
rect 117090 675680 117180 675920
rect 117420 675680 117510 675920
rect 117750 675680 117860 675920
rect 118100 675680 118190 675920
rect 118430 675680 118520 675920
rect 118760 675680 118850 675920
rect 119090 675680 119200 675920
rect 119440 675680 119530 675920
rect 119770 675680 119860 675920
rect 120100 675680 120190 675920
rect 120430 675680 120540 675920
rect 120780 675680 120870 675920
rect 121110 675680 121200 675920
rect 121440 675680 121530 675920
rect 121770 675680 121790 675920
rect 110790 675590 121790 675680
rect 110790 675350 110810 675590
rect 111050 675350 111160 675590
rect 111400 675350 111490 675590
rect 111730 675350 111820 675590
rect 112060 675350 112150 675590
rect 112390 675350 112500 675590
rect 112740 675350 112830 675590
rect 113070 675350 113160 675590
rect 113400 675350 113490 675590
rect 113730 675350 113840 675590
rect 114080 675350 114170 675590
rect 114410 675350 114500 675590
rect 114740 675350 114830 675590
rect 115070 675350 115180 675590
rect 115420 675350 115510 675590
rect 115750 675350 115840 675590
rect 116080 675350 116170 675590
rect 116410 675350 116520 675590
rect 116760 675350 116850 675590
rect 117090 675350 117180 675590
rect 117420 675350 117510 675590
rect 117750 675350 117860 675590
rect 118100 675350 118190 675590
rect 118430 675350 118520 675590
rect 118760 675350 118850 675590
rect 119090 675350 119200 675590
rect 119440 675350 119530 675590
rect 119770 675350 119860 675590
rect 120100 675350 120190 675590
rect 120430 675350 120540 675590
rect 120780 675350 120870 675590
rect 121110 675350 121200 675590
rect 121440 675350 121530 675590
rect 121770 675350 121790 675590
rect 110790 675240 121790 675350
rect 110790 675000 110810 675240
rect 111050 675000 111160 675240
rect 111400 675000 111490 675240
rect 111730 675000 111820 675240
rect 112060 675000 112150 675240
rect 112390 675000 112500 675240
rect 112740 675000 112830 675240
rect 113070 675000 113160 675240
rect 113400 675000 113490 675240
rect 113730 675000 113840 675240
rect 114080 675000 114170 675240
rect 114410 675000 114500 675240
rect 114740 675000 114830 675240
rect 115070 675000 115180 675240
rect 115420 675000 115510 675240
rect 115750 675000 115840 675240
rect 116080 675000 116170 675240
rect 116410 675000 116520 675240
rect 116760 675000 116850 675240
rect 117090 675000 117180 675240
rect 117420 675000 117510 675240
rect 117750 675000 117860 675240
rect 118100 675000 118190 675240
rect 118430 675000 118520 675240
rect 118760 675000 118850 675240
rect 119090 675000 119200 675240
rect 119440 675000 119530 675240
rect 119770 675000 119860 675240
rect 120100 675000 120190 675240
rect 120430 675000 120540 675240
rect 120780 675000 120870 675240
rect 121110 675000 121200 675240
rect 121440 675000 121530 675240
rect 121770 675000 121790 675240
rect 110790 674910 121790 675000
rect 110790 674670 110810 674910
rect 111050 674670 111160 674910
rect 111400 674670 111490 674910
rect 111730 674670 111820 674910
rect 112060 674670 112150 674910
rect 112390 674670 112500 674910
rect 112740 674670 112830 674910
rect 113070 674670 113160 674910
rect 113400 674670 113490 674910
rect 113730 674670 113840 674910
rect 114080 674670 114170 674910
rect 114410 674670 114500 674910
rect 114740 674670 114830 674910
rect 115070 674670 115180 674910
rect 115420 674670 115510 674910
rect 115750 674670 115840 674910
rect 116080 674670 116170 674910
rect 116410 674670 116520 674910
rect 116760 674670 116850 674910
rect 117090 674670 117180 674910
rect 117420 674670 117510 674910
rect 117750 674670 117860 674910
rect 118100 674670 118190 674910
rect 118430 674670 118520 674910
rect 118760 674670 118850 674910
rect 119090 674670 119200 674910
rect 119440 674670 119530 674910
rect 119770 674670 119860 674910
rect 120100 674670 120190 674910
rect 120430 674670 120540 674910
rect 120780 674670 120870 674910
rect 121110 674670 121200 674910
rect 121440 674670 121530 674910
rect 121770 674670 121790 674910
rect 110790 674580 121790 674670
rect 110790 674340 110810 674580
rect 111050 674340 111160 674580
rect 111400 674340 111490 674580
rect 111730 674340 111820 674580
rect 112060 674340 112150 674580
rect 112390 674340 112500 674580
rect 112740 674340 112830 674580
rect 113070 674340 113160 674580
rect 113400 674340 113490 674580
rect 113730 674340 113840 674580
rect 114080 674340 114170 674580
rect 114410 674340 114500 674580
rect 114740 674340 114830 674580
rect 115070 674340 115180 674580
rect 115420 674340 115510 674580
rect 115750 674340 115840 674580
rect 116080 674340 116170 674580
rect 116410 674340 116520 674580
rect 116760 674340 116850 674580
rect 117090 674340 117180 674580
rect 117420 674340 117510 674580
rect 117750 674340 117860 674580
rect 118100 674340 118190 674580
rect 118430 674340 118520 674580
rect 118760 674340 118850 674580
rect 119090 674340 119200 674580
rect 119440 674340 119530 674580
rect 119770 674340 119860 674580
rect 120100 674340 120190 674580
rect 120430 674340 120540 674580
rect 120780 674340 120870 674580
rect 121110 674340 121200 674580
rect 121440 674340 121530 674580
rect 121770 674340 121790 674580
rect 110790 674250 121790 674340
rect 110790 674010 110810 674250
rect 111050 674010 111160 674250
rect 111400 674010 111490 674250
rect 111730 674010 111820 674250
rect 112060 674010 112150 674250
rect 112390 674010 112500 674250
rect 112740 674010 112830 674250
rect 113070 674010 113160 674250
rect 113400 674010 113490 674250
rect 113730 674010 113840 674250
rect 114080 674010 114170 674250
rect 114410 674010 114500 674250
rect 114740 674010 114830 674250
rect 115070 674010 115180 674250
rect 115420 674010 115510 674250
rect 115750 674010 115840 674250
rect 116080 674010 116170 674250
rect 116410 674010 116520 674250
rect 116760 674010 116850 674250
rect 117090 674010 117180 674250
rect 117420 674010 117510 674250
rect 117750 674010 117860 674250
rect 118100 674010 118190 674250
rect 118430 674010 118520 674250
rect 118760 674010 118850 674250
rect 119090 674010 119200 674250
rect 119440 674010 119530 674250
rect 119770 674010 119860 674250
rect 120100 674010 120190 674250
rect 120430 674010 120540 674250
rect 120780 674010 120870 674250
rect 121110 674010 121200 674250
rect 121440 674010 121530 674250
rect 121770 674010 121790 674250
rect 110790 673900 121790 674010
rect 110790 673660 110810 673900
rect 111050 673660 111160 673900
rect 111400 673660 111490 673900
rect 111730 673660 111820 673900
rect 112060 673660 112150 673900
rect 112390 673660 112500 673900
rect 112740 673660 112830 673900
rect 113070 673660 113160 673900
rect 113400 673660 113490 673900
rect 113730 673660 113840 673900
rect 114080 673660 114170 673900
rect 114410 673660 114500 673900
rect 114740 673660 114830 673900
rect 115070 673660 115180 673900
rect 115420 673660 115510 673900
rect 115750 673660 115840 673900
rect 116080 673660 116170 673900
rect 116410 673660 116520 673900
rect 116760 673660 116850 673900
rect 117090 673660 117180 673900
rect 117420 673660 117510 673900
rect 117750 673660 117860 673900
rect 118100 673660 118190 673900
rect 118430 673660 118520 673900
rect 118760 673660 118850 673900
rect 119090 673660 119200 673900
rect 119440 673660 119530 673900
rect 119770 673660 119860 673900
rect 120100 673660 120190 673900
rect 120430 673660 120540 673900
rect 120780 673660 120870 673900
rect 121110 673660 121200 673900
rect 121440 673660 121530 673900
rect 121770 673660 121790 673900
rect 110790 673570 121790 673660
rect 110790 673330 110810 673570
rect 111050 673330 111160 673570
rect 111400 673330 111490 673570
rect 111730 673330 111820 673570
rect 112060 673330 112150 673570
rect 112390 673330 112500 673570
rect 112740 673330 112830 673570
rect 113070 673330 113160 673570
rect 113400 673330 113490 673570
rect 113730 673330 113840 673570
rect 114080 673330 114170 673570
rect 114410 673330 114500 673570
rect 114740 673330 114830 673570
rect 115070 673330 115180 673570
rect 115420 673330 115510 673570
rect 115750 673330 115840 673570
rect 116080 673330 116170 673570
rect 116410 673330 116520 673570
rect 116760 673330 116850 673570
rect 117090 673330 117180 673570
rect 117420 673330 117510 673570
rect 117750 673330 117860 673570
rect 118100 673330 118190 673570
rect 118430 673330 118520 673570
rect 118760 673330 118850 673570
rect 119090 673330 119200 673570
rect 119440 673330 119530 673570
rect 119770 673330 119860 673570
rect 120100 673330 120190 673570
rect 120430 673330 120540 673570
rect 120780 673330 120870 673570
rect 121110 673330 121200 673570
rect 121440 673330 121530 673570
rect 121770 673330 121790 673570
rect 110790 673240 121790 673330
rect 110790 673000 110810 673240
rect 111050 673000 111160 673240
rect 111400 673000 111490 673240
rect 111730 673000 111820 673240
rect 112060 673000 112150 673240
rect 112390 673000 112500 673240
rect 112740 673000 112830 673240
rect 113070 673000 113160 673240
rect 113400 673000 113490 673240
rect 113730 673000 113840 673240
rect 114080 673000 114170 673240
rect 114410 673000 114500 673240
rect 114740 673000 114830 673240
rect 115070 673000 115180 673240
rect 115420 673000 115510 673240
rect 115750 673000 115840 673240
rect 116080 673000 116170 673240
rect 116410 673000 116520 673240
rect 116760 673000 116850 673240
rect 117090 673000 117180 673240
rect 117420 673000 117510 673240
rect 117750 673000 117860 673240
rect 118100 673000 118190 673240
rect 118430 673000 118520 673240
rect 118760 673000 118850 673240
rect 119090 673000 119200 673240
rect 119440 673000 119530 673240
rect 119770 673000 119860 673240
rect 120100 673000 120190 673240
rect 120430 673000 120540 673240
rect 120780 673000 120870 673240
rect 121110 673000 121200 673240
rect 121440 673000 121530 673240
rect 121770 673000 121790 673240
rect 110790 672910 121790 673000
rect 110790 672670 110810 672910
rect 111050 672670 111160 672910
rect 111400 672670 111490 672910
rect 111730 672670 111820 672910
rect 112060 672670 112150 672910
rect 112390 672670 112500 672910
rect 112740 672670 112830 672910
rect 113070 672670 113160 672910
rect 113400 672670 113490 672910
rect 113730 672670 113840 672910
rect 114080 672670 114170 672910
rect 114410 672670 114500 672910
rect 114740 672670 114830 672910
rect 115070 672670 115180 672910
rect 115420 672670 115510 672910
rect 115750 672670 115840 672910
rect 116080 672670 116170 672910
rect 116410 672670 116520 672910
rect 116760 672670 116850 672910
rect 117090 672670 117180 672910
rect 117420 672670 117510 672910
rect 117750 672670 117860 672910
rect 118100 672670 118190 672910
rect 118430 672670 118520 672910
rect 118760 672670 118850 672910
rect 119090 672670 119200 672910
rect 119440 672670 119530 672910
rect 119770 672670 119860 672910
rect 120100 672670 120190 672910
rect 120430 672670 120540 672910
rect 120780 672670 120870 672910
rect 121110 672670 121200 672910
rect 121440 672670 121530 672910
rect 121770 672670 121790 672910
rect 110790 672560 121790 672670
rect 110790 672320 110810 672560
rect 111050 672320 111160 672560
rect 111400 672320 111490 672560
rect 111730 672320 111820 672560
rect 112060 672320 112150 672560
rect 112390 672320 112500 672560
rect 112740 672320 112830 672560
rect 113070 672320 113160 672560
rect 113400 672320 113490 672560
rect 113730 672320 113840 672560
rect 114080 672320 114170 672560
rect 114410 672320 114500 672560
rect 114740 672320 114830 672560
rect 115070 672320 115180 672560
rect 115420 672320 115510 672560
rect 115750 672320 115840 672560
rect 116080 672320 116170 672560
rect 116410 672320 116520 672560
rect 116760 672320 116850 672560
rect 117090 672320 117180 672560
rect 117420 672320 117510 672560
rect 117750 672320 117860 672560
rect 118100 672320 118190 672560
rect 118430 672320 118520 672560
rect 118760 672320 118850 672560
rect 119090 672320 119200 672560
rect 119440 672320 119530 672560
rect 119770 672320 119860 672560
rect 120100 672320 120190 672560
rect 120430 672320 120540 672560
rect 120780 672320 120870 672560
rect 121110 672320 121200 672560
rect 121440 672320 121530 672560
rect 121770 672320 121790 672560
rect 110790 672300 121790 672320
rect 122170 683280 133170 683300
rect 122170 683040 122190 683280
rect 122430 683040 122540 683280
rect 122780 683040 122870 683280
rect 123110 683040 123200 683280
rect 123440 683040 123530 683280
rect 123770 683040 123880 683280
rect 124120 683040 124210 683280
rect 124450 683040 124540 683280
rect 124780 683040 124870 683280
rect 125110 683040 125220 683280
rect 125460 683040 125550 683280
rect 125790 683040 125880 683280
rect 126120 683040 126210 683280
rect 126450 683040 126560 683280
rect 126800 683040 126890 683280
rect 127130 683040 127220 683280
rect 127460 683040 127550 683280
rect 127790 683040 127900 683280
rect 128140 683040 128230 683280
rect 128470 683040 128560 683280
rect 128800 683040 128890 683280
rect 129130 683040 129240 683280
rect 129480 683040 129570 683280
rect 129810 683040 129900 683280
rect 130140 683040 130230 683280
rect 130470 683040 130580 683280
rect 130820 683040 130910 683280
rect 131150 683040 131240 683280
rect 131480 683040 131570 683280
rect 131810 683040 131920 683280
rect 132160 683040 132250 683280
rect 132490 683040 132580 683280
rect 132820 683040 132910 683280
rect 133150 683040 133170 683280
rect 122170 682950 133170 683040
rect 122170 682710 122190 682950
rect 122430 682710 122540 682950
rect 122780 682710 122870 682950
rect 123110 682710 123200 682950
rect 123440 682710 123530 682950
rect 123770 682710 123880 682950
rect 124120 682710 124210 682950
rect 124450 682710 124540 682950
rect 124780 682710 124870 682950
rect 125110 682710 125220 682950
rect 125460 682710 125550 682950
rect 125790 682710 125880 682950
rect 126120 682710 126210 682950
rect 126450 682710 126560 682950
rect 126800 682710 126890 682950
rect 127130 682710 127220 682950
rect 127460 682710 127550 682950
rect 127790 682710 127900 682950
rect 128140 682710 128230 682950
rect 128470 682710 128560 682950
rect 128800 682710 128890 682950
rect 129130 682710 129240 682950
rect 129480 682710 129570 682950
rect 129810 682710 129900 682950
rect 130140 682710 130230 682950
rect 130470 682710 130580 682950
rect 130820 682710 130910 682950
rect 131150 682710 131240 682950
rect 131480 682710 131570 682950
rect 131810 682710 131920 682950
rect 132160 682710 132250 682950
rect 132490 682710 132580 682950
rect 132820 682710 132910 682950
rect 133150 682710 133170 682950
rect 122170 682620 133170 682710
rect 122170 682380 122190 682620
rect 122430 682380 122540 682620
rect 122780 682380 122870 682620
rect 123110 682380 123200 682620
rect 123440 682380 123530 682620
rect 123770 682380 123880 682620
rect 124120 682380 124210 682620
rect 124450 682380 124540 682620
rect 124780 682380 124870 682620
rect 125110 682380 125220 682620
rect 125460 682380 125550 682620
rect 125790 682380 125880 682620
rect 126120 682380 126210 682620
rect 126450 682380 126560 682620
rect 126800 682380 126890 682620
rect 127130 682380 127220 682620
rect 127460 682380 127550 682620
rect 127790 682380 127900 682620
rect 128140 682380 128230 682620
rect 128470 682380 128560 682620
rect 128800 682380 128890 682620
rect 129130 682380 129240 682620
rect 129480 682380 129570 682620
rect 129810 682380 129900 682620
rect 130140 682380 130230 682620
rect 130470 682380 130580 682620
rect 130820 682380 130910 682620
rect 131150 682380 131240 682620
rect 131480 682380 131570 682620
rect 131810 682380 131920 682620
rect 132160 682380 132250 682620
rect 132490 682380 132580 682620
rect 132820 682380 132910 682620
rect 133150 682380 133170 682620
rect 122170 682290 133170 682380
rect 122170 682050 122190 682290
rect 122430 682050 122540 682290
rect 122780 682050 122870 682290
rect 123110 682050 123200 682290
rect 123440 682050 123530 682290
rect 123770 682050 123880 682290
rect 124120 682050 124210 682290
rect 124450 682050 124540 682290
rect 124780 682050 124870 682290
rect 125110 682050 125220 682290
rect 125460 682050 125550 682290
rect 125790 682050 125880 682290
rect 126120 682050 126210 682290
rect 126450 682050 126560 682290
rect 126800 682050 126890 682290
rect 127130 682050 127220 682290
rect 127460 682050 127550 682290
rect 127790 682050 127900 682290
rect 128140 682050 128230 682290
rect 128470 682050 128560 682290
rect 128800 682050 128890 682290
rect 129130 682050 129240 682290
rect 129480 682050 129570 682290
rect 129810 682050 129900 682290
rect 130140 682050 130230 682290
rect 130470 682050 130580 682290
rect 130820 682050 130910 682290
rect 131150 682050 131240 682290
rect 131480 682050 131570 682290
rect 131810 682050 131920 682290
rect 132160 682050 132250 682290
rect 132490 682050 132580 682290
rect 132820 682050 132910 682290
rect 133150 682050 133170 682290
rect 122170 681940 133170 682050
rect 122170 681700 122190 681940
rect 122430 681700 122540 681940
rect 122780 681700 122870 681940
rect 123110 681700 123200 681940
rect 123440 681700 123530 681940
rect 123770 681700 123880 681940
rect 124120 681700 124210 681940
rect 124450 681700 124540 681940
rect 124780 681700 124870 681940
rect 125110 681700 125220 681940
rect 125460 681700 125550 681940
rect 125790 681700 125880 681940
rect 126120 681700 126210 681940
rect 126450 681700 126560 681940
rect 126800 681700 126890 681940
rect 127130 681700 127220 681940
rect 127460 681700 127550 681940
rect 127790 681700 127900 681940
rect 128140 681700 128230 681940
rect 128470 681700 128560 681940
rect 128800 681700 128890 681940
rect 129130 681700 129240 681940
rect 129480 681700 129570 681940
rect 129810 681700 129900 681940
rect 130140 681700 130230 681940
rect 130470 681700 130580 681940
rect 130820 681700 130910 681940
rect 131150 681700 131240 681940
rect 131480 681700 131570 681940
rect 131810 681700 131920 681940
rect 132160 681700 132250 681940
rect 132490 681700 132580 681940
rect 132820 681700 132910 681940
rect 133150 681700 133170 681940
rect 122170 681610 133170 681700
rect 122170 681370 122190 681610
rect 122430 681370 122540 681610
rect 122780 681370 122870 681610
rect 123110 681370 123200 681610
rect 123440 681370 123530 681610
rect 123770 681370 123880 681610
rect 124120 681370 124210 681610
rect 124450 681370 124540 681610
rect 124780 681370 124870 681610
rect 125110 681370 125220 681610
rect 125460 681370 125550 681610
rect 125790 681370 125880 681610
rect 126120 681370 126210 681610
rect 126450 681370 126560 681610
rect 126800 681370 126890 681610
rect 127130 681370 127220 681610
rect 127460 681370 127550 681610
rect 127790 681370 127900 681610
rect 128140 681370 128230 681610
rect 128470 681370 128560 681610
rect 128800 681370 128890 681610
rect 129130 681370 129240 681610
rect 129480 681370 129570 681610
rect 129810 681370 129900 681610
rect 130140 681370 130230 681610
rect 130470 681370 130580 681610
rect 130820 681370 130910 681610
rect 131150 681370 131240 681610
rect 131480 681370 131570 681610
rect 131810 681370 131920 681610
rect 132160 681370 132250 681610
rect 132490 681370 132580 681610
rect 132820 681370 132910 681610
rect 133150 681370 133170 681610
rect 122170 681280 133170 681370
rect 122170 681040 122190 681280
rect 122430 681040 122540 681280
rect 122780 681040 122870 681280
rect 123110 681040 123200 681280
rect 123440 681040 123530 681280
rect 123770 681040 123880 681280
rect 124120 681040 124210 681280
rect 124450 681040 124540 681280
rect 124780 681040 124870 681280
rect 125110 681040 125220 681280
rect 125460 681040 125550 681280
rect 125790 681040 125880 681280
rect 126120 681040 126210 681280
rect 126450 681040 126560 681280
rect 126800 681040 126890 681280
rect 127130 681040 127220 681280
rect 127460 681040 127550 681280
rect 127790 681040 127900 681280
rect 128140 681040 128230 681280
rect 128470 681040 128560 681280
rect 128800 681040 128890 681280
rect 129130 681040 129240 681280
rect 129480 681040 129570 681280
rect 129810 681040 129900 681280
rect 130140 681040 130230 681280
rect 130470 681040 130580 681280
rect 130820 681040 130910 681280
rect 131150 681040 131240 681280
rect 131480 681040 131570 681280
rect 131810 681040 131920 681280
rect 132160 681040 132250 681280
rect 132490 681040 132580 681280
rect 132820 681040 132910 681280
rect 133150 681040 133170 681280
rect 122170 680950 133170 681040
rect 122170 680710 122190 680950
rect 122430 680710 122540 680950
rect 122780 680710 122870 680950
rect 123110 680710 123200 680950
rect 123440 680710 123530 680950
rect 123770 680710 123880 680950
rect 124120 680710 124210 680950
rect 124450 680710 124540 680950
rect 124780 680710 124870 680950
rect 125110 680710 125220 680950
rect 125460 680710 125550 680950
rect 125790 680710 125880 680950
rect 126120 680710 126210 680950
rect 126450 680710 126560 680950
rect 126800 680710 126890 680950
rect 127130 680710 127220 680950
rect 127460 680710 127550 680950
rect 127790 680710 127900 680950
rect 128140 680710 128230 680950
rect 128470 680710 128560 680950
rect 128800 680710 128890 680950
rect 129130 680710 129240 680950
rect 129480 680710 129570 680950
rect 129810 680710 129900 680950
rect 130140 680710 130230 680950
rect 130470 680710 130580 680950
rect 130820 680710 130910 680950
rect 131150 680710 131240 680950
rect 131480 680710 131570 680950
rect 131810 680710 131920 680950
rect 132160 680710 132250 680950
rect 132490 680710 132580 680950
rect 132820 680710 132910 680950
rect 133150 680710 133170 680950
rect 122170 680600 133170 680710
rect 122170 680360 122190 680600
rect 122430 680360 122540 680600
rect 122780 680360 122870 680600
rect 123110 680360 123200 680600
rect 123440 680360 123530 680600
rect 123770 680360 123880 680600
rect 124120 680360 124210 680600
rect 124450 680360 124540 680600
rect 124780 680360 124870 680600
rect 125110 680360 125220 680600
rect 125460 680360 125550 680600
rect 125790 680360 125880 680600
rect 126120 680360 126210 680600
rect 126450 680360 126560 680600
rect 126800 680360 126890 680600
rect 127130 680360 127220 680600
rect 127460 680360 127550 680600
rect 127790 680360 127900 680600
rect 128140 680360 128230 680600
rect 128470 680360 128560 680600
rect 128800 680360 128890 680600
rect 129130 680360 129240 680600
rect 129480 680360 129570 680600
rect 129810 680360 129900 680600
rect 130140 680360 130230 680600
rect 130470 680360 130580 680600
rect 130820 680360 130910 680600
rect 131150 680360 131240 680600
rect 131480 680360 131570 680600
rect 131810 680360 131920 680600
rect 132160 680360 132250 680600
rect 132490 680360 132580 680600
rect 132820 680360 132910 680600
rect 133150 680360 133170 680600
rect 122170 680270 133170 680360
rect 122170 680030 122190 680270
rect 122430 680030 122540 680270
rect 122780 680030 122870 680270
rect 123110 680030 123200 680270
rect 123440 680030 123530 680270
rect 123770 680030 123880 680270
rect 124120 680030 124210 680270
rect 124450 680030 124540 680270
rect 124780 680030 124870 680270
rect 125110 680030 125220 680270
rect 125460 680030 125550 680270
rect 125790 680030 125880 680270
rect 126120 680030 126210 680270
rect 126450 680030 126560 680270
rect 126800 680030 126890 680270
rect 127130 680030 127220 680270
rect 127460 680030 127550 680270
rect 127790 680030 127900 680270
rect 128140 680030 128230 680270
rect 128470 680030 128560 680270
rect 128800 680030 128890 680270
rect 129130 680030 129240 680270
rect 129480 680030 129570 680270
rect 129810 680030 129900 680270
rect 130140 680030 130230 680270
rect 130470 680030 130580 680270
rect 130820 680030 130910 680270
rect 131150 680030 131240 680270
rect 131480 680030 131570 680270
rect 131810 680030 131920 680270
rect 132160 680030 132250 680270
rect 132490 680030 132580 680270
rect 132820 680030 132910 680270
rect 133150 680030 133170 680270
rect 122170 679940 133170 680030
rect 122170 679700 122190 679940
rect 122430 679700 122540 679940
rect 122780 679700 122870 679940
rect 123110 679700 123200 679940
rect 123440 679700 123530 679940
rect 123770 679700 123880 679940
rect 124120 679700 124210 679940
rect 124450 679700 124540 679940
rect 124780 679700 124870 679940
rect 125110 679700 125220 679940
rect 125460 679700 125550 679940
rect 125790 679700 125880 679940
rect 126120 679700 126210 679940
rect 126450 679700 126560 679940
rect 126800 679700 126890 679940
rect 127130 679700 127220 679940
rect 127460 679700 127550 679940
rect 127790 679700 127900 679940
rect 128140 679700 128230 679940
rect 128470 679700 128560 679940
rect 128800 679700 128890 679940
rect 129130 679700 129240 679940
rect 129480 679700 129570 679940
rect 129810 679700 129900 679940
rect 130140 679700 130230 679940
rect 130470 679700 130580 679940
rect 130820 679700 130910 679940
rect 131150 679700 131240 679940
rect 131480 679700 131570 679940
rect 131810 679700 131920 679940
rect 132160 679700 132250 679940
rect 132490 679700 132580 679940
rect 132820 679700 132910 679940
rect 133150 679700 133170 679940
rect 122170 679610 133170 679700
rect 122170 679370 122190 679610
rect 122430 679370 122540 679610
rect 122780 679370 122870 679610
rect 123110 679370 123200 679610
rect 123440 679370 123530 679610
rect 123770 679370 123880 679610
rect 124120 679370 124210 679610
rect 124450 679370 124540 679610
rect 124780 679370 124870 679610
rect 125110 679370 125220 679610
rect 125460 679370 125550 679610
rect 125790 679370 125880 679610
rect 126120 679370 126210 679610
rect 126450 679370 126560 679610
rect 126800 679370 126890 679610
rect 127130 679370 127220 679610
rect 127460 679370 127550 679610
rect 127790 679370 127900 679610
rect 128140 679370 128230 679610
rect 128470 679370 128560 679610
rect 128800 679370 128890 679610
rect 129130 679370 129240 679610
rect 129480 679370 129570 679610
rect 129810 679370 129900 679610
rect 130140 679370 130230 679610
rect 130470 679370 130580 679610
rect 130820 679370 130910 679610
rect 131150 679370 131240 679610
rect 131480 679370 131570 679610
rect 131810 679370 131920 679610
rect 132160 679370 132250 679610
rect 132490 679370 132580 679610
rect 132820 679370 132910 679610
rect 133150 679370 133170 679610
rect 122170 679260 133170 679370
rect 122170 679020 122190 679260
rect 122430 679020 122540 679260
rect 122780 679020 122870 679260
rect 123110 679020 123200 679260
rect 123440 679020 123530 679260
rect 123770 679020 123880 679260
rect 124120 679020 124210 679260
rect 124450 679020 124540 679260
rect 124780 679020 124870 679260
rect 125110 679020 125220 679260
rect 125460 679020 125550 679260
rect 125790 679020 125880 679260
rect 126120 679020 126210 679260
rect 126450 679020 126560 679260
rect 126800 679020 126890 679260
rect 127130 679020 127220 679260
rect 127460 679020 127550 679260
rect 127790 679020 127900 679260
rect 128140 679020 128230 679260
rect 128470 679020 128560 679260
rect 128800 679020 128890 679260
rect 129130 679020 129240 679260
rect 129480 679020 129570 679260
rect 129810 679020 129900 679260
rect 130140 679020 130230 679260
rect 130470 679020 130580 679260
rect 130820 679020 130910 679260
rect 131150 679020 131240 679260
rect 131480 679020 131570 679260
rect 131810 679020 131920 679260
rect 132160 679020 132250 679260
rect 132490 679020 132580 679260
rect 132820 679020 132910 679260
rect 133150 679020 133170 679260
rect 122170 678930 133170 679020
rect 122170 678690 122190 678930
rect 122430 678690 122540 678930
rect 122780 678690 122870 678930
rect 123110 678690 123200 678930
rect 123440 678690 123530 678930
rect 123770 678690 123880 678930
rect 124120 678690 124210 678930
rect 124450 678690 124540 678930
rect 124780 678690 124870 678930
rect 125110 678690 125220 678930
rect 125460 678690 125550 678930
rect 125790 678690 125880 678930
rect 126120 678690 126210 678930
rect 126450 678690 126560 678930
rect 126800 678690 126890 678930
rect 127130 678690 127220 678930
rect 127460 678690 127550 678930
rect 127790 678690 127900 678930
rect 128140 678690 128230 678930
rect 128470 678690 128560 678930
rect 128800 678690 128890 678930
rect 129130 678690 129240 678930
rect 129480 678690 129570 678930
rect 129810 678690 129900 678930
rect 130140 678690 130230 678930
rect 130470 678690 130580 678930
rect 130820 678690 130910 678930
rect 131150 678690 131240 678930
rect 131480 678690 131570 678930
rect 131810 678690 131920 678930
rect 132160 678690 132250 678930
rect 132490 678690 132580 678930
rect 132820 678690 132910 678930
rect 133150 678690 133170 678930
rect 122170 678600 133170 678690
rect 122170 678360 122190 678600
rect 122430 678360 122540 678600
rect 122780 678360 122870 678600
rect 123110 678360 123200 678600
rect 123440 678360 123530 678600
rect 123770 678360 123880 678600
rect 124120 678360 124210 678600
rect 124450 678360 124540 678600
rect 124780 678360 124870 678600
rect 125110 678360 125220 678600
rect 125460 678360 125550 678600
rect 125790 678360 125880 678600
rect 126120 678360 126210 678600
rect 126450 678360 126560 678600
rect 126800 678360 126890 678600
rect 127130 678360 127220 678600
rect 127460 678360 127550 678600
rect 127790 678360 127900 678600
rect 128140 678360 128230 678600
rect 128470 678360 128560 678600
rect 128800 678360 128890 678600
rect 129130 678360 129240 678600
rect 129480 678360 129570 678600
rect 129810 678360 129900 678600
rect 130140 678360 130230 678600
rect 130470 678360 130580 678600
rect 130820 678360 130910 678600
rect 131150 678360 131240 678600
rect 131480 678360 131570 678600
rect 131810 678360 131920 678600
rect 132160 678360 132250 678600
rect 132490 678360 132580 678600
rect 132820 678360 132910 678600
rect 133150 678360 133170 678600
rect 122170 678270 133170 678360
rect 122170 678030 122190 678270
rect 122430 678030 122540 678270
rect 122780 678030 122870 678270
rect 123110 678030 123200 678270
rect 123440 678030 123530 678270
rect 123770 678030 123880 678270
rect 124120 678030 124210 678270
rect 124450 678030 124540 678270
rect 124780 678030 124870 678270
rect 125110 678030 125220 678270
rect 125460 678030 125550 678270
rect 125790 678030 125880 678270
rect 126120 678030 126210 678270
rect 126450 678030 126560 678270
rect 126800 678030 126890 678270
rect 127130 678030 127220 678270
rect 127460 678030 127550 678270
rect 127790 678030 127900 678270
rect 128140 678030 128230 678270
rect 128470 678030 128560 678270
rect 128800 678030 128890 678270
rect 129130 678030 129240 678270
rect 129480 678030 129570 678270
rect 129810 678030 129900 678270
rect 130140 678030 130230 678270
rect 130470 678030 130580 678270
rect 130820 678030 130910 678270
rect 131150 678030 131240 678270
rect 131480 678030 131570 678270
rect 131810 678030 131920 678270
rect 132160 678030 132250 678270
rect 132490 678030 132580 678270
rect 132820 678030 132910 678270
rect 133150 678030 133170 678270
rect 122170 677920 133170 678030
rect 122170 677680 122190 677920
rect 122430 677680 122540 677920
rect 122780 677680 122870 677920
rect 123110 677680 123200 677920
rect 123440 677680 123530 677920
rect 123770 677680 123880 677920
rect 124120 677680 124210 677920
rect 124450 677680 124540 677920
rect 124780 677680 124870 677920
rect 125110 677680 125220 677920
rect 125460 677680 125550 677920
rect 125790 677680 125880 677920
rect 126120 677680 126210 677920
rect 126450 677680 126560 677920
rect 126800 677680 126890 677920
rect 127130 677680 127220 677920
rect 127460 677680 127550 677920
rect 127790 677680 127900 677920
rect 128140 677680 128230 677920
rect 128470 677680 128560 677920
rect 128800 677680 128890 677920
rect 129130 677680 129240 677920
rect 129480 677680 129570 677920
rect 129810 677680 129900 677920
rect 130140 677680 130230 677920
rect 130470 677680 130580 677920
rect 130820 677680 130910 677920
rect 131150 677680 131240 677920
rect 131480 677680 131570 677920
rect 131810 677680 131920 677920
rect 132160 677680 132250 677920
rect 132490 677680 132580 677920
rect 132820 677680 132910 677920
rect 133150 677680 133170 677920
rect 122170 677590 133170 677680
rect 122170 677350 122190 677590
rect 122430 677350 122540 677590
rect 122780 677350 122870 677590
rect 123110 677350 123200 677590
rect 123440 677350 123530 677590
rect 123770 677350 123880 677590
rect 124120 677350 124210 677590
rect 124450 677350 124540 677590
rect 124780 677350 124870 677590
rect 125110 677350 125220 677590
rect 125460 677350 125550 677590
rect 125790 677350 125880 677590
rect 126120 677350 126210 677590
rect 126450 677350 126560 677590
rect 126800 677350 126890 677590
rect 127130 677350 127220 677590
rect 127460 677350 127550 677590
rect 127790 677350 127900 677590
rect 128140 677350 128230 677590
rect 128470 677350 128560 677590
rect 128800 677350 128890 677590
rect 129130 677350 129240 677590
rect 129480 677350 129570 677590
rect 129810 677350 129900 677590
rect 130140 677350 130230 677590
rect 130470 677350 130580 677590
rect 130820 677350 130910 677590
rect 131150 677350 131240 677590
rect 131480 677350 131570 677590
rect 131810 677350 131920 677590
rect 132160 677350 132250 677590
rect 132490 677350 132580 677590
rect 132820 677350 132910 677590
rect 133150 677350 133170 677590
rect 122170 677260 133170 677350
rect 122170 677020 122190 677260
rect 122430 677020 122540 677260
rect 122780 677020 122870 677260
rect 123110 677020 123200 677260
rect 123440 677020 123530 677260
rect 123770 677020 123880 677260
rect 124120 677020 124210 677260
rect 124450 677020 124540 677260
rect 124780 677020 124870 677260
rect 125110 677020 125220 677260
rect 125460 677020 125550 677260
rect 125790 677020 125880 677260
rect 126120 677020 126210 677260
rect 126450 677020 126560 677260
rect 126800 677020 126890 677260
rect 127130 677020 127220 677260
rect 127460 677020 127550 677260
rect 127790 677020 127900 677260
rect 128140 677020 128230 677260
rect 128470 677020 128560 677260
rect 128800 677020 128890 677260
rect 129130 677020 129240 677260
rect 129480 677020 129570 677260
rect 129810 677020 129900 677260
rect 130140 677020 130230 677260
rect 130470 677020 130580 677260
rect 130820 677020 130910 677260
rect 131150 677020 131240 677260
rect 131480 677020 131570 677260
rect 131810 677020 131920 677260
rect 132160 677020 132250 677260
rect 132490 677020 132580 677260
rect 132820 677020 132910 677260
rect 133150 677020 133170 677260
rect 122170 676930 133170 677020
rect 122170 676690 122190 676930
rect 122430 676690 122540 676930
rect 122780 676690 122870 676930
rect 123110 676690 123200 676930
rect 123440 676690 123530 676930
rect 123770 676690 123880 676930
rect 124120 676690 124210 676930
rect 124450 676690 124540 676930
rect 124780 676690 124870 676930
rect 125110 676690 125220 676930
rect 125460 676690 125550 676930
rect 125790 676690 125880 676930
rect 126120 676690 126210 676930
rect 126450 676690 126560 676930
rect 126800 676690 126890 676930
rect 127130 676690 127220 676930
rect 127460 676690 127550 676930
rect 127790 676690 127900 676930
rect 128140 676690 128230 676930
rect 128470 676690 128560 676930
rect 128800 676690 128890 676930
rect 129130 676690 129240 676930
rect 129480 676690 129570 676930
rect 129810 676690 129900 676930
rect 130140 676690 130230 676930
rect 130470 676690 130580 676930
rect 130820 676690 130910 676930
rect 131150 676690 131240 676930
rect 131480 676690 131570 676930
rect 131810 676690 131920 676930
rect 132160 676690 132250 676930
rect 132490 676690 132580 676930
rect 132820 676690 132910 676930
rect 133150 676690 133170 676930
rect 122170 676580 133170 676690
rect 122170 676340 122190 676580
rect 122430 676340 122540 676580
rect 122780 676340 122870 676580
rect 123110 676340 123200 676580
rect 123440 676340 123530 676580
rect 123770 676340 123880 676580
rect 124120 676340 124210 676580
rect 124450 676340 124540 676580
rect 124780 676340 124870 676580
rect 125110 676340 125220 676580
rect 125460 676340 125550 676580
rect 125790 676340 125880 676580
rect 126120 676340 126210 676580
rect 126450 676340 126560 676580
rect 126800 676340 126890 676580
rect 127130 676340 127220 676580
rect 127460 676340 127550 676580
rect 127790 676340 127900 676580
rect 128140 676340 128230 676580
rect 128470 676340 128560 676580
rect 128800 676340 128890 676580
rect 129130 676340 129240 676580
rect 129480 676340 129570 676580
rect 129810 676340 129900 676580
rect 130140 676340 130230 676580
rect 130470 676340 130580 676580
rect 130820 676340 130910 676580
rect 131150 676340 131240 676580
rect 131480 676340 131570 676580
rect 131810 676340 131920 676580
rect 132160 676340 132250 676580
rect 132490 676340 132580 676580
rect 132820 676340 132910 676580
rect 133150 676340 133170 676580
rect 122170 676250 133170 676340
rect 122170 676010 122190 676250
rect 122430 676010 122540 676250
rect 122780 676010 122870 676250
rect 123110 676010 123200 676250
rect 123440 676010 123530 676250
rect 123770 676010 123880 676250
rect 124120 676010 124210 676250
rect 124450 676010 124540 676250
rect 124780 676010 124870 676250
rect 125110 676010 125220 676250
rect 125460 676010 125550 676250
rect 125790 676010 125880 676250
rect 126120 676010 126210 676250
rect 126450 676010 126560 676250
rect 126800 676010 126890 676250
rect 127130 676010 127220 676250
rect 127460 676010 127550 676250
rect 127790 676010 127900 676250
rect 128140 676010 128230 676250
rect 128470 676010 128560 676250
rect 128800 676010 128890 676250
rect 129130 676010 129240 676250
rect 129480 676010 129570 676250
rect 129810 676010 129900 676250
rect 130140 676010 130230 676250
rect 130470 676010 130580 676250
rect 130820 676010 130910 676250
rect 131150 676010 131240 676250
rect 131480 676010 131570 676250
rect 131810 676010 131920 676250
rect 132160 676010 132250 676250
rect 132490 676010 132580 676250
rect 132820 676010 132910 676250
rect 133150 676010 133170 676250
rect 122170 675920 133170 676010
rect 122170 675680 122190 675920
rect 122430 675680 122540 675920
rect 122780 675680 122870 675920
rect 123110 675680 123200 675920
rect 123440 675680 123530 675920
rect 123770 675680 123880 675920
rect 124120 675680 124210 675920
rect 124450 675680 124540 675920
rect 124780 675680 124870 675920
rect 125110 675680 125220 675920
rect 125460 675680 125550 675920
rect 125790 675680 125880 675920
rect 126120 675680 126210 675920
rect 126450 675680 126560 675920
rect 126800 675680 126890 675920
rect 127130 675680 127220 675920
rect 127460 675680 127550 675920
rect 127790 675680 127900 675920
rect 128140 675680 128230 675920
rect 128470 675680 128560 675920
rect 128800 675680 128890 675920
rect 129130 675680 129240 675920
rect 129480 675680 129570 675920
rect 129810 675680 129900 675920
rect 130140 675680 130230 675920
rect 130470 675680 130580 675920
rect 130820 675680 130910 675920
rect 131150 675680 131240 675920
rect 131480 675680 131570 675920
rect 131810 675680 131920 675920
rect 132160 675680 132250 675920
rect 132490 675680 132580 675920
rect 132820 675680 132910 675920
rect 133150 675680 133170 675920
rect 122170 675590 133170 675680
rect 122170 675350 122190 675590
rect 122430 675350 122540 675590
rect 122780 675350 122870 675590
rect 123110 675350 123200 675590
rect 123440 675350 123530 675590
rect 123770 675350 123880 675590
rect 124120 675350 124210 675590
rect 124450 675350 124540 675590
rect 124780 675350 124870 675590
rect 125110 675350 125220 675590
rect 125460 675350 125550 675590
rect 125790 675350 125880 675590
rect 126120 675350 126210 675590
rect 126450 675350 126560 675590
rect 126800 675350 126890 675590
rect 127130 675350 127220 675590
rect 127460 675350 127550 675590
rect 127790 675350 127900 675590
rect 128140 675350 128230 675590
rect 128470 675350 128560 675590
rect 128800 675350 128890 675590
rect 129130 675350 129240 675590
rect 129480 675350 129570 675590
rect 129810 675350 129900 675590
rect 130140 675350 130230 675590
rect 130470 675350 130580 675590
rect 130820 675350 130910 675590
rect 131150 675350 131240 675590
rect 131480 675350 131570 675590
rect 131810 675350 131920 675590
rect 132160 675350 132250 675590
rect 132490 675350 132580 675590
rect 132820 675350 132910 675590
rect 133150 675350 133170 675590
rect 122170 675240 133170 675350
rect 122170 675000 122190 675240
rect 122430 675000 122540 675240
rect 122780 675000 122870 675240
rect 123110 675000 123200 675240
rect 123440 675000 123530 675240
rect 123770 675000 123880 675240
rect 124120 675000 124210 675240
rect 124450 675000 124540 675240
rect 124780 675000 124870 675240
rect 125110 675000 125220 675240
rect 125460 675000 125550 675240
rect 125790 675000 125880 675240
rect 126120 675000 126210 675240
rect 126450 675000 126560 675240
rect 126800 675000 126890 675240
rect 127130 675000 127220 675240
rect 127460 675000 127550 675240
rect 127790 675000 127900 675240
rect 128140 675000 128230 675240
rect 128470 675000 128560 675240
rect 128800 675000 128890 675240
rect 129130 675000 129240 675240
rect 129480 675000 129570 675240
rect 129810 675000 129900 675240
rect 130140 675000 130230 675240
rect 130470 675000 130580 675240
rect 130820 675000 130910 675240
rect 131150 675000 131240 675240
rect 131480 675000 131570 675240
rect 131810 675000 131920 675240
rect 132160 675000 132250 675240
rect 132490 675000 132580 675240
rect 132820 675000 132910 675240
rect 133150 675000 133170 675240
rect 122170 674910 133170 675000
rect 122170 674670 122190 674910
rect 122430 674670 122540 674910
rect 122780 674670 122870 674910
rect 123110 674670 123200 674910
rect 123440 674670 123530 674910
rect 123770 674670 123880 674910
rect 124120 674670 124210 674910
rect 124450 674670 124540 674910
rect 124780 674670 124870 674910
rect 125110 674670 125220 674910
rect 125460 674670 125550 674910
rect 125790 674670 125880 674910
rect 126120 674670 126210 674910
rect 126450 674670 126560 674910
rect 126800 674670 126890 674910
rect 127130 674670 127220 674910
rect 127460 674670 127550 674910
rect 127790 674670 127900 674910
rect 128140 674670 128230 674910
rect 128470 674670 128560 674910
rect 128800 674670 128890 674910
rect 129130 674670 129240 674910
rect 129480 674670 129570 674910
rect 129810 674670 129900 674910
rect 130140 674670 130230 674910
rect 130470 674670 130580 674910
rect 130820 674670 130910 674910
rect 131150 674670 131240 674910
rect 131480 674670 131570 674910
rect 131810 674670 131920 674910
rect 132160 674670 132250 674910
rect 132490 674670 132580 674910
rect 132820 674670 132910 674910
rect 133150 674670 133170 674910
rect 122170 674580 133170 674670
rect 122170 674340 122190 674580
rect 122430 674340 122540 674580
rect 122780 674340 122870 674580
rect 123110 674340 123200 674580
rect 123440 674340 123530 674580
rect 123770 674340 123880 674580
rect 124120 674340 124210 674580
rect 124450 674340 124540 674580
rect 124780 674340 124870 674580
rect 125110 674340 125220 674580
rect 125460 674340 125550 674580
rect 125790 674340 125880 674580
rect 126120 674340 126210 674580
rect 126450 674340 126560 674580
rect 126800 674340 126890 674580
rect 127130 674340 127220 674580
rect 127460 674340 127550 674580
rect 127790 674340 127900 674580
rect 128140 674340 128230 674580
rect 128470 674340 128560 674580
rect 128800 674340 128890 674580
rect 129130 674340 129240 674580
rect 129480 674340 129570 674580
rect 129810 674340 129900 674580
rect 130140 674340 130230 674580
rect 130470 674340 130580 674580
rect 130820 674340 130910 674580
rect 131150 674340 131240 674580
rect 131480 674340 131570 674580
rect 131810 674340 131920 674580
rect 132160 674340 132250 674580
rect 132490 674340 132580 674580
rect 132820 674340 132910 674580
rect 133150 674340 133170 674580
rect 122170 674250 133170 674340
rect 122170 674010 122190 674250
rect 122430 674010 122540 674250
rect 122780 674010 122870 674250
rect 123110 674010 123200 674250
rect 123440 674010 123530 674250
rect 123770 674010 123880 674250
rect 124120 674010 124210 674250
rect 124450 674010 124540 674250
rect 124780 674010 124870 674250
rect 125110 674010 125220 674250
rect 125460 674010 125550 674250
rect 125790 674010 125880 674250
rect 126120 674010 126210 674250
rect 126450 674010 126560 674250
rect 126800 674010 126890 674250
rect 127130 674010 127220 674250
rect 127460 674010 127550 674250
rect 127790 674010 127900 674250
rect 128140 674010 128230 674250
rect 128470 674010 128560 674250
rect 128800 674010 128890 674250
rect 129130 674010 129240 674250
rect 129480 674010 129570 674250
rect 129810 674010 129900 674250
rect 130140 674010 130230 674250
rect 130470 674010 130580 674250
rect 130820 674010 130910 674250
rect 131150 674010 131240 674250
rect 131480 674010 131570 674250
rect 131810 674010 131920 674250
rect 132160 674010 132250 674250
rect 132490 674010 132580 674250
rect 132820 674010 132910 674250
rect 133150 674010 133170 674250
rect 122170 673900 133170 674010
rect 122170 673660 122190 673900
rect 122430 673660 122540 673900
rect 122780 673660 122870 673900
rect 123110 673660 123200 673900
rect 123440 673660 123530 673900
rect 123770 673660 123880 673900
rect 124120 673660 124210 673900
rect 124450 673660 124540 673900
rect 124780 673660 124870 673900
rect 125110 673660 125220 673900
rect 125460 673660 125550 673900
rect 125790 673660 125880 673900
rect 126120 673660 126210 673900
rect 126450 673660 126560 673900
rect 126800 673660 126890 673900
rect 127130 673660 127220 673900
rect 127460 673660 127550 673900
rect 127790 673660 127900 673900
rect 128140 673660 128230 673900
rect 128470 673660 128560 673900
rect 128800 673660 128890 673900
rect 129130 673660 129240 673900
rect 129480 673660 129570 673900
rect 129810 673660 129900 673900
rect 130140 673660 130230 673900
rect 130470 673660 130580 673900
rect 130820 673660 130910 673900
rect 131150 673660 131240 673900
rect 131480 673660 131570 673900
rect 131810 673660 131920 673900
rect 132160 673660 132250 673900
rect 132490 673660 132580 673900
rect 132820 673660 132910 673900
rect 133150 673660 133170 673900
rect 122170 673570 133170 673660
rect 122170 673330 122190 673570
rect 122430 673330 122540 673570
rect 122780 673330 122870 673570
rect 123110 673330 123200 673570
rect 123440 673330 123530 673570
rect 123770 673330 123880 673570
rect 124120 673330 124210 673570
rect 124450 673330 124540 673570
rect 124780 673330 124870 673570
rect 125110 673330 125220 673570
rect 125460 673330 125550 673570
rect 125790 673330 125880 673570
rect 126120 673330 126210 673570
rect 126450 673330 126560 673570
rect 126800 673330 126890 673570
rect 127130 673330 127220 673570
rect 127460 673330 127550 673570
rect 127790 673330 127900 673570
rect 128140 673330 128230 673570
rect 128470 673330 128560 673570
rect 128800 673330 128890 673570
rect 129130 673330 129240 673570
rect 129480 673330 129570 673570
rect 129810 673330 129900 673570
rect 130140 673330 130230 673570
rect 130470 673330 130580 673570
rect 130820 673330 130910 673570
rect 131150 673330 131240 673570
rect 131480 673330 131570 673570
rect 131810 673330 131920 673570
rect 132160 673330 132250 673570
rect 132490 673330 132580 673570
rect 132820 673330 132910 673570
rect 133150 673330 133170 673570
rect 122170 673240 133170 673330
rect 122170 673000 122190 673240
rect 122430 673000 122540 673240
rect 122780 673000 122870 673240
rect 123110 673000 123200 673240
rect 123440 673000 123530 673240
rect 123770 673000 123880 673240
rect 124120 673000 124210 673240
rect 124450 673000 124540 673240
rect 124780 673000 124870 673240
rect 125110 673000 125220 673240
rect 125460 673000 125550 673240
rect 125790 673000 125880 673240
rect 126120 673000 126210 673240
rect 126450 673000 126560 673240
rect 126800 673000 126890 673240
rect 127130 673000 127220 673240
rect 127460 673000 127550 673240
rect 127790 673000 127900 673240
rect 128140 673000 128230 673240
rect 128470 673000 128560 673240
rect 128800 673000 128890 673240
rect 129130 673000 129240 673240
rect 129480 673000 129570 673240
rect 129810 673000 129900 673240
rect 130140 673000 130230 673240
rect 130470 673000 130580 673240
rect 130820 673000 130910 673240
rect 131150 673000 131240 673240
rect 131480 673000 131570 673240
rect 131810 673000 131920 673240
rect 132160 673000 132250 673240
rect 132490 673000 132580 673240
rect 132820 673000 132910 673240
rect 133150 673000 133170 673240
rect 122170 672910 133170 673000
rect 122170 672670 122190 672910
rect 122430 672670 122540 672910
rect 122780 672670 122870 672910
rect 123110 672670 123200 672910
rect 123440 672670 123530 672910
rect 123770 672670 123880 672910
rect 124120 672670 124210 672910
rect 124450 672670 124540 672910
rect 124780 672670 124870 672910
rect 125110 672670 125220 672910
rect 125460 672670 125550 672910
rect 125790 672670 125880 672910
rect 126120 672670 126210 672910
rect 126450 672670 126560 672910
rect 126800 672670 126890 672910
rect 127130 672670 127220 672910
rect 127460 672670 127550 672910
rect 127790 672670 127900 672910
rect 128140 672670 128230 672910
rect 128470 672670 128560 672910
rect 128800 672670 128890 672910
rect 129130 672670 129240 672910
rect 129480 672670 129570 672910
rect 129810 672670 129900 672910
rect 130140 672670 130230 672910
rect 130470 672670 130580 672910
rect 130820 672670 130910 672910
rect 131150 672670 131240 672910
rect 131480 672670 131570 672910
rect 131810 672670 131920 672910
rect 132160 672670 132250 672910
rect 132490 672670 132580 672910
rect 132820 672670 132910 672910
rect 133150 672670 133170 672910
rect 122170 672560 133170 672670
rect 122170 672320 122190 672560
rect 122430 672320 122540 672560
rect 122780 672320 122870 672560
rect 123110 672320 123200 672560
rect 123440 672320 123530 672560
rect 123770 672320 123880 672560
rect 124120 672320 124210 672560
rect 124450 672320 124540 672560
rect 124780 672320 124870 672560
rect 125110 672320 125220 672560
rect 125460 672320 125550 672560
rect 125790 672320 125880 672560
rect 126120 672320 126210 672560
rect 126450 672320 126560 672560
rect 126800 672320 126890 672560
rect 127130 672320 127220 672560
rect 127460 672320 127550 672560
rect 127790 672320 127900 672560
rect 128140 672320 128230 672560
rect 128470 672320 128560 672560
rect 128800 672320 128890 672560
rect 129130 672320 129240 672560
rect 129480 672320 129570 672560
rect 129810 672320 129900 672560
rect 130140 672320 130230 672560
rect 130470 672320 130580 672560
rect 130820 672320 130910 672560
rect 131150 672320 131240 672560
rect 131480 672320 131570 672560
rect 131810 672320 131920 672560
rect 132160 672320 132250 672560
rect 132490 672320 132580 672560
rect 132820 672320 132910 672560
rect 133150 672320 133170 672560
rect 122170 672300 133170 672320
rect 133550 683280 144550 683300
rect 133550 683040 133570 683280
rect 133810 683040 133920 683280
rect 134160 683040 134250 683280
rect 134490 683040 134580 683280
rect 134820 683040 134910 683280
rect 135150 683040 135260 683280
rect 135500 683040 135590 683280
rect 135830 683040 135920 683280
rect 136160 683040 136250 683280
rect 136490 683040 136600 683280
rect 136840 683040 136930 683280
rect 137170 683040 137260 683280
rect 137500 683040 137590 683280
rect 137830 683040 137940 683280
rect 138180 683040 138270 683280
rect 138510 683040 138600 683280
rect 138840 683040 138930 683280
rect 139170 683040 139280 683280
rect 139520 683040 139610 683280
rect 139850 683040 139940 683280
rect 140180 683040 140270 683280
rect 140510 683040 140620 683280
rect 140860 683040 140950 683280
rect 141190 683040 141280 683280
rect 141520 683040 141610 683280
rect 141850 683040 141960 683280
rect 142200 683040 142290 683280
rect 142530 683040 142620 683280
rect 142860 683040 142950 683280
rect 143190 683040 143300 683280
rect 143540 683040 143630 683280
rect 143870 683040 143960 683280
rect 144200 683040 144290 683280
rect 144530 683040 144550 683280
rect 133550 682950 144550 683040
rect 133550 682710 133570 682950
rect 133810 682710 133920 682950
rect 134160 682710 134250 682950
rect 134490 682710 134580 682950
rect 134820 682710 134910 682950
rect 135150 682710 135260 682950
rect 135500 682710 135590 682950
rect 135830 682710 135920 682950
rect 136160 682710 136250 682950
rect 136490 682710 136600 682950
rect 136840 682710 136930 682950
rect 137170 682710 137260 682950
rect 137500 682710 137590 682950
rect 137830 682710 137940 682950
rect 138180 682710 138270 682950
rect 138510 682710 138600 682950
rect 138840 682710 138930 682950
rect 139170 682710 139280 682950
rect 139520 682710 139610 682950
rect 139850 682710 139940 682950
rect 140180 682710 140270 682950
rect 140510 682710 140620 682950
rect 140860 682710 140950 682950
rect 141190 682710 141280 682950
rect 141520 682710 141610 682950
rect 141850 682710 141960 682950
rect 142200 682710 142290 682950
rect 142530 682710 142620 682950
rect 142860 682710 142950 682950
rect 143190 682710 143300 682950
rect 143540 682710 143630 682950
rect 143870 682710 143960 682950
rect 144200 682710 144290 682950
rect 144530 682710 144550 682950
rect 133550 682620 144550 682710
rect 133550 682380 133570 682620
rect 133810 682380 133920 682620
rect 134160 682380 134250 682620
rect 134490 682380 134580 682620
rect 134820 682380 134910 682620
rect 135150 682380 135260 682620
rect 135500 682380 135590 682620
rect 135830 682380 135920 682620
rect 136160 682380 136250 682620
rect 136490 682380 136600 682620
rect 136840 682380 136930 682620
rect 137170 682380 137260 682620
rect 137500 682380 137590 682620
rect 137830 682380 137940 682620
rect 138180 682380 138270 682620
rect 138510 682380 138600 682620
rect 138840 682380 138930 682620
rect 139170 682380 139280 682620
rect 139520 682380 139610 682620
rect 139850 682380 139940 682620
rect 140180 682380 140270 682620
rect 140510 682380 140620 682620
rect 140860 682380 140950 682620
rect 141190 682380 141280 682620
rect 141520 682380 141610 682620
rect 141850 682380 141960 682620
rect 142200 682380 142290 682620
rect 142530 682380 142620 682620
rect 142860 682380 142950 682620
rect 143190 682380 143300 682620
rect 143540 682380 143630 682620
rect 143870 682380 143960 682620
rect 144200 682380 144290 682620
rect 144530 682380 144550 682620
rect 133550 682290 144550 682380
rect 133550 682050 133570 682290
rect 133810 682050 133920 682290
rect 134160 682050 134250 682290
rect 134490 682050 134580 682290
rect 134820 682050 134910 682290
rect 135150 682050 135260 682290
rect 135500 682050 135590 682290
rect 135830 682050 135920 682290
rect 136160 682050 136250 682290
rect 136490 682050 136600 682290
rect 136840 682050 136930 682290
rect 137170 682050 137260 682290
rect 137500 682050 137590 682290
rect 137830 682050 137940 682290
rect 138180 682050 138270 682290
rect 138510 682050 138600 682290
rect 138840 682050 138930 682290
rect 139170 682050 139280 682290
rect 139520 682050 139610 682290
rect 139850 682050 139940 682290
rect 140180 682050 140270 682290
rect 140510 682050 140620 682290
rect 140860 682050 140950 682290
rect 141190 682050 141280 682290
rect 141520 682050 141610 682290
rect 141850 682050 141960 682290
rect 142200 682050 142290 682290
rect 142530 682050 142620 682290
rect 142860 682050 142950 682290
rect 143190 682050 143300 682290
rect 143540 682050 143630 682290
rect 143870 682050 143960 682290
rect 144200 682050 144290 682290
rect 144530 682050 144550 682290
rect 133550 681940 144550 682050
rect 133550 681700 133570 681940
rect 133810 681700 133920 681940
rect 134160 681700 134250 681940
rect 134490 681700 134580 681940
rect 134820 681700 134910 681940
rect 135150 681700 135260 681940
rect 135500 681700 135590 681940
rect 135830 681700 135920 681940
rect 136160 681700 136250 681940
rect 136490 681700 136600 681940
rect 136840 681700 136930 681940
rect 137170 681700 137260 681940
rect 137500 681700 137590 681940
rect 137830 681700 137940 681940
rect 138180 681700 138270 681940
rect 138510 681700 138600 681940
rect 138840 681700 138930 681940
rect 139170 681700 139280 681940
rect 139520 681700 139610 681940
rect 139850 681700 139940 681940
rect 140180 681700 140270 681940
rect 140510 681700 140620 681940
rect 140860 681700 140950 681940
rect 141190 681700 141280 681940
rect 141520 681700 141610 681940
rect 141850 681700 141960 681940
rect 142200 681700 142290 681940
rect 142530 681700 142620 681940
rect 142860 681700 142950 681940
rect 143190 681700 143300 681940
rect 143540 681700 143630 681940
rect 143870 681700 143960 681940
rect 144200 681700 144290 681940
rect 144530 681700 144550 681940
rect 133550 681610 144550 681700
rect 133550 681370 133570 681610
rect 133810 681370 133920 681610
rect 134160 681370 134250 681610
rect 134490 681370 134580 681610
rect 134820 681370 134910 681610
rect 135150 681370 135260 681610
rect 135500 681370 135590 681610
rect 135830 681370 135920 681610
rect 136160 681370 136250 681610
rect 136490 681370 136600 681610
rect 136840 681370 136930 681610
rect 137170 681370 137260 681610
rect 137500 681370 137590 681610
rect 137830 681370 137940 681610
rect 138180 681370 138270 681610
rect 138510 681370 138600 681610
rect 138840 681370 138930 681610
rect 139170 681370 139280 681610
rect 139520 681370 139610 681610
rect 139850 681370 139940 681610
rect 140180 681370 140270 681610
rect 140510 681370 140620 681610
rect 140860 681370 140950 681610
rect 141190 681370 141280 681610
rect 141520 681370 141610 681610
rect 141850 681370 141960 681610
rect 142200 681370 142290 681610
rect 142530 681370 142620 681610
rect 142860 681370 142950 681610
rect 143190 681370 143300 681610
rect 143540 681370 143630 681610
rect 143870 681370 143960 681610
rect 144200 681370 144290 681610
rect 144530 681370 144550 681610
rect 133550 681280 144550 681370
rect 133550 681040 133570 681280
rect 133810 681040 133920 681280
rect 134160 681040 134250 681280
rect 134490 681040 134580 681280
rect 134820 681040 134910 681280
rect 135150 681040 135260 681280
rect 135500 681040 135590 681280
rect 135830 681040 135920 681280
rect 136160 681040 136250 681280
rect 136490 681040 136600 681280
rect 136840 681040 136930 681280
rect 137170 681040 137260 681280
rect 137500 681040 137590 681280
rect 137830 681040 137940 681280
rect 138180 681040 138270 681280
rect 138510 681040 138600 681280
rect 138840 681040 138930 681280
rect 139170 681040 139280 681280
rect 139520 681040 139610 681280
rect 139850 681040 139940 681280
rect 140180 681040 140270 681280
rect 140510 681040 140620 681280
rect 140860 681040 140950 681280
rect 141190 681040 141280 681280
rect 141520 681040 141610 681280
rect 141850 681040 141960 681280
rect 142200 681040 142290 681280
rect 142530 681040 142620 681280
rect 142860 681040 142950 681280
rect 143190 681040 143300 681280
rect 143540 681040 143630 681280
rect 143870 681040 143960 681280
rect 144200 681040 144290 681280
rect 144530 681040 144550 681280
rect 133550 680950 144550 681040
rect 133550 680710 133570 680950
rect 133810 680710 133920 680950
rect 134160 680710 134250 680950
rect 134490 680710 134580 680950
rect 134820 680710 134910 680950
rect 135150 680710 135260 680950
rect 135500 680710 135590 680950
rect 135830 680710 135920 680950
rect 136160 680710 136250 680950
rect 136490 680710 136600 680950
rect 136840 680710 136930 680950
rect 137170 680710 137260 680950
rect 137500 680710 137590 680950
rect 137830 680710 137940 680950
rect 138180 680710 138270 680950
rect 138510 680710 138600 680950
rect 138840 680710 138930 680950
rect 139170 680710 139280 680950
rect 139520 680710 139610 680950
rect 139850 680710 139940 680950
rect 140180 680710 140270 680950
rect 140510 680710 140620 680950
rect 140860 680710 140950 680950
rect 141190 680710 141280 680950
rect 141520 680710 141610 680950
rect 141850 680710 141960 680950
rect 142200 680710 142290 680950
rect 142530 680710 142620 680950
rect 142860 680710 142950 680950
rect 143190 680710 143300 680950
rect 143540 680710 143630 680950
rect 143870 680710 143960 680950
rect 144200 680710 144290 680950
rect 144530 680710 144550 680950
rect 133550 680600 144550 680710
rect 133550 680360 133570 680600
rect 133810 680360 133920 680600
rect 134160 680360 134250 680600
rect 134490 680360 134580 680600
rect 134820 680360 134910 680600
rect 135150 680360 135260 680600
rect 135500 680360 135590 680600
rect 135830 680360 135920 680600
rect 136160 680360 136250 680600
rect 136490 680360 136600 680600
rect 136840 680360 136930 680600
rect 137170 680360 137260 680600
rect 137500 680360 137590 680600
rect 137830 680360 137940 680600
rect 138180 680360 138270 680600
rect 138510 680360 138600 680600
rect 138840 680360 138930 680600
rect 139170 680360 139280 680600
rect 139520 680360 139610 680600
rect 139850 680360 139940 680600
rect 140180 680360 140270 680600
rect 140510 680360 140620 680600
rect 140860 680360 140950 680600
rect 141190 680360 141280 680600
rect 141520 680360 141610 680600
rect 141850 680360 141960 680600
rect 142200 680360 142290 680600
rect 142530 680360 142620 680600
rect 142860 680360 142950 680600
rect 143190 680360 143300 680600
rect 143540 680360 143630 680600
rect 143870 680360 143960 680600
rect 144200 680360 144290 680600
rect 144530 680360 144550 680600
rect 133550 680270 144550 680360
rect 133550 680030 133570 680270
rect 133810 680030 133920 680270
rect 134160 680030 134250 680270
rect 134490 680030 134580 680270
rect 134820 680030 134910 680270
rect 135150 680030 135260 680270
rect 135500 680030 135590 680270
rect 135830 680030 135920 680270
rect 136160 680030 136250 680270
rect 136490 680030 136600 680270
rect 136840 680030 136930 680270
rect 137170 680030 137260 680270
rect 137500 680030 137590 680270
rect 137830 680030 137940 680270
rect 138180 680030 138270 680270
rect 138510 680030 138600 680270
rect 138840 680030 138930 680270
rect 139170 680030 139280 680270
rect 139520 680030 139610 680270
rect 139850 680030 139940 680270
rect 140180 680030 140270 680270
rect 140510 680030 140620 680270
rect 140860 680030 140950 680270
rect 141190 680030 141280 680270
rect 141520 680030 141610 680270
rect 141850 680030 141960 680270
rect 142200 680030 142290 680270
rect 142530 680030 142620 680270
rect 142860 680030 142950 680270
rect 143190 680030 143300 680270
rect 143540 680030 143630 680270
rect 143870 680030 143960 680270
rect 144200 680030 144290 680270
rect 144530 680030 144550 680270
rect 133550 679940 144550 680030
rect 133550 679700 133570 679940
rect 133810 679700 133920 679940
rect 134160 679700 134250 679940
rect 134490 679700 134580 679940
rect 134820 679700 134910 679940
rect 135150 679700 135260 679940
rect 135500 679700 135590 679940
rect 135830 679700 135920 679940
rect 136160 679700 136250 679940
rect 136490 679700 136600 679940
rect 136840 679700 136930 679940
rect 137170 679700 137260 679940
rect 137500 679700 137590 679940
rect 137830 679700 137940 679940
rect 138180 679700 138270 679940
rect 138510 679700 138600 679940
rect 138840 679700 138930 679940
rect 139170 679700 139280 679940
rect 139520 679700 139610 679940
rect 139850 679700 139940 679940
rect 140180 679700 140270 679940
rect 140510 679700 140620 679940
rect 140860 679700 140950 679940
rect 141190 679700 141280 679940
rect 141520 679700 141610 679940
rect 141850 679700 141960 679940
rect 142200 679700 142290 679940
rect 142530 679700 142620 679940
rect 142860 679700 142950 679940
rect 143190 679700 143300 679940
rect 143540 679700 143630 679940
rect 143870 679700 143960 679940
rect 144200 679700 144290 679940
rect 144530 679700 144550 679940
rect 133550 679610 144550 679700
rect 133550 679370 133570 679610
rect 133810 679370 133920 679610
rect 134160 679370 134250 679610
rect 134490 679370 134580 679610
rect 134820 679370 134910 679610
rect 135150 679370 135260 679610
rect 135500 679370 135590 679610
rect 135830 679370 135920 679610
rect 136160 679370 136250 679610
rect 136490 679370 136600 679610
rect 136840 679370 136930 679610
rect 137170 679370 137260 679610
rect 137500 679370 137590 679610
rect 137830 679370 137940 679610
rect 138180 679370 138270 679610
rect 138510 679370 138600 679610
rect 138840 679370 138930 679610
rect 139170 679370 139280 679610
rect 139520 679370 139610 679610
rect 139850 679370 139940 679610
rect 140180 679370 140270 679610
rect 140510 679370 140620 679610
rect 140860 679370 140950 679610
rect 141190 679370 141280 679610
rect 141520 679370 141610 679610
rect 141850 679370 141960 679610
rect 142200 679370 142290 679610
rect 142530 679370 142620 679610
rect 142860 679370 142950 679610
rect 143190 679370 143300 679610
rect 143540 679370 143630 679610
rect 143870 679370 143960 679610
rect 144200 679370 144290 679610
rect 144530 679370 144550 679610
rect 133550 679260 144550 679370
rect 133550 679020 133570 679260
rect 133810 679020 133920 679260
rect 134160 679020 134250 679260
rect 134490 679020 134580 679260
rect 134820 679020 134910 679260
rect 135150 679020 135260 679260
rect 135500 679020 135590 679260
rect 135830 679020 135920 679260
rect 136160 679020 136250 679260
rect 136490 679020 136600 679260
rect 136840 679020 136930 679260
rect 137170 679020 137260 679260
rect 137500 679020 137590 679260
rect 137830 679020 137940 679260
rect 138180 679020 138270 679260
rect 138510 679020 138600 679260
rect 138840 679020 138930 679260
rect 139170 679020 139280 679260
rect 139520 679020 139610 679260
rect 139850 679020 139940 679260
rect 140180 679020 140270 679260
rect 140510 679020 140620 679260
rect 140860 679020 140950 679260
rect 141190 679020 141280 679260
rect 141520 679020 141610 679260
rect 141850 679020 141960 679260
rect 142200 679020 142290 679260
rect 142530 679020 142620 679260
rect 142860 679020 142950 679260
rect 143190 679020 143300 679260
rect 143540 679020 143630 679260
rect 143870 679020 143960 679260
rect 144200 679020 144290 679260
rect 144530 679020 144550 679260
rect 133550 678930 144550 679020
rect 133550 678690 133570 678930
rect 133810 678690 133920 678930
rect 134160 678690 134250 678930
rect 134490 678690 134580 678930
rect 134820 678690 134910 678930
rect 135150 678690 135260 678930
rect 135500 678690 135590 678930
rect 135830 678690 135920 678930
rect 136160 678690 136250 678930
rect 136490 678690 136600 678930
rect 136840 678690 136930 678930
rect 137170 678690 137260 678930
rect 137500 678690 137590 678930
rect 137830 678690 137940 678930
rect 138180 678690 138270 678930
rect 138510 678690 138600 678930
rect 138840 678690 138930 678930
rect 139170 678690 139280 678930
rect 139520 678690 139610 678930
rect 139850 678690 139940 678930
rect 140180 678690 140270 678930
rect 140510 678690 140620 678930
rect 140860 678690 140950 678930
rect 141190 678690 141280 678930
rect 141520 678690 141610 678930
rect 141850 678690 141960 678930
rect 142200 678690 142290 678930
rect 142530 678690 142620 678930
rect 142860 678690 142950 678930
rect 143190 678690 143300 678930
rect 143540 678690 143630 678930
rect 143870 678690 143960 678930
rect 144200 678690 144290 678930
rect 144530 678690 144550 678930
rect 133550 678600 144550 678690
rect 133550 678360 133570 678600
rect 133810 678360 133920 678600
rect 134160 678360 134250 678600
rect 134490 678360 134580 678600
rect 134820 678360 134910 678600
rect 135150 678360 135260 678600
rect 135500 678360 135590 678600
rect 135830 678360 135920 678600
rect 136160 678360 136250 678600
rect 136490 678360 136600 678600
rect 136840 678360 136930 678600
rect 137170 678360 137260 678600
rect 137500 678360 137590 678600
rect 137830 678360 137940 678600
rect 138180 678360 138270 678600
rect 138510 678360 138600 678600
rect 138840 678360 138930 678600
rect 139170 678360 139280 678600
rect 139520 678360 139610 678600
rect 139850 678360 139940 678600
rect 140180 678360 140270 678600
rect 140510 678360 140620 678600
rect 140860 678360 140950 678600
rect 141190 678360 141280 678600
rect 141520 678360 141610 678600
rect 141850 678360 141960 678600
rect 142200 678360 142290 678600
rect 142530 678360 142620 678600
rect 142860 678360 142950 678600
rect 143190 678360 143300 678600
rect 143540 678360 143630 678600
rect 143870 678360 143960 678600
rect 144200 678360 144290 678600
rect 144530 678360 144550 678600
rect 133550 678270 144550 678360
rect 133550 678030 133570 678270
rect 133810 678030 133920 678270
rect 134160 678030 134250 678270
rect 134490 678030 134580 678270
rect 134820 678030 134910 678270
rect 135150 678030 135260 678270
rect 135500 678030 135590 678270
rect 135830 678030 135920 678270
rect 136160 678030 136250 678270
rect 136490 678030 136600 678270
rect 136840 678030 136930 678270
rect 137170 678030 137260 678270
rect 137500 678030 137590 678270
rect 137830 678030 137940 678270
rect 138180 678030 138270 678270
rect 138510 678030 138600 678270
rect 138840 678030 138930 678270
rect 139170 678030 139280 678270
rect 139520 678030 139610 678270
rect 139850 678030 139940 678270
rect 140180 678030 140270 678270
rect 140510 678030 140620 678270
rect 140860 678030 140950 678270
rect 141190 678030 141280 678270
rect 141520 678030 141610 678270
rect 141850 678030 141960 678270
rect 142200 678030 142290 678270
rect 142530 678030 142620 678270
rect 142860 678030 142950 678270
rect 143190 678030 143300 678270
rect 143540 678030 143630 678270
rect 143870 678030 143960 678270
rect 144200 678030 144290 678270
rect 144530 678030 144550 678270
rect 133550 677920 144550 678030
rect 133550 677680 133570 677920
rect 133810 677680 133920 677920
rect 134160 677680 134250 677920
rect 134490 677680 134580 677920
rect 134820 677680 134910 677920
rect 135150 677680 135260 677920
rect 135500 677680 135590 677920
rect 135830 677680 135920 677920
rect 136160 677680 136250 677920
rect 136490 677680 136600 677920
rect 136840 677680 136930 677920
rect 137170 677680 137260 677920
rect 137500 677680 137590 677920
rect 137830 677680 137940 677920
rect 138180 677680 138270 677920
rect 138510 677680 138600 677920
rect 138840 677680 138930 677920
rect 139170 677680 139280 677920
rect 139520 677680 139610 677920
rect 139850 677680 139940 677920
rect 140180 677680 140270 677920
rect 140510 677680 140620 677920
rect 140860 677680 140950 677920
rect 141190 677680 141280 677920
rect 141520 677680 141610 677920
rect 141850 677680 141960 677920
rect 142200 677680 142290 677920
rect 142530 677680 142620 677920
rect 142860 677680 142950 677920
rect 143190 677680 143300 677920
rect 143540 677680 143630 677920
rect 143870 677680 143960 677920
rect 144200 677680 144290 677920
rect 144530 677680 144550 677920
rect 133550 677590 144550 677680
rect 133550 677350 133570 677590
rect 133810 677350 133920 677590
rect 134160 677350 134250 677590
rect 134490 677350 134580 677590
rect 134820 677350 134910 677590
rect 135150 677350 135260 677590
rect 135500 677350 135590 677590
rect 135830 677350 135920 677590
rect 136160 677350 136250 677590
rect 136490 677350 136600 677590
rect 136840 677350 136930 677590
rect 137170 677350 137260 677590
rect 137500 677350 137590 677590
rect 137830 677350 137940 677590
rect 138180 677350 138270 677590
rect 138510 677350 138600 677590
rect 138840 677350 138930 677590
rect 139170 677350 139280 677590
rect 139520 677350 139610 677590
rect 139850 677350 139940 677590
rect 140180 677350 140270 677590
rect 140510 677350 140620 677590
rect 140860 677350 140950 677590
rect 141190 677350 141280 677590
rect 141520 677350 141610 677590
rect 141850 677350 141960 677590
rect 142200 677350 142290 677590
rect 142530 677350 142620 677590
rect 142860 677350 142950 677590
rect 143190 677350 143300 677590
rect 143540 677350 143630 677590
rect 143870 677350 143960 677590
rect 144200 677350 144290 677590
rect 144530 677350 144550 677590
rect 133550 677260 144550 677350
rect 133550 677020 133570 677260
rect 133810 677020 133920 677260
rect 134160 677020 134250 677260
rect 134490 677020 134580 677260
rect 134820 677020 134910 677260
rect 135150 677020 135260 677260
rect 135500 677020 135590 677260
rect 135830 677020 135920 677260
rect 136160 677020 136250 677260
rect 136490 677020 136600 677260
rect 136840 677020 136930 677260
rect 137170 677020 137260 677260
rect 137500 677020 137590 677260
rect 137830 677020 137940 677260
rect 138180 677020 138270 677260
rect 138510 677020 138600 677260
rect 138840 677020 138930 677260
rect 139170 677020 139280 677260
rect 139520 677020 139610 677260
rect 139850 677020 139940 677260
rect 140180 677020 140270 677260
rect 140510 677020 140620 677260
rect 140860 677020 140950 677260
rect 141190 677020 141280 677260
rect 141520 677020 141610 677260
rect 141850 677020 141960 677260
rect 142200 677020 142290 677260
rect 142530 677020 142620 677260
rect 142860 677020 142950 677260
rect 143190 677020 143300 677260
rect 143540 677020 143630 677260
rect 143870 677020 143960 677260
rect 144200 677020 144290 677260
rect 144530 677020 144550 677260
rect 133550 676930 144550 677020
rect 133550 676690 133570 676930
rect 133810 676690 133920 676930
rect 134160 676690 134250 676930
rect 134490 676690 134580 676930
rect 134820 676690 134910 676930
rect 135150 676690 135260 676930
rect 135500 676690 135590 676930
rect 135830 676690 135920 676930
rect 136160 676690 136250 676930
rect 136490 676690 136600 676930
rect 136840 676690 136930 676930
rect 137170 676690 137260 676930
rect 137500 676690 137590 676930
rect 137830 676690 137940 676930
rect 138180 676690 138270 676930
rect 138510 676690 138600 676930
rect 138840 676690 138930 676930
rect 139170 676690 139280 676930
rect 139520 676690 139610 676930
rect 139850 676690 139940 676930
rect 140180 676690 140270 676930
rect 140510 676690 140620 676930
rect 140860 676690 140950 676930
rect 141190 676690 141280 676930
rect 141520 676690 141610 676930
rect 141850 676690 141960 676930
rect 142200 676690 142290 676930
rect 142530 676690 142620 676930
rect 142860 676690 142950 676930
rect 143190 676690 143300 676930
rect 143540 676690 143630 676930
rect 143870 676690 143960 676930
rect 144200 676690 144290 676930
rect 144530 676690 144550 676930
rect 133550 676580 144550 676690
rect 133550 676340 133570 676580
rect 133810 676340 133920 676580
rect 134160 676340 134250 676580
rect 134490 676340 134580 676580
rect 134820 676340 134910 676580
rect 135150 676340 135260 676580
rect 135500 676340 135590 676580
rect 135830 676340 135920 676580
rect 136160 676340 136250 676580
rect 136490 676340 136600 676580
rect 136840 676340 136930 676580
rect 137170 676340 137260 676580
rect 137500 676340 137590 676580
rect 137830 676340 137940 676580
rect 138180 676340 138270 676580
rect 138510 676340 138600 676580
rect 138840 676340 138930 676580
rect 139170 676340 139280 676580
rect 139520 676340 139610 676580
rect 139850 676340 139940 676580
rect 140180 676340 140270 676580
rect 140510 676340 140620 676580
rect 140860 676340 140950 676580
rect 141190 676340 141280 676580
rect 141520 676340 141610 676580
rect 141850 676340 141960 676580
rect 142200 676340 142290 676580
rect 142530 676340 142620 676580
rect 142860 676340 142950 676580
rect 143190 676340 143300 676580
rect 143540 676340 143630 676580
rect 143870 676340 143960 676580
rect 144200 676340 144290 676580
rect 144530 676340 144550 676580
rect 133550 676250 144550 676340
rect 133550 676010 133570 676250
rect 133810 676010 133920 676250
rect 134160 676010 134250 676250
rect 134490 676010 134580 676250
rect 134820 676010 134910 676250
rect 135150 676010 135260 676250
rect 135500 676010 135590 676250
rect 135830 676010 135920 676250
rect 136160 676010 136250 676250
rect 136490 676010 136600 676250
rect 136840 676010 136930 676250
rect 137170 676010 137260 676250
rect 137500 676010 137590 676250
rect 137830 676010 137940 676250
rect 138180 676010 138270 676250
rect 138510 676010 138600 676250
rect 138840 676010 138930 676250
rect 139170 676010 139280 676250
rect 139520 676010 139610 676250
rect 139850 676010 139940 676250
rect 140180 676010 140270 676250
rect 140510 676010 140620 676250
rect 140860 676010 140950 676250
rect 141190 676010 141280 676250
rect 141520 676010 141610 676250
rect 141850 676010 141960 676250
rect 142200 676010 142290 676250
rect 142530 676010 142620 676250
rect 142860 676010 142950 676250
rect 143190 676010 143300 676250
rect 143540 676010 143630 676250
rect 143870 676010 143960 676250
rect 144200 676010 144290 676250
rect 144530 676010 144550 676250
rect 133550 675920 144550 676010
rect 133550 675680 133570 675920
rect 133810 675680 133920 675920
rect 134160 675680 134250 675920
rect 134490 675680 134580 675920
rect 134820 675680 134910 675920
rect 135150 675680 135260 675920
rect 135500 675680 135590 675920
rect 135830 675680 135920 675920
rect 136160 675680 136250 675920
rect 136490 675680 136600 675920
rect 136840 675680 136930 675920
rect 137170 675680 137260 675920
rect 137500 675680 137590 675920
rect 137830 675680 137940 675920
rect 138180 675680 138270 675920
rect 138510 675680 138600 675920
rect 138840 675680 138930 675920
rect 139170 675680 139280 675920
rect 139520 675680 139610 675920
rect 139850 675680 139940 675920
rect 140180 675680 140270 675920
rect 140510 675680 140620 675920
rect 140860 675680 140950 675920
rect 141190 675680 141280 675920
rect 141520 675680 141610 675920
rect 141850 675680 141960 675920
rect 142200 675680 142290 675920
rect 142530 675680 142620 675920
rect 142860 675680 142950 675920
rect 143190 675680 143300 675920
rect 143540 675680 143630 675920
rect 143870 675680 143960 675920
rect 144200 675680 144290 675920
rect 144530 675680 144550 675920
rect 133550 675590 144550 675680
rect 133550 675350 133570 675590
rect 133810 675350 133920 675590
rect 134160 675350 134250 675590
rect 134490 675350 134580 675590
rect 134820 675350 134910 675590
rect 135150 675350 135260 675590
rect 135500 675350 135590 675590
rect 135830 675350 135920 675590
rect 136160 675350 136250 675590
rect 136490 675350 136600 675590
rect 136840 675350 136930 675590
rect 137170 675350 137260 675590
rect 137500 675350 137590 675590
rect 137830 675350 137940 675590
rect 138180 675350 138270 675590
rect 138510 675350 138600 675590
rect 138840 675350 138930 675590
rect 139170 675350 139280 675590
rect 139520 675350 139610 675590
rect 139850 675350 139940 675590
rect 140180 675350 140270 675590
rect 140510 675350 140620 675590
rect 140860 675350 140950 675590
rect 141190 675350 141280 675590
rect 141520 675350 141610 675590
rect 141850 675350 141960 675590
rect 142200 675350 142290 675590
rect 142530 675350 142620 675590
rect 142860 675350 142950 675590
rect 143190 675350 143300 675590
rect 143540 675350 143630 675590
rect 143870 675350 143960 675590
rect 144200 675350 144290 675590
rect 144530 675350 144550 675590
rect 133550 675240 144550 675350
rect 133550 675000 133570 675240
rect 133810 675000 133920 675240
rect 134160 675000 134250 675240
rect 134490 675000 134580 675240
rect 134820 675000 134910 675240
rect 135150 675000 135260 675240
rect 135500 675000 135590 675240
rect 135830 675000 135920 675240
rect 136160 675000 136250 675240
rect 136490 675000 136600 675240
rect 136840 675000 136930 675240
rect 137170 675000 137260 675240
rect 137500 675000 137590 675240
rect 137830 675000 137940 675240
rect 138180 675000 138270 675240
rect 138510 675000 138600 675240
rect 138840 675000 138930 675240
rect 139170 675000 139280 675240
rect 139520 675000 139610 675240
rect 139850 675000 139940 675240
rect 140180 675000 140270 675240
rect 140510 675000 140620 675240
rect 140860 675000 140950 675240
rect 141190 675000 141280 675240
rect 141520 675000 141610 675240
rect 141850 675000 141960 675240
rect 142200 675000 142290 675240
rect 142530 675000 142620 675240
rect 142860 675000 142950 675240
rect 143190 675000 143300 675240
rect 143540 675000 143630 675240
rect 143870 675000 143960 675240
rect 144200 675000 144290 675240
rect 144530 675000 144550 675240
rect 133550 674910 144550 675000
rect 133550 674670 133570 674910
rect 133810 674670 133920 674910
rect 134160 674670 134250 674910
rect 134490 674670 134580 674910
rect 134820 674670 134910 674910
rect 135150 674670 135260 674910
rect 135500 674670 135590 674910
rect 135830 674670 135920 674910
rect 136160 674670 136250 674910
rect 136490 674670 136600 674910
rect 136840 674670 136930 674910
rect 137170 674670 137260 674910
rect 137500 674670 137590 674910
rect 137830 674670 137940 674910
rect 138180 674670 138270 674910
rect 138510 674670 138600 674910
rect 138840 674670 138930 674910
rect 139170 674670 139280 674910
rect 139520 674670 139610 674910
rect 139850 674670 139940 674910
rect 140180 674670 140270 674910
rect 140510 674670 140620 674910
rect 140860 674670 140950 674910
rect 141190 674670 141280 674910
rect 141520 674670 141610 674910
rect 141850 674670 141960 674910
rect 142200 674670 142290 674910
rect 142530 674670 142620 674910
rect 142860 674670 142950 674910
rect 143190 674670 143300 674910
rect 143540 674670 143630 674910
rect 143870 674670 143960 674910
rect 144200 674670 144290 674910
rect 144530 674670 144550 674910
rect 133550 674580 144550 674670
rect 133550 674340 133570 674580
rect 133810 674340 133920 674580
rect 134160 674340 134250 674580
rect 134490 674340 134580 674580
rect 134820 674340 134910 674580
rect 135150 674340 135260 674580
rect 135500 674340 135590 674580
rect 135830 674340 135920 674580
rect 136160 674340 136250 674580
rect 136490 674340 136600 674580
rect 136840 674340 136930 674580
rect 137170 674340 137260 674580
rect 137500 674340 137590 674580
rect 137830 674340 137940 674580
rect 138180 674340 138270 674580
rect 138510 674340 138600 674580
rect 138840 674340 138930 674580
rect 139170 674340 139280 674580
rect 139520 674340 139610 674580
rect 139850 674340 139940 674580
rect 140180 674340 140270 674580
rect 140510 674340 140620 674580
rect 140860 674340 140950 674580
rect 141190 674340 141280 674580
rect 141520 674340 141610 674580
rect 141850 674340 141960 674580
rect 142200 674340 142290 674580
rect 142530 674340 142620 674580
rect 142860 674340 142950 674580
rect 143190 674340 143300 674580
rect 143540 674340 143630 674580
rect 143870 674340 143960 674580
rect 144200 674340 144290 674580
rect 144530 674340 144550 674580
rect 133550 674250 144550 674340
rect 133550 674010 133570 674250
rect 133810 674010 133920 674250
rect 134160 674010 134250 674250
rect 134490 674010 134580 674250
rect 134820 674010 134910 674250
rect 135150 674010 135260 674250
rect 135500 674010 135590 674250
rect 135830 674010 135920 674250
rect 136160 674010 136250 674250
rect 136490 674010 136600 674250
rect 136840 674010 136930 674250
rect 137170 674010 137260 674250
rect 137500 674010 137590 674250
rect 137830 674010 137940 674250
rect 138180 674010 138270 674250
rect 138510 674010 138600 674250
rect 138840 674010 138930 674250
rect 139170 674010 139280 674250
rect 139520 674010 139610 674250
rect 139850 674010 139940 674250
rect 140180 674010 140270 674250
rect 140510 674010 140620 674250
rect 140860 674010 140950 674250
rect 141190 674010 141280 674250
rect 141520 674010 141610 674250
rect 141850 674010 141960 674250
rect 142200 674010 142290 674250
rect 142530 674010 142620 674250
rect 142860 674010 142950 674250
rect 143190 674010 143300 674250
rect 143540 674010 143630 674250
rect 143870 674010 143960 674250
rect 144200 674010 144290 674250
rect 144530 674010 144550 674250
rect 133550 673900 144550 674010
rect 133550 673660 133570 673900
rect 133810 673660 133920 673900
rect 134160 673660 134250 673900
rect 134490 673660 134580 673900
rect 134820 673660 134910 673900
rect 135150 673660 135260 673900
rect 135500 673660 135590 673900
rect 135830 673660 135920 673900
rect 136160 673660 136250 673900
rect 136490 673660 136600 673900
rect 136840 673660 136930 673900
rect 137170 673660 137260 673900
rect 137500 673660 137590 673900
rect 137830 673660 137940 673900
rect 138180 673660 138270 673900
rect 138510 673660 138600 673900
rect 138840 673660 138930 673900
rect 139170 673660 139280 673900
rect 139520 673660 139610 673900
rect 139850 673660 139940 673900
rect 140180 673660 140270 673900
rect 140510 673660 140620 673900
rect 140860 673660 140950 673900
rect 141190 673660 141280 673900
rect 141520 673660 141610 673900
rect 141850 673660 141960 673900
rect 142200 673660 142290 673900
rect 142530 673660 142620 673900
rect 142860 673660 142950 673900
rect 143190 673660 143300 673900
rect 143540 673660 143630 673900
rect 143870 673660 143960 673900
rect 144200 673660 144290 673900
rect 144530 673660 144550 673900
rect 133550 673570 144550 673660
rect 133550 673330 133570 673570
rect 133810 673330 133920 673570
rect 134160 673330 134250 673570
rect 134490 673330 134580 673570
rect 134820 673330 134910 673570
rect 135150 673330 135260 673570
rect 135500 673330 135590 673570
rect 135830 673330 135920 673570
rect 136160 673330 136250 673570
rect 136490 673330 136600 673570
rect 136840 673330 136930 673570
rect 137170 673330 137260 673570
rect 137500 673330 137590 673570
rect 137830 673330 137940 673570
rect 138180 673330 138270 673570
rect 138510 673330 138600 673570
rect 138840 673330 138930 673570
rect 139170 673330 139280 673570
rect 139520 673330 139610 673570
rect 139850 673330 139940 673570
rect 140180 673330 140270 673570
rect 140510 673330 140620 673570
rect 140860 673330 140950 673570
rect 141190 673330 141280 673570
rect 141520 673330 141610 673570
rect 141850 673330 141960 673570
rect 142200 673330 142290 673570
rect 142530 673330 142620 673570
rect 142860 673330 142950 673570
rect 143190 673330 143300 673570
rect 143540 673330 143630 673570
rect 143870 673330 143960 673570
rect 144200 673330 144290 673570
rect 144530 673330 144550 673570
rect 133550 673240 144550 673330
rect 133550 673000 133570 673240
rect 133810 673000 133920 673240
rect 134160 673000 134250 673240
rect 134490 673000 134580 673240
rect 134820 673000 134910 673240
rect 135150 673000 135260 673240
rect 135500 673000 135590 673240
rect 135830 673000 135920 673240
rect 136160 673000 136250 673240
rect 136490 673000 136600 673240
rect 136840 673000 136930 673240
rect 137170 673000 137260 673240
rect 137500 673000 137590 673240
rect 137830 673000 137940 673240
rect 138180 673000 138270 673240
rect 138510 673000 138600 673240
rect 138840 673000 138930 673240
rect 139170 673000 139280 673240
rect 139520 673000 139610 673240
rect 139850 673000 139940 673240
rect 140180 673000 140270 673240
rect 140510 673000 140620 673240
rect 140860 673000 140950 673240
rect 141190 673000 141280 673240
rect 141520 673000 141610 673240
rect 141850 673000 141960 673240
rect 142200 673000 142290 673240
rect 142530 673000 142620 673240
rect 142860 673000 142950 673240
rect 143190 673000 143300 673240
rect 143540 673000 143630 673240
rect 143870 673000 143960 673240
rect 144200 673000 144290 673240
rect 144530 673000 144550 673240
rect 133550 672910 144550 673000
rect 133550 672670 133570 672910
rect 133810 672670 133920 672910
rect 134160 672670 134250 672910
rect 134490 672670 134580 672910
rect 134820 672670 134910 672910
rect 135150 672670 135260 672910
rect 135500 672670 135590 672910
rect 135830 672670 135920 672910
rect 136160 672670 136250 672910
rect 136490 672670 136600 672910
rect 136840 672670 136930 672910
rect 137170 672670 137260 672910
rect 137500 672670 137590 672910
rect 137830 672670 137940 672910
rect 138180 672670 138270 672910
rect 138510 672670 138600 672910
rect 138840 672670 138930 672910
rect 139170 672670 139280 672910
rect 139520 672670 139610 672910
rect 139850 672670 139940 672910
rect 140180 672670 140270 672910
rect 140510 672670 140620 672910
rect 140860 672670 140950 672910
rect 141190 672670 141280 672910
rect 141520 672670 141610 672910
rect 141850 672670 141960 672910
rect 142200 672670 142290 672910
rect 142530 672670 142620 672910
rect 142860 672670 142950 672910
rect 143190 672670 143300 672910
rect 143540 672670 143630 672910
rect 143870 672670 143960 672910
rect 144200 672670 144290 672910
rect 144530 672670 144550 672910
rect 133550 672560 144550 672670
rect 133550 672320 133570 672560
rect 133810 672320 133920 672560
rect 134160 672320 134250 672560
rect 134490 672320 134580 672560
rect 134820 672320 134910 672560
rect 135150 672320 135260 672560
rect 135500 672320 135590 672560
rect 135830 672320 135920 672560
rect 136160 672320 136250 672560
rect 136490 672320 136600 672560
rect 136840 672320 136930 672560
rect 137170 672320 137260 672560
rect 137500 672320 137590 672560
rect 137830 672320 137940 672560
rect 138180 672320 138270 672560
rect 138510 672320 138600 672560
rect 138840 672320 138930 672560
rect 139170 672320 139280 672560
rect 139520 672320 139610 672560
rect 139850 672320 139940 672560
rect 140180 672320 140270 672560
rect 140510 672320 140620 672560
rect 140860 672320 140950 672560
rect 141190 672320 141280 672560
rect 141520 672320 141610 672560
rect 141850 672320 141960 672560
rect 142200 672320 142290 672560
rect 142530 672320 142620 672560
rect 142860 672320 142950 672560
rect 143190 672320 143300 672560
rect 143540 672320 143630 672560
rect 143870 672320 143960 672560
rect 144200 672320 144290 672560
rect 144530 672320 144550 672560
rect 133550 672300 144550 672320
rect 144930 683280 155930 683300
rect 144930 683040 144950 683280
rect 145190 683040 145300 683280
rect 145540 683040 145630 683280
rect 145870 683040 145960 683280
rect 146200 683040 146290 683280
rect 146530 683040 146640 683280
rect 146880 683040 146970 683280
rect 147210 683040 147300 683280
rect 147540 683040 147630 683280
rect 147870 683040 147980 683280
rect 148220 683040 148310 683280
rect 148550 683040 148640 683280
rect 148880 683040 148970 683280
rect 149210 683040 149320 683280
rect 149560 683040 149650 683280
rect 149890 683040 149980 683280
rect 150220 683040 150310 683280
rect 150550 683040 150660 683280
rect 150900 683040 150990 683280
rect 151230 683040 151320 683280
rect 151560 683040 151650 683280
rect 151890 683040 152000 683280
rect 152240 683040 152330 683280
rect 152570 683040 152660 683280
rect 152900 683040 152990 683280
rect 153230 683040 153340 683280
rect 153580 683040 153670 683280
rect 153910 683040 154000 683280
rect 154240 683040 154330 683280
rect 154570 683040 154680 683280
rect 154920 683040 155010 683280
rect 155250 683040 155340 683280
rect 155580 683040 155670 683280
rect 155910 683040 155930 683280
rect 144930 682950 155930 683040
rect 144930 682710 144950 682950
rect 145190 682710 145300 682950
rect 145540 682710 145630 682950
rect 145870 682710 145960 682950
rect 146200 682710 146290 682950
rect 146530 682710 146640 682950
rect 146880 682710 146970 682950
rect 147210 682710 147300 682950
rect 147540 682710 147630 682950
rect 147870 682710 147980 682950
rect 148220 682710 148310 682950
rect 148550 682710 148640 682950
rect 148880 682710 148970 682950
rect 149210 682710 149320 682950
rect 149560 682710 149650 682950
rect 149890 682710 149980 682950
rect 150220 682710 150310 682950
rect 150550 682710 150660 682950
rect 150900 682710 150990 682950
rect 151230 682710 151320 682950
rect 151560 682710 151650 682950
rect 151890 682710 152000 682950
rect 152240 682710 152330 682950
rect 152570 682710 152660 682950
rect 152900 682710 152990 682950
rect 153230 682710 153340 682950
rect 153580 682710 153670 682950
rect 153910 682710 154000 682950
rect 154240 682710 154330 682950
rect 154570 682710 154680 682950
rect 154920 682710 155010 682950
rect 155250 682710 155340 682950
rect 155580 682710 155670 682950
rect 155910 682710 155930 682950
rect 144930 682620 155930 682710
rect 144930 682380 144950 682620
rect 145190 682380 145300 682620
rect 145540 682380 145630 682620
rect 145870 682380 145960 682620
rect 146200 682380 146290 682620
rect 146530 682380 146640 682620
rect 146880 682380 146970 682620
rect 147210 682380 147300 682620
rect 147540 682380 147630 682620
rect 147870 682380 147980 682620
rect 148220 682380 148310 682620
rect 148550 682380 148640 682620
rect 148880 682380 148970 682620
rect 149210 682380 149320 682620
rect 149560 682380 149650 682620
rect 149890 682380 149980 682620
rect 150220 682380 150310 682620
rect 150550 682380 150660 682620
rect 150900 682380 150990 682620
rect 151230 682380 151320 682620
rect 151560 682380 151650 682620
rect 151890 682380 152000 682620
rect 152240 682380 152330 682620
rect 152570 682380 152660 682620
rect 152900 682380 152990 682620
rect 153230 682380 153340 682620
rect 153580 682380 153670 682620
rect 153910 682380 154000 682620
rect 154240 682380 154330 682620
rect 154570 682380 154680 682620
rect 154920 682380 155010 682620
rect 155250 682380 155340 682620
rect 155580 682380 155670 682620
rect 155910 682380 155930 682620
rect 144930 682290 155930 682380
rect 144930 682050 144950 682290
rect 145190 682050 145300 682290
rect 145540 682050 145630 682290
rect 145870 682050 145960 682290
rect 146200 682050 146290 682290
rect 146530 682050 146640 682290
rect 146880 682050 146970 682290
rect 147210 682050 147300 682290
rect 147540 682050 147630 682290
rect 147870 682050 147980 682290
rect 148220 682050 148310 682290
rect 148550 682050 148640 682290
rect 148880 682050 148970 682290
rect 149210 682050 149320 682290
rect 149560 682050 149650 682290
rect 149890 682050 149980 682290
rect 150220 682050 150310 682290
rect 150550 682050 150660 682290
rect 150900 682050 150990 682290
rect 151230 682050 151320 682290
rect 151560 682050 151650 682290
rect 151890 682050 152000 682290
rect 152240 682050 152330 682290
rect 152570 682050 152660 682290
rect 152900 682050 152990 682290
rect 153230 682050 153340 682290
rect 153580 682050 153670 682290
rect 153910 682050 154000 682290
rect 154240 682050 154330 682290
rect 154570 682050 154680 682290
rect 154920 682050 155010 682290
rect 155250 682050 155340 682290
rect 155580 682050 155670 682290
rect 155910 682050 155930 682290
rect 144930 681940 155930 682050
rect 144930 681700 144950 681940
rect 145190 681700 145300 681940
rect 145540 681700 145630 681940
rect 145870 681700 145960 681940
rect 146200 681700 146290 681940
rect 146530 681700 146640 681940
rect 146880 681700 146970 681940
rect 147210 681700 147300 681940
rect 147540 681700 147630 681940
rect 147870 681700 147980 681940
rect 148220 681700 148310 681940
rect 148550 681700 148640 681940
rect 148880 681700 148970 681940
rect 149210 681700 149320 681940
rect 149560 681700 149650 681940
rect 149890 681700 149980 681940
rect 150220 681700 150310 681940
rect 150550 681700 150660 681940
rect 150900 681700 150990 681940
rect 151230 681700 151320 681940
rect 151560 681700 151650 681940
rect 151890 681700 152000 681940
rect 152240 681700 152330 681940
rect 152570 681700 152660 681940
rect 152900 681700 152990 681940
rect 153230 681700 153340 681940
rect 153580 681700 153670 681940
rect 153910 681700 154000 681940
rect 154240 681700 154330 681940
rect 154570 681700 154680 681940
rect 154920 681700 155010 681940
rect 155250 681700 155340 681940
rect 155580 681700 155670 681940
rect 155910 681700 155930 681940
rect 144930 681610 155930 681700
rect 144930 681370 144950 681610
rect 145190 681370 145300 681610
rect 145540 681370 145630 681610
rect 145870 681370 145960 681610
rect 146200 681370 146290 681610
rect 146530 681370 146640 681610
rect 146880 681370 146970 681610
rect 147210 681370 147300 681610
rect 147540 681370 147630 681610
rect 147870 681370 147980 681610
rect 148220 681370 148310 681610
rect 148550 681370 148640 681610
rect 148880 681370 148970 681610
rect 149210 681370 149320 681610
rect 149560 681370 149650 681610
rect 149890 681370 149980 681610
rect 150220 681370 150310 681610
rect 150550 681370 150660 681610
rect 150900 681370 150990 681610
rect 151230 681370 151320 681610
rect 151560 681370 151650 681610
rect 151890 681370 152000 681610
rect 152240 681370 152330 681610
rect 152570 681370 152660 681610
rect 152900 681370 152990 681610
rect 153230 681370 153340 681610
rect 153580 681370 153670 681610
rect 153910 681370 154000 681610
rect 154240 681370 154330 681610
rect 154570 681370 154680 681610
rect 154920 681370 155010 681610
rect 155250 681370 155340 681610
rect 155580 681370 155670 681610
rect 155910 681370 155930 681610
rect 144930 681280 155930 681370
rect 144930 681040 144950 681280
rect 145190 681040 145300 681280
rect 145540 681040 145630 681280
rect 145870 681040 145960 681280
rect 146200 681040 146290 681280
rect 146530 681040 146640 681280
rect 146880 681040 146970 681280
rect 147210 681040 147300 681280
rect 147540 681040 147630 681280
rect 147870 681040 147980 681280
rect 148220 681040 148310 681280
rect 148550 681040 148640 681280
rect 148880 681040 148970 681280
rect 149210 681040 149320 681280
rect 149560 681040 149650 681280
rect 149890 681040 149980 681280
rect 150220 681040 150310 681280
rect 150550 681040 150660 681280
rect 150900 681040 150990 681280
rect 151230 681040 151320 681280
rect 151560 681040 151650 681280
rect 151890 681040 152000 681280
rect 152240 681040 152330 681280
rect 152570 681040 152660 681280
rect 152900 681040 152990 681280
rect 153230 681040 153340 681280
rect 153580 681040 153670 681280
rect 153910 681040 154000 681280
rect 154240 681040 154330 681280
rect 154570 681040 154680 681280
rect 154920 681040 155010 681280
rect 155250 681040 155340 681280
rect 155580 681040 155670 681280
rect 155910 681040 155930 681280
rect 144930 680950 155930 681040
rect 144930 680710 144950 680950
rect 145190 680710 145300 680950
rect 145540 680710 145630 680950
rect 145870 680710 145960 680950
rect 146200 680710 146290 680950
rect 146530 680710 146640 680950
rect 146880 680710 146970 680950
rect 147210 680710 147300 680950
rect 147540 680710 147630 680950
rect 147870 680710 147980 680950
rect 148220 680710 148310 680950
rect 148550 680710 148640 680950
rect 148880 680710 148970 680950
rect 149210 680710 149320 680950
rect 149560 680710 149650 680950
rect 149890 680710 149980 680950
rect 150220 680710 150310 680950
rect 150550 680710 150660 680950
rect 150900 680710 150990 680950
rect 151230 680710 151320 680950
rect 151560 680710 151650 680950
rect 151890 680710 152000 680950
rect 152240 680710 152330 680950
rect 152570 680710 152660 680950
rect 152900 680710 152990 680950
rect 153230 680710 153340 680950
rect 153580 680710 153670 680950
rect 153910 680710 154000 680950
rect 154240 680710 154330 680950
rect 154570 680710 154680 680950
rect 154920 680710 155010 680950
rect 155250 680710 155340 680950
rect 155580 680710 155670 680950
rect 155910 680710 155930 680950
rect 144930 680600 155930 680710
rect 144930 680360 144950 680600
rect 145190 680360 145300 680600
rect 145540 680360 145630 680600
rect 145870 680360 145960 680600
rect 146200 680360 146290 680600
rect 146530 680360 146640 680600
rect 146880 680360 146970 680600
rect 147210 680360 147300 680600
rect 147540 680360 147630 680600
rect 147870 680360 147980 680600
rect 148220 680360 148310 680600
rect 148550 680360 148640 680600
rect 148880 680360 148970 680600
rect 149210 680360 149320 680600
rect 149560 680360 149650 680600
rect 149890 680360 149980 680600
rect 150220 680360 150310 680600
rect 150550 680360 150660 680600
rect 150900 680360 150990 680600
rect 151230 680360 151320 680600
rect 151560 680360 151650 680600
rect 151890 680360 152000 680600
rect 152240 680360 152330 680600
rect 152570 680360 152660 680600
rect 152900 680360 152990 680600
rect 153230 680360 153340 680600
rect 153580 680360 153670 680600
rect 153910 680360 154000 680600
rect 154240 680360 154330 680600
rect 154570 680360 154680 680600
rect 154920 680360 155010 680600
rect 155250 680360 155340 680600
rect 155580 680360 155670 680600
rect 155910 680360 155930 680600
rect 144930 680270 155930 680360
rect 144930 680030 144950 680270
rect 145190 680030 145300 680270
rect 145540 680030 145630 680270
rect 145870 680030 145960 680270
rect 146200 680030 146290 680270
rect 146530 680030 146640 680270
rect 146880 680030 146970 680270
rect 147210 680030 147300 680270
rect 147540 680030 147630 680270
rect 147870 680030 147980 680270
rect 148220 680030 148310 680270
rect 148550 680030 148640 680270
rect 148880 680030 148970 680270
rect 149210 680030 149320 680270
rect 149560 680030 149650 680270
rect 149890 680030 149980 680270
rect 150220 680030 150310 680270
rect 150550 680030 150660 680270
rect 150900 680030 150990 680270
rect 151230 680030 151320 680270
rect 151560 680030 151650 680270
rect 151890 680030 152000 680270
rect 152240 680030 152330 680270
rect 152570 680030 152660 680270
rect 152900 680030 152990 680270
rect 153230 680030 153340 680270
rect 153580 680030 153670 680270
rect 153910 680030 154000 680270
rect 154240 680030 154330 680270
rect 154570 680030 154680 680270
rect 154920 680030 155010 680270
rect 155250 680030 155340 680270
rect 155580 680030 155670 680270
rect 155910 680030 155930 680270
rect 144930 679940 155930 680030
rect 144930 679700 144950 679940
rect 145190 679700 145300 679940
rect 145540 679700 145630 679940
rect 145870 679700 145960 679940
rect 146200 679700 146290 679940
rect 146530 679700 146640 679940
rect 146880 679700 146970 679940
rect 147210 679700 147300 679940
rect 147540 679700 147630 679940
rect 147870 679700 147980 679940
rect 148220 679700 148310 679940
rect 148550 679700 148640 679940
rect 148880 679700 148970 679940
rect 149210 679700 149320 679940
rect 149560 679700 149650 679940
rect 149890 679700 149980 679940
rect 150220 679700 150310 679940
rect 150550 679700 150660 679940
rect 150900 679700 150990 679940
rect 151230 679700 151320 679940
rect 151560 679700 151650 679940
rect 151890 679700 152000 679940
rect 152240 679700 152330 679940
rect 152570 679700 152660 679940
rect 152900 679700 152990 679940
rect 153230 679700 153340 679940
rect 153580 679700 153670 679940
rect 153910 679700 154000 679940
rect 154240 679700 154330 679940
rect 154570 679700 154680 679940
rect 154920 679700 155010 679940
rect 155250 679700 155340 679940
rect 155580 679700 155670 679940
rect 155910 679700 155930 679940
rect 144930 679610 155930 679700
rect 144930 679370 144950 679610
rect 145190 679370 145300 679610
rect 145540 679370 145630 679610
rect 145870 679370 145960 679610
rect 146200 679370 146290 679610
rect 146530 679370 146640 679610
rect 146880 679370 146970 679610
rect 147210 679370 147300 679610
rect 147540 679370 147630 679610
rect 147870 679370 147980 679610
rect 148220 679370 148310 679610
rect 148550 679370 148640 679610
rect 148880 679370 148970 679610
rect 149210 679370 149320 679610
rect 149560 679370 149650 679610
rect 149890 679370 149980 679610
rect 150220 679370 150310 679610
rect 150550 679370 150660 679610
rect 150900 679370 150990 679610
rect 151230 679370 151320 679610
rect 151560 679370 151650 679610
rect 151890 679370 152000 679610
rect 152240 679370 152330 679610
rect 152570 679370 152660 679610
rect 152900 679370 152990 679610
rect 153230 679370 153340 679610
rect 153580 679370 153670 679610
rect 153910 679370 154000 679610
rect 154240 679370 154330 679610
rect 154570 679370 154680 679610
rect 154920 679370 155010 679610
rect 155250 679370 155340 679610
rect 155580 679370 155670 679610
rect 155910 679370 155930 679610
rect 144930 679260 155930 679370
rect 144930 679020 144950 679260
rect 145190 679020 145300 679260
rect 145540 679020 145630 679260
rect 145870 679020 145960 679260
rect 146200 679020 146290 679260
rect 146530 679020 146640 679260
rect 146880 679020 146970 679260
rect 147210 679020 147300 679260
rect 147540 679020 147630 679260
rect 147870 679020 147980 679260
rect 148220 679020 148310 679260
rect 148550 679020 148640 679260
rect 148880 679020 148970 679260
rect 149210 679020 149320 679260
rect 149560 679020 149650 679260
rect 149890 679020 149980 679260
rect 150220 679020 150310 679260
rect 150550 679020 150660 679260
rect 150900 679020 150990 679260
rect 151230 679020 151320 679260
rect 151560 679020 151650 679260
rect 151890 679020 152000 679260
rect 152240 679020 152330 679260
rect 152570 679020 152660 679260
rect 152900 679020 152990 679260
rect 153230 679020 153340 679260
rect 153580 679020 153670 679260
rect 153910 679020 154000 679260
rect 154240 679020 154330 679260
rect 154570 679020 154680 679260
rect 154920 679020 155010 679260
rect 155250 679020 155340 679260
rect 155580 679020 155670 679260
rect 155910 679020 155930 679260
rect 144930 678930 155930 679020
rect 144930 678690 144950 678930
rect 145190 678690 145300 678930
rect 145540 678690 145630 678930
rect 145870 678690 145960 678930
rect 146200 678690 146290 678930
rect 146530 678690 146640 678930
rect 146880 678690 146970 678930
rect 147210 678690 147300 678930
rect 147540 678690 147630 678930
rect 147870 678690 147980 678930
rect 148220 678690 148310 678930
rect 148550 678690 148640 678930
rect 148880 678690 148970 678930
rect 149210 678690 149320 678930
rect 149560 678690 149650 678930
rect 149890 678690 149980 678930
rect 150220 678690 150310 678930
rect 150550 678690 150660 678930
rect 150900 678690 150990 678930
rect 151230 678690 151320 678930
rect 151560 678690 151650 678930
rect 151890 678690 152000 678930
rect 152240 678690 152330 678930
rect 152570 678690 152660 678930
rect 152900 678690 152990 678930
rect 153230 678690 153340 678930
rect 153580 678690 153670 678930
rect 153910 678690 154000 678930
rect 154240 678690 154330 678930
rect 154570 678690 154680 678930
rect 154920 678690 155010 678930
rect 155250 678690 155340 678930
rect 155580 678690 155670 678930
rect 155910 678690 155930 678930
rect 144930 678600 155930 678690
rect 144930 678360 144950 678600
rect 145190 678360 145300 678600
rect 145540 678360 145630 678600
rect 145870 678360 145960 678600
rect 146200 678360 146290 678600
rect 146530 678360 146640 678600
rect 146880 678360 146970 678600
rect 147210 678360 147300 678600
rect 147540 678360 147630 678600
rect 147870 678360 147980 678600
rect 148220 678360 148310 678600
rect 148550 678360 148640 678600
rect 148880 678360 148970 678600
rect 149210 678360 149320 678600
rect 149560 678360 149650 678600
rect 149890 678360 149980 678600
rect 150220 678360 150310 678600
rect 150550 678360 150660 678600
rect 150900 678360 150990 678600
rect 151230 678360 151320 678600
rect 151560 678360 151650 678600
rect 151890 678360 152000 678600
rect 152240 678360 152330 678600
rect 152570 678360 152660 678600
rect 152900 678360 152990 678600
rect 153230 678360 153340 678600
rect 153580 678360 153670 678600
rect 153910 678360 154000 678600
rect 154240 678360 154330 678600
rect 154570 678360 154680 678600
rect 154920 678360 155010 678600
rect 155250 678360 155340 678600
rect 155580 678360 155670 678600
rect 155910 678360 155930 678600
rect 144930 678270 155930 678360
rect 144930 678030 144950 678270
rect 145190 678030 145300 678270
rect 145540 678030 145630 678270
rect 145870 678030 145960 678270
rect 146200 678030 146290 678270
rect 146530 678030 146640 678270
rect 146880 678030 146970 678270
rect 147210 678030 147300 678270
rect 147540 678030 147630 678270
rect 147870 678030 147980 678270
rect 148220 678030 148310 678270
rect 148550 678030 148640 678270
rect 148880 678030 148970 678270
rect 149210 678030 149320 678270
rect 149560 678030 149650 678270
rect 149890 678030 149980 678270
rect 150220 678030 150310 678270
rect 150550 678030 150660 678270
rect 150900 678030 150990 678270
rect 151230 678030 151320 678270
rect 151560 678030 151650 678270
rect 151890 678030 152000 678270
rect 152240 678030 152330 678270
rect 152570 678030 152660 678270
rect 152900 678030 152990 678270
rect 153230 678030 153340 678270
rect 153580 678030 153670 678270
rect 153910 678030 154000 678270
rect 154240 678030 154330 678270
rect 154570 678030 154680 678270
rect 154920 678030 155010 678270
rect 155250 678030 155340 678270
rect 155580 678030 155670 678270
rect 155910 678030 155930 678270
rect 144930 677920 155930 678030
rect 144930 677680 144950 677920
rect 145190 677680 145300 677920
rect 145540 677680 145630 677920
rect 145870 677680 145960 677920
rect 146200 677680 146290 677920
rect 146530 677680 146640 677920
rect 146880 677680 146970 677920
rect 147210 677680 147300 677920
rect 147540 677680 147630 677920
rect 147870 677680 147980 677920
rect 148220 677680 148310 677920
rect 148550 677680 148640 677920
rect 148880 677680 148970 677920
rect 149210 677680 149320 677920
rect 149560 677680 149650 677920
rect 149890 677680 149980 677920
rect 150220 677680 150310 677920
rect 150550 677680 150660 677920
rect 150900 677680 150990 677920
rect 151230 677680 151320 677920
rect 151560 677680 151650 677920
rect 151890 677680 152000 677920
rect 152240 677680 152330 677920
rect 152570 677680 152660 677920
rect 152900 677680 152990 677920
rect 153230 677680 153340 677920
rect 153580 677680 153670 677920
rect 153910 677680 154000 677920
rect 154240 677680 154330 677920
rect 154570 677680 154680 677920
rect 154920 677680 155010 677920
rect 155250 677680 155340 677920
rect 155580 677680 155670 677920
rect 155910 677680 155930 677920
rect 144930 677590 155930 677680
rect 144930 677350 144950 677590
rect 145190 677350 145300 677590
rect 145540 677350 145630 677590
rect 145870 677350 145960 677590
rect 146200 677350 146290 677590
rect 146530 677350 146640 677590
rect 146880 677350 146970 677590
rect 147210 677350 147300 677590
rect 147540 677350 147630 677590
rect 147870 677350 147980 677590
rect 148220 677350 148310 677590
rect 148550 677350 148640 677590
rect 148880 677350 148970 677590
rect 149210 677350 149320 677590
rect 149560 677350 149650 677590
rect 149890 677350 149980 677590
rect 150220 677350 150310 677590
rect 150550 677350 150660 677590
rect 150900 677350 150990 677590
rect 151230 677350 151320 677590
rect 151560 677350 151650 677590
rect 151890 677350 152000 677590
rect 152240 677350 152330 677590
rect 152570 677350 152660 677590
rect 152900 677350 152990 677590
rect 153230 677350 153340 677590
rect 153580 677350 153670 677590
rect 153910 677350 154000 677590
rect 154240 677350 154330 677590
rect 154570 677350 154680 677590
rect 154920 677350 155010 677590
rect 155250 677350 155340 677590
rect 155580 677350 155670 677590
rect 155910 677350 155930 677590
rect 144930 677260 155930 677350
rect 144930 677020 144950 677260
rect 145190 677020 145300 677260
rect 145540 677020 145630 677260
rect 145870 677020 145960 677260
rect 146200 677020 146290 677260
rect 146530 677020 146640 677260
rect 146880 677020 146970 677260
rect 147210 677020 147300 677260
rect 147540 677020 147630 677260
rect 147870 677020 147980 677260
rect 148220 677020 148310 677260
rect 148550 677020 148640 677260
rect 148880 677020 148970 677260
rect 149210 677020 149320 677260
rect 149560 677020 149650 677260
rect 149890 677020 149980 677260
rect 150220 677020 150310 677260
rect 150550 677020 150660 677260
rect 150900 677020 150990 677260
rect 151230 677020 151320 677260
rect 151560 677020 151650 677260
rect 151890 677020 152000 677260
rect 152240 677020 152330 677260
rect 152570 677020 152660 677260
rect 152900 677020 152990 677260
rect 153230 677020 153340 677260
rect 153580 677020 153670 677260
rect 153910 677020 154000 677260
rect 154240 677020 154330 677260
rect 154570 677020 154680 677260
rect 154920 677020 155010 677260
rect 155250 677020 155340 677260
rect 155580 677020 155670 677260
rect 155910 677020 155930 677260
rect 144930 676930 155930 677020
rect 144930 676690 144950 676930
rect 145190 676690 145300 676930
rect 145540 676690 145630 676930
rect 145870 676690 145960 676930
rect 146200 676690 146290 676930
rect 146530 676690 146640 676930
rect 146880 676690 146970 676930
rect 147210 676690 147300 676930
rect 147540 676690 147630 676930
rect 147870 676690 147980 676930
rect 148220 676690 148310 676930
rect 148550 676690 148640 676930
rect 148880 676690 148970 676930
rect 149210 676690 149320 676930
rect 149560 676690 149650 676930
rect 149890 676690 149980 676930
rect 150220 676690 150310 676930
rect 150550 676690 150660 676930
rect 150900 676690 150990 676930
rect 151230 676690 151320 676930
rect 151560 676690 151650 676930
rect 151890 676690 152000 676930
rect 152240 676690 152330 676930
rect 152570 676690 152660 676930
rect 152900 676690 152990 676930
rect 153230 676690 153340 676930
rect 153580 676690 153670 676930
rect 153910 676690 154000 676930
rect 154240 676690 154330 676930
rect 154570 676690 154680 676930
rect 154920 676690 155010 676930
rect 155250 676690 155340 676930
rect 155580 676690 155670 676930
rect 155910 676690 155930 676930
rect 144930 676580 155930 676690
rect 144930 676340 144950 676580
rect 145190 676340 145300 676580
rect 145540 676340 145630 676580
rect 145870 676340 145960 676580
rect 146200 676340 146290 676580
rect 146530 676340 146640 676580
rect 146880 676340 146970 676580
rect 147210 676340 147300 676580
rect 147540 676340 147630 676580
rect 147870 676340 147980 676580
rect 148220 676340 148310 676580
rect 148550 676340 148640 676580
rect 148880 676340 148970 676580
rect 149210 676340 149320 676580
rect 149560 676340 149650 676580
rect 149890 676340 149980 676580
rect 150220 676340 150310 676580
rect 150550 676340 150660 676580
rect 150900 676340 150990 676580
rect 151230 676340 151320 676580
rect 151560 676340 151650 676580
rect 151890 676340 152000 676580
rect 152240 676340 152330 676580
rect 152570 676340 152660 676580
rect 152900 676340 152990 676580
rect 153230 676340 153340 676580
rect 153580 676340 153670 676580
rect 153910 676340 154000 676580
rect 154240 676340 154330 676580
rect 154570 676340 154680 676580
rect 154920 676340 155010 676580
rect 155250 676340 155340 676580
rect 155580 676340 155670 676580
rect 155910 676340 155930 676580
rect 144930 676250 155930 676340
rect 144930 676010 144950 676250
rect 145190 676010 145300 676250
rect 145540 676010 145630 676250
rect 145870 676010 145960 676250
rect 146200 676010 146290 676250
rect 146530 676010 146640 676250
rect 146880 676010 146970 676250
rect 147210 676010 147300 676250
rect 147540 676010 147630 676250
rect 147870 676010 147980 676250
rect 148220 676010 148310 676250
rect 148550 676010 148640 676250
rect 148880 676010 148970 676250
rect 149210 676010 149320 676250
rect 149560 676010 149650 676250
rect 149890 676010 149980 676250
rect 150220 676010 150310 676250
rect 150550 676010 150660 676250
rect 150900 676010 150990 676250
rect 151230 676010 151320 676250
rect 151560 676010 151650 676250
rect 151890 676010 152000 676250
rect 152240 676010 152330 676250
rect 152570 676010 152660 676250
rect 152900 676010 152990 676250
rect 153230 676010 153340 676250
rect 153580 676010 153670 676250
rect 153910 676010 154000 676250
rect 154240 676010 154330 676250
rect 154570 676010 154680 676250
rect 154920 676010 155010 676250
rect 155250 676010 155340 676250
rect 155580 676010 155670 676250
rect 155910 676010 155930 676250
rect 144930 675920 155930 676010
rect 144930 675680 144950 675920
rect 145190 675680 145300 675920
rect 145540 675680 145630 675920
rect 145870 675680 145960 675920
rect 146200 675680 146290 675920
rect 146530 675680 146640 675920
rect 146880 675680 146970 675920
rect 147210 675680 147300 675920
rect 147540 675680 147630 675920
rect 147870 675680 147980 675920
rect 148220 675680 148310 675920
rect 148550 675680 148640 675920
rect 148880 675680 148970 675920
rect 149210 675680 149320 675920
rect 149560 675680 149650 675920
rect 149890 675680 149980 675920
rect 150220 675680 150310 675920
rect 150550 675680 150660 675920
rect 150900 675680 150990 675920
rect 151230 675680 151320 675920
rect 151560 675680 151650 675920
rect 151890 675680 152000 675920
rect 152240 675680 152330 675920
rect 152570 675680 152660 675920
rect 152900 675680 152990 675920
rect 153230 675680 153340 675920
rect 153580 675680 153670 675920
rect 153910 675680 154000 675920
rect 154240 675680 154330 675920
rect 154570 675680 154680 675920
rect 154920 675680 155010 675920
rect 155250 675680 155340 675920
rect 155580 675680 155670 675920
rect 155910 675680 155930 675920
rect 144930 675590 155930 675680
rect 144930 675350 144950 675590
rect 145190 675350 145300 675590
rect 145540 675350 145630 675590
rect 145870 675350 145960 675590
rect 146200 675350 146290 675590
rect 146530 675350 146640 675590
rect 146880 675350 146970 675590
rect 147210 675350 147300 675590
rect 147540 675350 147630 675590
rect 147870 675350 147980 675590
rect 148220 675350 148310 675590
rect 148550 675350 148640 675590
rect 148880 675350 148970 675590
rect 149210 675350 149320 675590
rect 149560 675350 149650 675590
rect 149890 675350 149980 675590
rect 150220 675350 150310 675590
rect 150550 675350 150660 675590
rect 150900 675350 150990 675590
rect 151230 675350 151320 675590
rect 151560 675350 151650 675590
rect 151890 675350 152000 675590
rect 152240 675350 152330 675590
rect 152570 675350 152660 675590
rect 152900 675350 152990 675590
rect 153230 675350 153340 675590
rect 153580 675350 153670 675590
rect 153910 675350 154000 675590
rect 154240 675350 154330 675590
rect 154570 675350 154680 675590
rect 154920 675350 155010 675590
rect 155250 675350 155340 675590
rect 155580 675350 155670 675590
rect 155910 675350 155930 675590
rect 144930 675240 155930 675350
rect 144930 675000 144950 675240
rect 145190 675000 145300 675240
rect 145540 675000 145630 675240
rect 145870 675000 145960 675240
rect 146200 675000 146290 675240
rect 146530 675000 146640 675240
rect 146880 675000 146970 675240
rect 147210 675000 147300 675240
rect 147540 675000 147630 675240
rect 147870 675000 147980 675240
rect 148220 675000 148310 675240
rect 148550 675000 148640 675240
rect 148880 675000 148970 675240
rect 149210 675000 149320 675240
rect 149560 675000 149650 675240
rect 149890 675000 149980 675240
rect 150220 675000 150310 675240
rect 150550 675000 150660 675240
rect 150900 675000 150990 675240
rect 151230 675000 151320 675240
rect 151560 675000 151650 675240
rect 151890 675000 152000 675240
rect 152240 675000 152330 675240
rect 152570 675000 152660 675240
rect 152900 675000 152990 675240
rect 153230 675000 153340 675240
rect 153580 675000 153670 675240
rect 153910 675000 154000 675240
rect 154240 675000 154330 675240
rect 154570 675000 154680 675240
rect 154920 675000 155010 675240
rect 155250 675000 155340 675240
rect 155580 675000 155670 675240
rect 155910 675000 155930 675240
rect 144930 674910 155930 675000
rect 144930 674670 144950 674910
rect 145190 674670 145300 674910
rect 145540 674670 145630 674910
rect 145870 674670 145960 674910
rect 146200 674670 146290 674910
rect 146530 674670 146640 674910
rect 146880 674670 146970 674910
rect 147210 674670 147300 674910
rect 147540 674670 147630 674910
rect 147870 674670 147980 674910
rect 148220 674670 148310 674910
rect 148550 674670 148640 674910
rect 148880 674670 148970 674910
rect 149210 674670 149320 674910
rect 149560 674670 149650 674910
rect 149890 674670 149980 674910
rect 150220 674670 150310 674910
rect 150550 674670 150660 674910
rect 150900 674670 150990 674910
rect 151230 674670 151320 674910
rect 151560 674670 151650 674910
rect 151890 674670 152000 674910
rect 152240 674670 152330 674910
rect 152570 674670 152660 674910
rect 152900 674670 152990 674910
rect 153230 674670 153340 674910
rect 153580 674670 153670 674910
rect 153910 674670 154000 674910
rect 154240 674670 154330 674910
rect 154570 674670 154680 674910
rect 154920 674670 155010 674910
rect 155250 674670 155340 674910
rect 155580 674670 155670 674910
rect 155910 674670 155930 674910
rect 144930 674580 155930 674670
rect 144930 674340 144950 674580
rect 145190 674340 145300 674580
rect 145540 674340 145630 674580
rect 145870 674340 145960 674580
rect 146200 674340 146290 674580
rect 146530 674340 146640 674580
rect 146880 674340 146970 674580
rect 147210 674340 147300 674580
rect 147540 674340 147630 674580
rect 147870 674340 147980 674580
rect 148220 674340 148310 674580
rect 148550 674340 148640 674580
rect 148880 674340 148970 674580
rect 149210 674340 149320 674580
rect 149560 674340 149650 674580
rect 149890 674340 149980 674580
rect 150220 674340 150310 674580
rect 150550 674340 150660 674580
rect 150900 674340 150990 674580
rect 151230 674340 151320 674580
rect 151560 674340 151650 674580
rect 151890 674340 152000 674580
rect 152240 674340 152330 674580
rect 152570 674340 152660 674580
rect 152900 674340 152990 674580
rect 153230 674340 153340 674580
rect 153580 674340 153670 674580
rect 153910 674340 154000 674580
rect 154240 674340 154330 674580
rect 154570 674340 154680 674580
rect 154920 674340 155010 674580
rect 155250 674340 155340 674580
rect 155580 674340 155670 674580
rect 155910 674340 155930 674580
rect 144930 674250 155930 674340
rect 144930 674010 144950 674250
rect 145190 674010 145300 674250
rect 145540 674010 145630 674250
rect 145870 674010 145960 674250
rect 146200 674010 146290 674250
rect 146530 674010 146640 674250
rect 146880 674010 146970 674250
rect 147210 674010 147300 674250
rect 147540 674010 147630 674250
rect 147870 674010 147980 674250
rect 148220 674010 148310 674250
rect 148550 674010 148640 674250
rect 148880 674010 148970 674250
rect 149210 674010 149320 674250
rect 149560 674010 149650 674250
rect 149890 674010 149980 674250
rect 150220 674010 150310 674250
rect 150550 674010 150660 674250
rect 150900 674010 150990 674250
rect 151230 674010 151320 674250
rect 151560 674010 151650 674250
rect 151890 674010 152000 674250
rect 152240 674010 152330 674250
rect 152570 674010 152660 674250
rect 152900 674010 152990 674250
rect 153230 674010 153340 674250
rect 153580 674010 153670 674250
rect 153910 674010 154000 674250
rect 154240 674010 154330 674250
rect 154570 674010 154680 674250
rect 154920 674010 155010 674250
rect 155250 674010 155340 674250
rect 155580 674010 155670 674250
rect 155910 674010 155930 674250
rect 144930 673900 155930 674010
rect 144930 673660 144950 673900
rect 145190 673660 145300 673900
rect 145540 673660 145630 673900
rect 145870 673660 145960 673900
rect 146200 673660 146290 673900
rect 146530 673660 146640 673900
rect 146880 673660 146970 673900
rect 147210 673660 147300 673900
rect 147540 673660 147630 673900
rect 147870 673660 147980 673900
rect 148220 673660 148310 673900
rect 148550 673660 148640 673900
rect 148880 673660 148970 673900
rect 149210 673660 149320 673900
rect 149560 673660 149650 673900
rect 149890 673660 149980 673900
rect 150220 673660 150310 673900
rect 150550 673660 150660 673900
rect 150900 673660 150990 673900
rect 151230 673660 151320 673900
rect 151560 673660 151650 673900
rect 151890 673660 152000 673900
rect 152240 673660 152330 673900
rect 152570 673660 152660 673900
rect 152900 673660 152990 673900
rect 153230 673660 153340 673900
rect 153580 673660 153670 673900
rect 153910 673660 154000 673900
rect 154240 673660 154330 673900
rect 154570 673660 154680 673900
rect 154920 673660 155010 673900
rect 155250 673660 155340 673900
rect 155580 673660 155670 673900
rect 155910 673660 155930 673900
rect 144930 673570 155930 673660
rect 144930 673330 144950 673570
rect 145190 673330 145300 673570
rect 145540 673330 145630 673570
rect 145870 673330 145960 673570
rect 146200 673330 146290 673570
rect 146530 673330 146640 673570
rect 146880 673330 146970 673570
rect 147210 673330 147300 673570
rect 147540 673330 147630 673570
rect 147870 673330 147980 673570
rect 148220 673330 148310 673570
rect 148550 673330 148640 673570
rect 148880 673330 148970 673570
rect 149210 673330 149320 673570
rect 149560 673330 149650 673570
rect 149890 673330 149980 673570
rect 150220 673330 150310 673570
rect 150550 673330 150660 673570
rect 150900 673330 150990 673570
rect 151230 673330 151320 673570
rect 151560 673330 151650 673570
rect 151890 673330 152000 673570
rect 152240 673330 152330 673570
rect 152570 673330 152660 673570
rect 152900 673330 152990 673570
rect 153230 673330 153340 673570
rect 153580 673330 153670 673570
rect 153910 673330 154000 673570
rect 154240 673330 154330 673570
rect 154570 673330 154680 673570
rect 154920 673330 155010 673570
rect 155250 673330 155340 673570
rect 155580 673330 155670 673570
rect 155910 673330 155930 673570
rect 144930 673240 155930 673330
rect 144930 673000 144950 673240
rect 145190 673000 145300 673240
rect 145540 673000 145630 673240
rect 145870 673000 145960 673240
rect 146200 673000 146290 673240
rect 146530 673000 146640 673240
rect 146880 673000 146970 673240
rect 147210 673000 147300 673240
rect 147540 673000 147630 673240
rect 147870 673000 147980 673240
rect 148220 673000 148310 673240
rect 148550 673000 148640 673240
rect 148880 673000 148970 673240
rect 149210 673000 149320 673240
rect 149560 673000 149650 673240
rect 149890 673000 149980 673240
rect 150220 673000 150310 673240
rect 150550 673000 150660 673240
rect 150900 673000 150990 673240
rect 151230 673000 151320 673240
rect 151560 673000 151650 673240
rect 151890 673000 152000 673240
rect 152240 673000 152330 673240
rect 152570 673000 152660 673240
rect 152900 673000 152990 673240
rect 153230 673000 153340 673240
rect 153580 673000 153670 673240
rect 153910 673000 154000 673240
rect 154240 673000 154330 673240
rect 154570 673000 154680 673240
rect 154920 673000 155010 673240
rect 155250 673000 155340 673240
rect 155580 673000 155670 673240
rect 155910 673000 155930 673240
rect 144930 672910 155930 673000
rect 144930 672670 144950 672910
rect 145190 672670 145300 672910
rect 145540 672670 145630 672910
rect 145870 672670 145960 672910
rect 146200 672670 146290 672910
rect 146530 672670 146640 672910
rect 146880 672670 146970 672910
rect 147210 672670 147300 672910
rect 147540 672670 147630 672910
rect 147870 672670 147980 672910
rect 148220 672670 148310 672910
rect 148550 672670 148640 672910
rect 148880 672670 148970 672910
rect 149210 672670 149320 672910
rect 149560 672670 149650 672910
rect 149890 672670 149980 672910
rect 150220 672670 150310 672910
rect 150550 672670 150660 672910
rect 150900 672670 150990 672910
rect 151230 672670 151320 672910
rect 151560 672670 151650 672910
rect 151890 672670 152000 672910
rect 152240 672670 152330 672910
rect 152570 672670 152660 672910
rect 152900 672670 152990 672910
rect 153230 672670 153340 672910
rect 153580 672670 153670 672910
rect 153910 672670 154000 672910
rect 154240 672670 154330 672910
rect 154570 672670 154680 672910
rect 154920 672670 155010 672910
rect 155250 672670 155340 672910
rect 155580 672670 155670 672910
rect 155910 672670 155930 672910
rect 144930 672560 155930 672670
rect 144930 672320 144950 672560
rect 145190 672320 145300 672560
rect 145540 672320 145630 672560
rect 145870 672320 145960 672560
rect 146200 672320 146290 672560
rect 146530 672320 146640 672560
rect 146880 672320 146970 672560
rect 147210 672320 147300 672560
rect 147540 672320 147630 672560
rect 147870 672320 147980 672560
rect 148220 672320 148310 672560
rect 148550 672320 148640 672560
rect 148880 672320 148970 672560
rect 149210 672320 149320 672560
rect 149560 672320 149650 672560
rect 149890 672320 149980 672560
rect 150220 672320 150310 672560
rect 150550 672320 150660 672560
rect 150900 672320 150990 672560
rect 151230 672320 151320 672560
rect 151560 672320 151650 672560
rect 151890 672320 152000 672560
rect 152240 672320 152330 672560
rect 152570 672320 152660 672560
rect 152900 672320 152990 672560
rect 153230 672320 153340 672560
rect 153580 672320 153670 672560
rect 153910 672320 154000 672560
rect 154240 672320 154330 672560
rect 154570 672320 154680 672560
rect 154920 672320 155010 672560
rect 155250 672320 155340 672560
rect 155580 672320 155670 672560
rect 155910 672320 155930 672560
rect 144930 672300 155930 672320
rect 110790 671900 121790 671920
rect 110790 671660 110810 671900
rect 111050 671660 111140 671900
rect 111380 671660 111470 671900
rect 111710 671660 111800 671900
rect 112040 671660 112150 671900
rect 112390 671660 112480 671900
rect 112720 671660 112810 671900
rect 113050 671660 113140 671900
rect 113380 671660 113490 671900
rect 113730 671660 113820 671900
rect 114060 671660 114150 671900
rect 114390 671660 114480 671900
rect 114720 671660 114830 671900
rect 115070 671660 115160 671900
rect 115400 671660 115490 671900
rect 115730 671660 115820 671900
rect 116060 671660 116170 671900
rect 116410 671660 116500 671900
rect 116740 671660 116830 671900
rect 117070 671660 117160 671900
rect 117400 671660 117510 671900
rect 117750 671660 117840 671900
rect 118080 671660 118170 671900
rect 118410 671660 118500 671900
rect 118740 671660 118850 671900
rect 119090 671660 119180 671900
rect 119420 671660 119510 671900
rect 119750 671660 119840 671900
rect 120080 671660 120190 671900
rect 120430 671660 120520 671900
rect 120760 671660 120850 671900
rect 121090 671660 121180 671900
rect 121420 671660 121530 671900
rect 121770 671660 121790 671900
rect 110790 671550 121790 671660
rect 110790 671310 110810 671550
rect 111050 671310 111140 671550
rect 111380 671310 111470 671550
rect 111710 671310 111800 671550
rect 112040 671310 112150 671550
rect 112390 671310 112480 671550
rect 112720 671310 112810 671550
rect 113050 671310 113140 671550
rect 113380 671310 113490 671550
rect 113730 671310 113820 671550
rect 114060 671310 114150 671550
rect 114390 671310 114480 671550
rect 114720 671310 114830 671550
rect 115070 671310 115160 671550
rect 115400 671310 115490 671550
rect 115730 671310 115820 671550
rect 116060 671310 116170 671550
rect 116410 671310 116500 671550
rect 116740 671310 116830 671550
rect 117070 671310 117160 671550
rect 117400 671310 117510 671550
rect 117750 671310 117840 671550
rect 118080 671310 118170 671550
rect 118410 671310 118500 671550
rect 118740 671310 118850 671550
rect 119090 671310 119180 671550
rect 119420 671310 119510 671550
rect 119750 671310 119840 671550
rect 120080 671310 120190 671550
rect 120430 671310 120520 671550
rect 120760 671310 120850 671550
rect 121090 671310 121180 671550
rect 121420 671310 121530 671550
rect 121770 671310 121790 671550
rect 110790 671220 121790 671310
rect 110790 670980 110810 671220
rect 111050 670980 111140 671220
rect 111380 670980 111470 671220
rect 111710 670980 111800 671220
rect 112040 670980 112150 671220
rect 112390 670980 112480 671220
rect 112720 670980 112810 671220
rect 113050 670980 113140 671220
rect 113380 670980 113490 671220
rect 113730 670980 113820 671220
rect 114060 670980 114150 671220
rect 114390 670980 114480 671220
rect 114720 670980 114830 671220
rect 115070 670980 115160 671220
rect 115400 670980 115490 671220
rect 115730 670980 115820 671220
rect 116060 670980 116170 671220
rect 116410 670980 116500 671220
rect 116740 670980 116830 671220
rect 117070 670980 117160 671220
rect 117400 670980 117510 671220
rect 117750 670980 117840 671220
rect 118080 670980 118170 671220
rect 118410 670980 118500 671220
rect 118740 670980 118850 671220
rect 119090 670980 119180 671220
rect 119420 670980 119510 671220
rect 119750 670980 119840 671220
rect 120080 670980 120190 671220
rect 120430 670980 120520 671220
rect 120760 670980 120850 671220
rect 121090 670980 121180 671220
rect 121420 670980 121530 671220
rect 121770 670980 121790 671220
rect 110790 670890 121790 670980
rect 110790 670650 110810 670890
rect 111050 670650 111140 670890
rect 111380 670650 111470 670890
rect 111710 670650 111800 670890
rect 112040 670650 112150 670890
rect 112390 670650 112480 670890
rect 112720 670650 112810 670890
rect 113050 670650 113140 670890
rect 113380 670650 113490 670890
rect 113730 670650 113820 670890
rect 114060 670650 114150 670890
rect 114390 670650 114480 670890
rect 114720 670650 114830 670890
rect 115070 670650 115160 670890
rect 115400 670650 115490 670890
rect 115730 670650 115820 670890
rect 116060 670650 116170 670890
rect 116410 670650 116500 670890
rect 116740 670650 116830 670890
rect 117070 670650 117160 670890
rect 117400 670650 117510 670890
rect 117750 670650 117840 670890
rect 118080 670650 118170 670890
rect 118410 670650 118500 670890
rect 118740 670650 118850 670890
rect 119090 670650 119180 670890
rect 119420 670650 119510 670890
rect 119750 670650 119840 670890
rect 120080 670650 120190 670890
rect 120430 670650 120520 670890
rect 120760 670650 120850 670890
rect 121090 670650 121180 670890
rect 121420 670650 121530 670890
rect 121770 670650 121790 670890
rect 110790 670560 121790 670650
rect 110790 670320 110810 670560
rect 111050 670320 111140 670560
rect 111380 670320 111470 670560
rect 111710 670320 111800 670560
rect 112040 670320 112150 670560
rect 112390 670320 112480 670560
rect 112720 670320 112810 670560
rect 113050 670320 113140 670560
rect 113380 670320 113490 670560
rect 113730 670320 113820 670560
rect 114060 670320 114150 670560
rect 114390 670320 114480 670560
rect 114720 670320 114830 670560
rect 115070 670320 115160 670560
rect 115400 670320 115490 670560
rect 115730 670320 115820 670560
rect 116060 670320 116170 670560
rect 116410 670320 116500 670560
rect 116740 670320 116830 670560
rect 117070 670320 117160 670560
rect 117400 670320 117510 670560
rect 117750 670320 117840 670560
rect 118080 670320 118170 670560
rect 118410 670320 118500 670560
rect 118740 670320 118850 670560
rect 119090 670320 119180 670560
rect 119420 670320 119510 670560
rect 119750 670320 119840 670560
rect 120080 670320 120190 670560
rect 120430 670320 120520 670560
rect 120760 670320 120850 670560
rect 121090 670320 121180 670560
rect 121420 670320 121530 670560
rect 121770 670320 121790 670560
rect 110790 670210 121790 670320
rect 110790 669970 110810 670210
rect 111050 669970 111140 670210
rect 111380 669970 111470 670210
rect 111710 669970 111800 670210
rect 112040 669970 112150 670210
rect 112390 669970 112480 670210
rect 112720 669970 112810 670210
rect 113050 669970 113140 670210
rect 113380 669970 113490 670210
rect 113730 669970 113820 670210
rect 114060 669970 114150 670210
rect 114390 669970 114480 670210
rect 114720 669970 114830 670210
rect 115070 669970 115160 670210
rect 115400 669970 115490 670210
rect 115730 669970 115820 670210
rect 116060 669970 116170 670210
rect 116410 669970 116500 670210
rect 116740 669970 116830 670210
rect 117070 669970 117160 670210
rect 117400 669970 117510 670210
rect 117750 669970 117840 670210
rect 118080 669970 118170 670210
rect 118410 669970 118500 670210
rect 118740 669970 118850 670210
rect 119090 669970 119180 670210
rect 119420 669970 119510 670210
rect 119750 669970 119840 670210
rect 120080 669970 120190 670210
rect 120430 669970 120520 670210
rect 120760 669970 120850 670210
rect 121090 669970 121180 670210
rect 121420 669970 121530 670210
rect 121770 669970 121790 670210
rect 110790 669880 121790 669970
rect 110790 669640 110810 669880
rect 111050 669640 111140 669880
rect 111380 669640 111470 669880
rect 111710 669640 111800 669880
rect 112040 669640 112150 669880
rect 112390 669640 112480 669880
rect 112720 669640 112810 669880
rect 113050 669640 113140 669880
rect 113380 669640 113490 669880
rect 113730 669640 113820 669880
rect 114060 669640 114150 669880
rect 114390 669640 114480 669880
rect 114720 669640 114830 669880
rect 115070 669640 115160 669880
rect 115400 669640 115490 669880
rect 115730 669640 115820 669880
rect 116060 669640 116170 669880
rect 116410 669640 116500 669880
rect 116740 669640 116830 669880
rect 117070 669640 117160 669880
rect 117400 669640 117510 669880
rect 117750 669640 117840 669880
rect 118080 669640 118170 669880
rect 118410 669640 118500 669880
rect 118740 669640 118850 669880
rect 119090 669640 119180 669880
rect 119420 669640 119510 669880
rect 119750 669640 119840 669880
rect 120080 669640 120190 669880
rect 120430 669640 120520 669880
rect 120760 669640 120850 669880
rect 121090 669640 121180 669880
rect 121420 669640 121530 669880
rect 121770 669640 121790 669880
rect 110790 669550 121790 669640
rect 110790 669310 110810 669550
rect 111050 669310 111140 669550
rect 111380 669310 111470 669550
rect 111710 669310 111800 669550
rect 112040 669310 112150 669550
rect 112390 669310 112480 669550
rect 112720 669310 112810 669550
rect 113050 669310 113140 669550
rect 113380 669310 113490 669550
rect 113730 669310 113820 669550
rect 114060 669310 114150 669550
rect 114390 669310 114480 669550
rect 114720 669310 114830 669550
rect 115070 669310 115160 669550
rect 115400 669310 115490 669550
rect 115730 669310 115820 669550
rect 116060 669310 116170 669550
rect 116410 669310 116500 669550
rect 116740 669310 116830 669550
rect 117070 669310 117160 669550
rect 117400 669310 117510 669550
rect 117750 669310 117840 669550
rect 118080 669310 118170 669550
rect 118410 669310 118500 669550
rect 118740 669310 118850 669550
rect 119090 669310 119180 669550
rect 119420 669310 119510 669550
rect 119750 669310 119840 669550
rect 120080 669310 120190 669550
rect 120430 669310 120520 669550
rect 120760 669310 120850 669550
rect 121090 669310 121180 669550
rect 121420 669310 121530 669550
rect 121770 669310 121790 669550
rect 110790 669220 121790 669310
rect 110790 668980 110810 669220
rect 111050 668980 111140 669220
rect 111380 668980 111470 669220
rect 111710 668980 111800 669220
rect 112040 668980 112150 669220
rect 112390 668980 112480 669220
rect 112720 668980 112810 669220
rect 113050 668980 113140 669220
rect 113380 668980 113490 669220
rect 113730 668980 113820 669220
rect 114060 668980 114150 669220
rect 114390 668980 114480 669220
rect 114720 668980 114830 669220
rect 115070 668980 115160 669220
rect 115400 668980 115490 669220
rect 115730 668980 115820 669220
rect 116060 668980 116170 669220
rect 116410 668980 116500 669220
rect 116740 668980 116830 669220
rect 117070 668980 117160 669220
rect 117400 668980 117510 669220
rect 117750 668980 117840 669220
rect 118080 668980 118170 669220
rect 118410 668980 118500 669220
rect 118740 668980 118850 669220
rect 119090 668980 119180 669220
rect 119420 668980 119510 669220
rect 119750 668980 119840 669220
rect 120080 668980 120190 669220
rect 120430 668980 120520 669220
rect 120760 668980 120850 669220
rect 121090 668980 121180 669220
rect 121420 668980 121530 669220
rect 121770 668980 121790 669220
rect 110790 668870 121790 668980
rect 110790 668630 110810 668870
rect 111050 668630 111140 668870
rect 111380 668630 111470 668870
rect 111710 668630 111800 668870
rect 112040 668630 112150 668870
rect 112390 668630 112480 668870
rect 112720 668630 112810 668870
rect 113050 668630 113140 668870
rect 113380 668630 113490 668870
rect 113730 668630 113820 668870
rect 114060 668630 114150 668870
rect 114390 668630 114480 668870
rect 114720 668630 114830 668870
rect 115070 668630 115160 668870
rect 115400 668630 115490 668870
rect 115730 668630 115820 668870
rect 116060 668630 116170 668870
rect 116410 668630 116500 668870
rect 116740 668630 116830 668870
rect 117070 668630 117160 668870
rect 117400 668630 117510 668870
rect 117750 668630 117840 668870
rect 118080 668630 118170 668870
rect 118410 668630 118500 668870
rect 118740 668630 118850 668870
rect 119090 668630 119180 668870
rect 119420 668630 119510 668870
rect 119750 668630 119840 668870
rect 120080 668630 120190 668870
rect 120430 668630 120520 668870
rect 120760 668630 120850 668870
rect 121090 668630 121180 668870
rect 121420 668630 121530 668870
rect 121770 668630 121790 668870
rect 110790 668540 121790 668630
rect 110790 668300 110810 668540
rect 111050 668300 111140 668540
rect 111380 668300 111470 668540
rect 111710 668300 111800 668540
rect 112040 668300 112150 668540
rect 112390 668300 112480 668540
rect 112720 668300 112810 668540
rect 113050 668300 113140 668540
rect 113380 668300 113490 668540
rect 113730 668300 113820 668540
rect 114060 668300 114150 668540
rect 114390 668300 114480 668540
rect 114720 668300 114830 668540
rect 115070 668300 115160 668540
rect 115400 668300 115490 668540
rect 115730 668300 115820 668540
rect 116060 668300 116170 668540
rect 116410 668300 116500 668540
rect 116740 668300 116830 668540
rect 117070 668300 117160 668540
rect 117400 668300 117510 668540
rect 117750 668300 117840 668540
rect 118080 668300 118170 668540
rect 118410 668300 118500 668540
rect 118740 668300 118850 668540
rect 119090 668300 119180 668540
rect 119420 668300 119510 668540
rect 119750 668300 119840 668540
rect 120080 668300 120190 668540
rect 120430 668300 120520 668540
rect 120760 668300 120850 668540
rect 121090 668300 121180 668540
rect 121420 668300 121530 668540
rect 121770 668300 121790 668540
rect 110790 668210 121790 668300
rect 110790 667970 110810 668210
rect 111050 667970 111140 668210
rect 111380 667970 111470 668210
rect 111710 667970 111800 668210
rect 112040 667970 112150 668210
rect 112390 667970 112480 668210
rect 112720 667970 112810 668210
rect 113050 667970 113140 668210
rect 113380 667970 113490 668210
rect 113730 667970 113820 668210
rect 114060 667970 114150 668210
rect 114390 667970 114480 668210
rect 114720 667970 114830 668210
rect 115070 667970 115160 668210
rect 115400 667970 115490 668210
rect 115730 667970 115820 668210
rect 116060 667970 116170 668210
rect 116410 667970 116500 668210
rect 116740 667970 116830 668210
rect 117070 667970 117160 668210
rect 117400 667970 117510 668210
rect 117750 667970 117840 668210
rect 118080 667970 118170 668210
rect 118410 667970 118500 668210
rect 118740 667970 118850 668210
rect 119090 667970 119180 668210
rect 119420 667970 119510 668210
rect 119750 667970 119840 668210
rect 120080 667970 120190 668210
rect 120430 667970 120520 668210
rect 120760 667970 120850 668210
rect 121090 667970 121180 668210
rect 121420 667970 121530 668210
rect 121770 667970 121790 668210
rect 110790 667880 121790 667970
rect 110790 667640 110810 667880
rect 111050 667640 111140 667880
rect 111380 667640 111470 667880
rect 111710 667640 111800 667880
rect 112040 667640 112150 667880
rect 112390 667640 112480 667880
rect 112720 667640 112810 667880
rect 113050 667640 113140 667880
rect 113380 667640 113490 667880
rect 113730 667640 113820 667880
rect 114060 667640 114150 667880
rect 114390 667640 114480 667880
rect 114720 667640 114830 667880
rect 115070 667640 115160 667880
rect 115400 667640 115490 667880
rect 115730 667640 115820 667880
rect 116060 667640 116170 667880
rect 116410 667640 116500 667880
rect 116740 667640 116830 667880
rect 117070 667640 117160 667880
rect 117400 667640 117510 667880
rect 117750 667640 117840 667880
rect 118080 667640 118170 667880
rect 118410 667640 118500 667880
rect 118740 667640 118850 667880
rect 119090 667640 119180 667880
rect 119420 667640 119510 667880
rect 119750 667640 119840 667880
rect 120080 667640 120190 667880
rect 120430 667640 120520 667880
rect 120760 667640 120850 667880
rect 121090 667640 121180 667880
rect 121420 667640 121530 667880
rect 121770 667640 121790 667880
rect 110790 667530 121790 667640
rect 110790 667290 110810 667530
rect 111050 667290 111140 667530
rect 111380 667290 111470 667530
rect 111710 667290 111800 667530
rect 112040 667290 112150 667530
rect 112390 667290 112480 667530
rect 112720 667290 112810 667530
rect 113050 667290 113140 667530
rect 113380 667290 113490 667530
rect 113730 667290 113820 667530
rect 114060 667290 114150 667530
rect 114390 667290 114480 667530
rect 114720 667290 114830 667530
rect 115070 667290 115160 667530
rect 115400 667290 115490 667530
rect 115730 667290 115820 667530
rect 116060 667290 116170 667530
rect 116410 667290 116500 667530
rect 116740 667290 116830 667530
rect 117070 667290 117160 667530
rect 117400 667290 117510 667530
rect 117750 667290 117840 667530
rect 118080 667290 118170 667530
rect 118410 667290 118500 667530
rect 118740 667290 118850 667530
rect 119090 667290 119180 667530
rect 119420 667290 119510 667530
rect 119750 667290 119840 667530
rect 120080 667290 120190 667530
rect 120430 667290 120520 667530
rect 120760 667290 120850 667530
rect 121090 667290 121180 667530
rect 121420 667290 121530 667530
rect 121770 667290 121790 667530
rect 110790 667200 121790 667290
rect 110790 666960 110810 667200
rect 111050 666960 111140 667200
rect 111380 666960 111470 667200
rect 111710 666960 111800 667200
rect 112040 666960 112150 667200
rect 112390 666960 112480 667200
rect 112720 666960 112810 667200
rect 113050 666960 113140 667200
rect 113380 666960 113490 667200
rect 113730 666960 113820 667200
rect 114060 666960 114150 667200
rect 114390 666960 114480 667200
rect 114720 666960 114830 667200
rect 115070 666960 115160 667200
rect 115400 666960 115490 667200
rect 115730 666960 115820 667200
rect 116060 666960 116170 667200
rect 116410 666960 116500 667200
rect 116740 666960 116830 667200
rect 117070 666960 117160 667200
rect 117400 666960 117510 667200
rect 117750 666960 117840 667200
rect 118080 666960 118170 667200
rect 118410 666960 118500 667200
rect 118740 666960 118850 667200
rect 119090 666960 119180 667200
rect 119420 666960 119510 667200
rect 119750 666960 119840 667200
rect 120080 666960 120190 667200
rect 120430 666960 120520 667200
rect 120760 666960 120850 667200
rect 121090 666960 121180 667200
rect 121420 666960 121530 667200
rect 121770 666960 121790 667200
rect 110790 666870 121790 666960
rect 110790 666630 110810 666870
rect 111050 666630 111140 666870
rect 111380 666630 111470 666870
rect 111710 666630 111800 666870
rect 112040 666630 112150 666870
rect 112390 666630 112480 666870
rect 112720 666630 112810 666870
rect 113050 666630 113140 666870
rect 113380 666630 113490 666870
rect 113730 666630 113820 666870
rect 114060 666630 114150 666870
rect 114390 666630 114480 666870
rect 114720 666630 114830 666870
rect 115070 666630 115160 666870
rect 115400 666630 115490 666870
rect 115730 666630 115820 666870
rect 116060 666630 116170 666870
rect 116410 666630 116500 666870
rect 116740 666630 116830 666870
rect 117070 666630 117160 666870
rect 117400 666630 117510 666870
rect 117750 666630 117840 666870
rect 118080 666630 118170 666870
rect 118410 666630 118500 666870
rect 118740 666630 118850 666870
rect 119090 666630 119180 666870
rect 119420 666630 119510 666870
rect 119750 666630 119840 666870
rect 120080 666630 120190 666870
rect 120430 666630 120520 666870
rect 120760 666630 120850 666870
rect 121090 666630 121180 666870
rect 121420 666630 121530 666870
rect 121770 666630 121790 666870
rect 110790 666540 121790 666630
rect 110790 666300 110810 666540
rect 111050 666300 111140 666540
rect 111380 666300 111470 666540
rect 111710 666300 111800 666540
rect 112040 666300 112150 666540
rect 112390 666300 112480 666540
rect 112720 666300 112810 666540
rect 113050 666300 113140 666540
rect 113380 666300 113490 666540
rect 113730 666300 113820 666540
rect 114060 666300 114150 666540
rect 114390 666300 114480 666540
rect 114720 666300 114830 666540
rect 115070 666300 115160 666540
rect 115400 666300 115490 666540
rect 115730 666300 115820 666540
rect 116060 666300 116170 666540
rect 116410 666300 116500 666540
rect 116740 666300 116830 666540
rect 117070 666300 117160 666540
rect 117400 666300 117510 666540
rect 117750 666300 117840 666540
rect 118080 666300 118170 666540
rect 118410 666300 118500 666540
rect 118740 666300 118850 666540
rect 119090 666300 119180 666540
rect 119420 666300 119510 666540
rect 119750 666300 119840 666540
rect 120080 666300 120190 666540
rect 120430 666300 120520 666540
rect 120760 666300 120850 666540
rect 121090 666300 121180 666540
rect 121420 666300 121530 666540
rect 121770 666300 121790 666540
rect 110790 666190 121790 666300
rect 110790 665950 110810 666190
rect 111050 665950 111140 666190
rect 111380 665950 111470 666190
rect 111710 665950 111800 666190
rect 112040 665950 112150 666190
rect 112390 665950 112480 666190
rect 112720 665950 112810 666190
rect 113050 665950 113140 666190
rect 113380 665950 113490 666190
rect 113730 665950 113820 666190
rect 114060 665950 114150 666190
rect 114390 665950 114480 666190
rect 114720 665950 114830 666190
rect 115070 665950 115160 666190
rect 115400 665950 115490 666190
rect 115730 665950 115820 666190
rect 116060 665950 116170 666190
rect 116410 665950 116500 666190
rect 116740 665950 116830 666190
rect 117070 665950 117160 666190
rect 117400 665950 117510 666190
rect 117750 665950 117840 666190
rect 118080 665950 118170 666190
rect 118410 665950 118500 666190
rect 118740 665950 118850 666190
rect 119090 665950 119180 666190
rect 119420 665950 119510 666190
rect 119750 665950 119840 666190
rect 120080 665950 120190 666190
rect 120430 665950 120520 666190
rect 120760 665950 120850 666190
rect 121090 665950 121180 666190
rect 121420 665950 121530 666190
rect 121770 665950 121790 666190
rect 110790 665860 121790 665950
rect 110790 665620 110810 665860
rect 111050 665620 111140 665860
rect 111380 665620 111470 665860
rect 111710 665620 111800 665860
rect 112040 665620 112150 665860
rect 112390 665620 112480 665860
rect 112720 665620 112810 665860
rect 113050 665620 113140 665860
rect 113380 665620 113490 665860
rect 113730 665620 113820 665860
rect 114060 665620 114150 665860
rect 114390 665620 114480 665860
rect 114720 665620 114830 665860
rect 115070 665620 115160 665860
rect 115400 665620 115490 665860
rect 115730 665620 115820 665860
rect 116060 665620 116170 665860
rect 116410 665620 116500 665860
rect 116740 665620 116830 665860
rect 117070 665620 117160 665860
rect 117400 665620 117510 665860
rect 117750 665620 117840 665860
rect 118080 665620 118170 665860
rect 118410 665620 118500 665860
rect 118740 665620 118850 665860
rect 119090 665620 119180 665860
rect 119420 665620 119510 665860
rect 119750 665620 119840 665860
rect 120080 665620 120190 665860
rect 120430 665620 120520 665860
rect 120760 665620 120850 665860
rect 121090 665620 121180 665860
rect 121420 665620 121530 665860
rect 121770 665620 121790 665860
rect 110790 665530 121790 665620
rect 110790 665290 110810 665530
rect 111050 665290 111140 665530
rect 111380 665290 111470 665530
rect 111710 665290 111800 665530
rect 112040 665290 112150 665530
rect 112390 665290 112480 665530
rect 112720 665290 112810 665530
rect 113050 665290 113140 665530
rect 113380 665290 113490 665530
rect 113730 665290 113820 665530
rect 114060 665290 114150 665530
rect 114390 665290 114480 665530
rect 114720 665290 114830 665530
rect 115070 665290 115160 665530
rect 115400 665290 115490 665530
rect 115730 665290 115820 665530
rect 116060 665290 116170 665530
rect 116410 665290 116500 665530
rect 116740 665290 116830 665530
rect 117070 665290 117160 665530
rect 117400 665290 117510 665530
rect 117750 665290 117840 665530
rect 118080 665290 118170 665530
rect 118410 665290 118500 665530
rect 118740 665290 118850 665530
rect 119090 665290 119180 665530
rect 119420 665290 119510 665530
rect 119750 665290 119840 665530
rect 120080 665290 120190 665530
rect 120430 665290 120520 665530
rect 120760 665290 120850 665530
rect 121090 665290 121180 665530
rect 121420 665290 121530 665530
rect 121770 665290 121790 665530
rect 110790 665200 121790 665290
rect 110790 664960 110810 665200
rect 111050 664960 111140 665200
rect 111380 664960 111470 665200
rect 111710 664960 111800 665200
rect 112040 664960 112150 665200
rect 112390 664960 112480 665200
rect 112720 664960 112810 665200
rect 113050 664960 113140 665200
rect 113380 664960 113490 665200
rect 113730 664960 113820 665200
rect 114060 664960 114150 665200
rect 114390 664960 114480 665200
rect 114720 664960 114830 665200
rect 115070 664960 115160 665200
rect 115400 664960 115490 665200
rect 115730 664960 115820 665200
rect 116060 664960 116170 665200
rect 116410 664960 116500 665200
rect 116740 664960 116830 665200
rect 117070 664960 117160 665200
rect 117400 664960 117510 665200
rect 117750 664960 117840 665200
rect 118080 664960 118170 665200
rect 118410 664960 118500 665200
rect 118740 664960 118850 665200
rect 119090 664960 119180 665200
rect 119420 664960 119510 665200
rect 119750 664960 119840 665200
rect 120080 664960 120190 665200
rect 120430 664960 120520 665200
rect 120760 664960 120850 665200
rect 121090 664960 121180 665200
rect 121420 664960 121530 665200
rect 121770 664960 121790 665200
rect 110790 664850 121790 664960
rect 110790 664610 110810 664850
rect 111050 664610 111140 664850
rect 111380 664610 111470 664850
rect 111710 664610 111800 664850
rect 112040 664610 112150 664850
rect 112390 664610 112480 664850
rect 112720 664610 112810 664850
rect 113050 664610 113140 664850
rect 113380 664610 113490 664850
rect 113730 664610 113820 664850
rect 114060 664610 114150 664850
rect 114390 664610 114480 664850
rect 114720 664610 114830 664850
rect 115070 664610 115160 664850
rect 115400 664610 115490 664850
rect 115730 664610 115820 664850
rect 116060 664610 116170 664850
rect 116410 664610 116500 664850
rect 116740 664610 116830 664850
rect 117070 664610 117160 664850
rect 117400 664610 117510 664850
rect 117750 664610 117840 664850
rect 118080 664610 118170 664850
rect 118410 664610 118500 664850
rect 118740 664610 118850 664850
rect 119090 664610 119180 664850
rect 119420 664610 119510 664850
rect 119750 664610 119840 664850
rect 120080 664610 120190 664850
rect 120430 664610 120520 664850
rect 120760 664610 120850 664850
rect 121090 664610 121180 664850
rect 121420 664610 121530 664850
rect 121770 664610 121790 664850
rect 110790 664520 121790 664610
rect 110790 664280 110810 664520
rect 111050 664280 111140 664520
rect 111380 664280 111470 664520
rect 111710 664280 111800 664520
rect 112040 664280 112150 664520
rect 112390 664280 112480 664520
rect 112720 664280 112810 664520
rect 113050 664280 113140 664520
rect 113380 664280 113490 664520
rect 113730 664280 113820 664520
rect 114060 664280 114150 664520
rect 114390 664280 114480 664520
rect 114720 664280 114830 664520
rect 115070 664280 115160 664520
rect 115400 664280 115490 664520
rect 115730 664280 115820 664520
rect 116060 664280 116170 664520
rect 116410 664280 116500 664520
rect 116740 664280 116830 664520
rect 117070 664280 117160 664520
rect 117400 664280 117510 664520
rect 117750 664280 117840 664520
rect 118080 664280 118170 664520
rect 118410 664280 118500 664520
rect 118740 664280 118850 664520
rect 119090 664280 119180 664520
rect 119420 664280 119510 664520
rect 119750 664280 119840 664520
rect 120080 664280 120190 664520
rect 120430 664280 120520 664520
rect 120760 664280 120850 664520
rect 121090 664280 121180 664520
rect 121420 664280 121530 664520
rect 121770 664280 121790 664520
rect 110790 664190 121790 664280
rect 110790 663950 110810 664190
rect 111050 663950 111140 664190
rect 111380 663950 111470 664190
rect 111710 663950 111800 664190
rect 112040 663950 112150 664190
rect 112390 663950 112480 664190
rect 112720 663950 112810 664190
rect 113050 663950 113140 664190
rect 113380 663950 113490 664190
rect 113730 663950 113820 664190
rect 114060 663950 114150 664190
rect 114390 663950 114480 664190
rect 114720 663950 114830 664190
rect 115070 663950 115160 664190
rect 115400 663950 115490 664190
rect 115730 663950 115820 664190
rect 116060 663950 116170 664190
rect 116410 663950 116500 664190
rect 116740 663950 116830 664190
rect 117070 663950 117160 664190
rect 117400 663950 117510 664190
rect 117750 663950 117840 664190
rect 118080 663950 118170 664190
rect 118410 663950 118500 664190
rect 118740 663950 118850 664190
rect 119090 663950 119180 664190
rect 119420 663950 119510 664190
rect 119750 663950 119840 664190
rect 120080 663950 120190 664190
rect 120430 663950 120520 664190
rect 120760 663950 120850 664190
rect 121090 663950 121180 664190
rect 121420 663950 121530 664190
rect 121770 663950 121790 664190
rect 110790 663860 121790 663950
rect 110790 663620 110810 663860
rect 111050 663620 111140 663860
rect 111380 663620 111470 663860
rect 111710 663620 111800 663860
rect 112040 663620 112150 663860
rect 112390 663620 112480 663860
rect 112720 663620 112810 663860
rect 113050 663620 113140 663860
rect 113380 663620 113490 663860
rect 113730 663620 113820 663860
rect 114060 663620 114150 663860
rect 114390 663620 114480 663860
rect 114720 663620 114830 663860
rect 115070 663620 115160 663860
rect 115400 663620 115490 663860
rect 115730 663620 115820 663860
rect 116060 663620 116170 663860
rect 116410 663620 116500 663860
rect 116740 663620 116830 663860
rect 117070 663620 117160 663860
rect 117400 663620 117510 663860
rect 117750 663620 117840 663860
rect 118080 663620 118170 663860
rect 118410 663620 118500 663860
rect 118740 663620 118850 663860
rect 119090 663620 119180 663860
rect 119420 663620 119510 663860
rect 119750 663620 119840 663860
rect 120080 663620 120190 663860
rect 120430 663620 120520 663860
rect 120760 663620 120850 663860
rect 121090 663620 121180 663860
rect 121420 663620 121530 663860
rect 121770 663620 121790 663860
rect 110790 663510 121790 663620
rect 110790 663270 110810 663510
rect 111050 663270 111140 663510
rect 111380 663270 111470 663510
rect 111710 663270 111800 663510
rect 112040 663270 112150 663510
rect 112390 663270 112480 663510
rect 112720 663270 112810 663510
rect 113050 663270 113140 663510
rect 113380 663270 113490 663510
rect 113730 663270 113820 663510
rect 114060 663270 114150 663510
rect 114390 663270 114480 663510
rect 114720 663270 114830 663510
rect 115070 663270 115160 663510
rect 115400 663270 115490 663510
rect 115730 663270 115820 663510
rect 116060 663270 116170 663510
rect 116410 663270 116500 663510
rect 116740 663270 116830 663510
rect 117070 663270 117160 663510
rect 117400 663270 117510 663510
rect 117750 663270 117840 663510
rect 118080 663270 118170 663510
rect 118410 663270 118500 663510
rect 118740 663270 118850 663510
rect 119090 663270 119180 663510
rect 119420 663270 119510 663510
rect 119750 663270 119840 663510
rect 120080 663270 120190 663510
rect 120430 663270 120520 663510
rect 120760 663270 120850 663510
rect 121090 663270 121180 663510
rect 121420 663270 121530 663510
rect 121770 663270 121790 663510
rect 110790 663180 121790 663270
rect 110790 662940 110810 663180
rect 111050 662940 111140 663180
rect 111380 662940 111470 663180
rect 111710 662940 111800 663180
rect 112040 662940 112150 663180
rect 112390 662940 112480 663180
rect 112720 662940 112810 663180
rect 113050 662940 113140 663180
rect 113380 662940 113490 663180
rect 113730 662940 113820 663180
rect 114060 662940 114150 663180
rect 114390 662940 114480 663180
rect 114720 662940 114830 663180
rect 115070 662940 115160 663180
rect 115400 662940 115490 663180
rect 115730 662940 115820 663180
rect 116060 662940 116170 663180
rect 116410 662940 116500 663180
rect 116740 662940 116830 663180
rect 117070 662940 117160 663180
rect 117400 662940 117510 663180
rect 117750 662940 117840 663180
rect 118080 662940 118170 663180
rect 118410 662940 118500 663180
rect 118740 662940 118850 663180
rect 119090 662940 119180 663180
rect 119420 662940 119510 663180
rect 119750 662940 119840 663180
rect 120080 662940 120190 663180
rect 120430 662940 120520 663180
rect 120760 662940 120850 663180
rect 121090 662940 121180 663180
rect 121420 662940 121530 663180
rect 121770 662940 121790 663180
rect 110790 662850 121790 662940
rect 110790 662610 110810 662850
rect 111050 662610 111140 662850
rect 111380 662610 111470 662850
rect 111710 662610 111800 662850
rect 112040 662610 112150 662850
rect 112390 662610 112480 662850
rect 112720 662610 112810 662850
rect 113050 662610 113140 662850
rect 113380 662610 113490 662850
rect 113730 662610 113820 662850
rect 114060 662610 114150 662850
rect 114390 662610 114480 662850
rect 114720 662610 114830 662850
rect 115070 662610 115160 662850
rect 115400 662610 115490 662850
rect 115730 662610 115820 662850
rect 116060 662610 116170 662850
rect 116410 662610 116500 662850
rect 116740 662610 116830 662850
rect 117070 662610 117160 662850
rect 117400 662610 117510 662850
rect 117750 662610 117840 662850
rect 118080 662610 118170 662850
rect 118410 662610 118500 662850
rect 118740 662610 118850 662850
rect 119090 662610 119180 662850
rect 119420 662610 119510 662850
rect 119750 662610 119840 662850
rect 120080 662610 120190 662850
rect 120430 662610 120520 662850
rect 120760 662610 120850 662850
rect 121090 662610 121180 662850
rect 121420 662610 121530 662850
rect 121770 662610 121790 662850
rect 110790 662520 121790 662610
rect 110790 662280 110810 662520
rect 111050 662280 111140 662520
rect 111380 662280 111470 662520
rect 111710 662280 111800 662520
rect 112040 662280 112150 662520
rect 112390 662280 112480 662520
rect 112720 662280 112810 662520
rect 113050 662280 113140 662520
rect 113380 662280 113490 662520
rect 113730 662280 113820 662520
rect 114060 662280 114150 662520
rect 114390 662280 114480 662520
rect 114720 662280 114830 662520
rect 115070 662280 115160 662520
rect 115400 662280 115490 662520
rect 115730 662280 115820 662520
rect 116060 662280 116170 662520
rect 116410 662280 116500 662520
rect 116740 662280 116830 662520
rect 117070 662280 117160 662520
rect 117400 662280 117510 662520
rect 117750 662280 117840 662520
rect 118080 662280 118170 662520
rect 118410 662280 118500 662520
rect 118740 662280 118850 662520
rect 119090 662280 119180 662520
rect 119420 662280 119510 662520
rect 119750 662280 119840 662520
rect 120080 662280 120190 662520
rect 120430 662280 120520 662520
rect 120760 662280 120850 662520
rect 121090 662280 121180 662520
rect 121420 662280 121530 662520
rect 121770 662280 121790 662520
rect 110790 662170 121790 662280
rect 110790 661930 110810 662170
rect 111050 661930 111140 662170
rect 111380 661930 111470 662170
rect 111710 661930 111800 662170
rect 112040 661930 112150 662170
rect 112390 661930 112480 662170
rect 112720 661930 112810 662170
rect 113050 661930 113140 662170
rect 113380 661930 113490 662170
rect 113730 661930 113820 662170
rect 114060 661930 114150 662170
rect 114390 661930 114480 662170
rect 114720 661930 114830 662170
rect 115070 661930 115160 662170
rect 115400 661930 115490 662170
rect 115730 661930 115820 662170
rect 116060 661930 116170 662170
rect 116410 661930 116500 662170
rect 116740 661930 116830 662170
rect 117070 661930 117160 662170
rect 117400 661930 117510 662170
rect 117750 661930 117840 662170
rect 118080 661930 118170 662170
rect 118410 661930 118500 662170
rect 118740 661930 118850 662170
rect 119090 661930 119180 662170
rect 119420 661930 119510 662170
rect 119750 661930 119840 662170
rect 120080 661930 120190 662170
rect 120430 661930 120520 662170
rect 120760 661930 120850 662170
rect 121090 661930 121180 662170
rect 121420 661930 121530 662170
rect 121770 661930 121790 662170
rect 110790 661840 121790 661930
rect 110790 661600 110810 661840
rect 111050 661600 111140 661840
rect 111380 661600 111470 661840
rect 111710 661600 111800 661840
rect 112040 661600 112150 661840
rect 112390 661600 112480 661840
rect 112720 661600 112810 661840
rect 113050 661600 113140 661840
rect 113380 661600 113490 661840
rect 113730 661600 113820 661840
rect 114060 661600 114150 661840
rect 114390 661600 114480 661840
rect 114720 661600 114830 661840
rect 115070 661600 115160 661840
rect 115400 661600 115490 661840
rect 115730 661600 115820 661840
rect 116060 661600 116170 661840
rect 116410 661600 116500 661840
rect 116740 661600 116830 661840
rect 117070 661600 117160 661840
rect 117400 661600 117510 661840
rect 117750 661600 117840 661840
rect 118080 661600 118170 661840
rect 118410 661600 118500 661840
rect 118740 661600 118850 661840
rect 119090 661600 119180 661840
rect 119420 661600 119510 661840
rect 119750 661600 119840 661840
rect 120080 661600 120190 661840
rect 120430 661600 120520 661840
rect 120760 661600 120850 661840
rect 121090 661600 121180 661840
rect 121420 661600 121530 661840
rect 121770 661600 121790 661840
rect 110790 661510 121790 661600
rect 110790 661270 110810 661510
rect 111050 661270 111140 661510
rect 111380 661270 111470 661510
rect 111710 661270 111800 661510
rect 112040 661270 112150 661510
rect 112390 661270 112480 661510
rect 112720 661270 112810 661510
rect 113050 661270 113140 661510
rect 113380 661270 113490 661510
rect 113730 661270 113820 661510
rect 114060 661270 114150 661510
rect 114390 661270 114480 661510
rect 114720 661270 114830 661510
rect 115070 661270 115160 661510
rect 115400 661270 115490 661510
rect 115730 661270 115820 661510
rect 116060 661270 116170 661510
rect 116410 661270 116500 661510
rect 116740 661270 116830 661510
rect 117070 661270 117160 661510
rect 117400 661270 117510 661510
rect 117750 661270 117840 661510
rect 118080 661270 118170 661510
rect 118410 661270 118500 661510
rect 118740 661270 118850 661510
rect 119090 661270 119180 661510
rect 119420 661270 119510 661510
rect 119750 661270 119840 661510
rect 120080 661270 120190 661510
rect 120430 661270 120520 661510
rect 120760 661270 120850 661510
rect 121090 661270 121180 661510
rect 121420 661270 121530 661510
rect 121770 661270 121790 661510
rect 110790 661180 121790 661270
rect 110790 660940 110810 661180
rect 111050 660940 111140 661180
rect 111380 660940 111470 661180
rect 111710 660940 111800 661180
rect 112040 660940 112150 661180
rect 112390 660940 112480 661180
rect 112720 660940 112810 661180
rect 113050 660940 113140 661180
rect 113380 660940 113490 661180
rect 113730 660940 113820 661180
rect 114060 660940 114150 661180
rect 114390 660940 114480 661180
rect 114720 660940 114830 661180
rect 115070 660940 115160 661180
rect 115400 660940 115490 661180
rect 115730 660940 115820 661180
rect 116060 660940 116170 661180
rect 116410 660940 116500 661180
rect 116740 660940 116830 661180
rect 117070 660940 117160 661180
rect 117400 660940 117510 661180
rect 117750 660940 117840 661180
rect 118080 660940 118170 661180
rect 118410 660940 118500 661180
rect 118740 660940 118850 661180
rect 119090 660940 119180 661180
rect 119420 660940 119510 661180
rect 119750 660940 119840 661180
rect 120080 660940 120190 661180
rect 120430 660940 120520 661180
rect 120760 660940 120850 661180
rect 121090 660940 121180 661180
rect 121420 660940 121530 661180
rect 121770 660940 121790 661180
rect 110790 660920 121790 660940
rect 122170 671900 133170 671920
rect 122170 671660 122190 671900
rect 122430 671660 122520 671900
rect 122760 671660 122850 671900
rect 123090 671660 123180 671900
rect 123420 671660 123530 671900
rect 123770 671660 123860 671900
rect 124100 671660 124190 671900
rect 124430 671660 124520 671900
rect 124760 671660 124870 671900
rect 125110 671660 125200 671900
rect 125440 671660 125530 671900
rect 125770 671660 125860 671900
rect 126100 671660 126210 671900
rect 126450 671660 126540 671900
rect 126780 671660 126870 671900
rect 127110 671660 127200 671900
rect 127440 671660 127550 671900
rect 127790 671660 127880 671900
rect 128120 671660 128210 671900
rect 128450 671660 128540 671900
rect 128780 671660 128890 671900
rect 129130 671660 129220 671900
rect 129460 671660 129550 671900
rect 129790 671660 129880 671900
rect 130120 671660 130230 671900
rect 130470 671660 130560 671900
rect 130800 671660 130890 671900
rect 131130 671660 131220 671900
rect 131460 671660 131570 671900
rect 131810 671660 131900 671900
rect 132140 671660 132230 671900
rect 132470 671660 132560 671900
rect 132800 671660 132910 671900
rect 133150 671660 133170 671900
rect 122170 671550 133170 671660
rect 122170 671310 122190 671550
rect 122430 671310 122520 671550
rect 122760 671310 122850 671550
rect 123090 671310 123180 671550
rect 123420 671310 123530 671550
rect 123770 671310 123860 671550
rect 124100 671310 124190 671550
rect 124430 671310 124520 671550
rect 124760 671310 124870 671550
rect 125110 671310 125200 671550
rect 125440 671310 125530 671550
rect 125770 671310 125860 671550
rect 126100 671310 126210 671550
rect 126450 671310 126540 671550
rect 126780 671310 126870 671550
rect 127110 671310 127200 671550
rect 127440 671310 127550 671550
rect 127790 671310 127880 671550
rect 128120 671310 128210 671550
rect 128450 671310 128540 671550
rect 128780 671310 128890 671550
rect 129130 671310 129220 671550
rect 129460 671310 129550 671550
rect 129790 671310 129880 671550
rect 130120 671310 130230 671550
rect 130470 671310 130560 671550
rect 130800 671310 130890 671550
rect 131130 671310 131220 671550
rect 131460 671310 131570 671550
rect 131810 671310 131900 671550
rect 132140 671310 132230 671550
rect 132470 671310 132560 671550
rect 132800 671310 132910 671550
rect 133150 671310 133170 671550
rect 122170 671220 133170 671310
rect 122170 670980 122190 671220
rect 122430 670980 122520 671220
rect 122760 670980 122850 671220
rect 123090 670980 123180 671220
rect 123420 670980 123530 671220
rect 123770 670980 123860 671220
rect 124100 670980 124190 671220
rect 124430 670980 124520 671220
rect 124760 670980 124870 671220
rect 125110 670980 125200 671220
rect 125440 670980 125530 671220
rect 125770 670980 125860 671220
rect 126100 670980 126210 671220
rect 126450 670980 126540 671220
rect 126780 670980 126870 671220
rect 127110 670980 127200 671220
rect 127440 670980 127550 671220
rect 127790 670980 127880 671220
rect 128120 670980 128210 671220
rect 128450 670980 128540 671220
rect 128780 670980 128890 671220
rect 129130 670980 129220 671220
rect 129460 670980 129550 671220
rect 129790 670980 129880 671220
rect 130120 670980 130230 671220
rect 130470 670980 130560 671220
rect 130800 670980 130890 671220
rect 131130 670980 131220 671220
rect 131460 670980 131570 671220
rect 131810 670980 131900 671220
rect 132140 670980 132230 671220
rect 132470 670980 132560 671220
rect 132800 670980 132910 671220
rect 133150 670980 133170 671220
rect 122170 670890 133170 670980
rect 122170 670650 122190 670890
rect 122430 670650 122520 670890
rect 122760 670650 122850 670890
rect 123090 670650 123180 670890
rect 123420 670650 123530 670890
rect 123770 670650 123860 670890
rect 124100 670650 124190 670890
rect 124430 670650 124520 670890
rect 124760 670650 124870 670890
rect 125110 670650 125200 670890
rect 125440 670650 125530 670890
rect 125770 670650 125860 670890
rect 126100 670650 126210 670890
rect 126450 670650 126540 670890
rect 126780 670650 126870 670890
rect 127110 670650 127200 670890
rect 127440 670650 127550 670890
rect 127790 670650 127880 670890
rect 128120 670650 128210 670890
rect 128450 670650 128540 670890
rect 128780 670650 128890 670890
rect 129130 670650 129220 670890
rect 129460 670650 129550 670890
rect 129790 670650 129880 670890
rect 130120 670650 130230 670890
rect 130470 670650 130560 670890
rect 130800 670650 130890 670890
rect 131130 670650 131220 670890
rect 131460 670650 131570 670890
rect 131810 670650 131900 670890
rect 132140 670650 132230 670890
rect 132470 670650 132560 670890
rect 132800 670650 132910 670890
rect 133150 670650 133170 670890
rect 122170 670560 133170 670650
rect 122170 670320 122190 670560
rect 122430 670320 122520 670560
rect 122760 670320 122850 670560
rect 123090 670320 123180 670560
rect 123420 670320 123530 670560
rect 123770 670320 123860 670560
rect 124100 670320 124190 670560
rect 124430 670320 124520 670560
rect 124760 670320 124870 670560
rect 125110 670320 125200 670560
rect 125440 670320 125530 670560
rect 125770 670320 125860 670560
rect 126100 670320 126210 670560
rect 126450 670320 126540 670560
rect 126780 670320 126870 670560
rect 127110 670320 127200 670560
rect 127440 670320 127550 670560
rect 127790 670320 127880 670560
rect 128120 670320 128210 670560
rect 128450 670320 128540 670560
rect 128780 670320 128890 670560
rect 129130 670320 129220 670560
rect 129460 670320 129550 670560
rect 129790 670320 129880 670560
rect 130120 670320 130230 670560
rect 130470 670320 130560 670560
rect 130800 670320 130890 670560
rect 131130 670320 131220 670560
rect 131460 670320 131570 670560
rect 131810 670320 131900 670560
rect 132140 670320 132230 670560
rect 132470 670320 132560 670560
rect 132800 670320 132910 670560
rect 133150 670320 133170 670560
rect 122170 670210 133170 670320
rect 122170 669970 122190 670210
rect 122430 669970 122520 670210
rect 122760 669970 122850 670210
rect 123090 669970 123180 670210
rect 123420 669970 123530 670210
rect 123770 669970 123860 670210
rect 124100 669970 124190 670210
rect 124430 669970 124520 670210
rect 124760 669970 124870 670210
rect 125110 669970 125200 670210
rect 125440 669970 125530 670210
rect 125770 669970 125860 670210
rect 126100 669970 126210 670210
rect 126450 669970 126540 670210
rect 126780 669970 126870 670210
rect 127110 669970 127200 670210
rect 127440 669970 127550 670210
rect 127790 669970 127880 670210
rect 128120 669970 128210 670210
rect 128450 669970 128540 670210
rect 128780 669970 128890 670210
rect 129130 669970 129220 670210
rect 129460 669970 129550 670210
rect 129790 669970 129880 670210
rect 130120 669970 130230 670210
rect 130470 669970 130560 670210
rect 130800 669970 130890 670210
rect 131130 669970 131220 670210
rect 131460 669970 131570 670210
rect 131810 669970 131900 670210
rect 132140 669970 132230 670210
rect 132470 669970 132560 670210
rect 132800 669970 132910 670210
rect 133150 669970 133170 670210
rect 122170 669880 133170 669970
rect 122170 669640 122190 669880
rect 122430 669640 122520 669880
rect 122760 669640 122850 669880
rect 123090 669640 123180 669880
rect 123420 669640 123530 669880
rect 123770 669640 123860 669880
rect 124100 669640 124190 669880
rect 124430 669640 124520 669880
rect 124760 669640 124870 669880
rect 125110 669640 125200 669880
rect 125440 669640 125530 669880
rect 125770 669640 125860 669880
rect 126100 669640 126210 669880
rect 126450 669640 126540 669880
rect 126780 669640 126870 669880
rect 127110 669640 127200 669880
rect 127440 669640 127550 669880
rect 127790 669640 127880 669880
rect 128120 669640 128210 669880
rect 128450 669640 128540 669880
rect 128780 669640 128890 669880
rect 129130 669640 129220 669880
rect 129460 669640 129550 669880
rect 129790 669640 129880 669880
rect 130120 669640 130230 669880
rect 130470 669640 130560 669880
rect 130800 669640 130890 669880
rect 131130 669640 131220 669880
rect 131460 669640 131570 669880
rect 131810 669640 131900 669880
rect 132140 669640 132230 669880
rect 132470 669640 132560 669880
rect 132800 669640 132910 669880
rect 133150 669640 133170 669880
rect 122170 669550 133170 669640
rect 122170 669310 122190 669550
rect 122430 669310 122520 669550
rect 122760 669310 122850 669550
rect 123090 669310 123180 669550
rect 123420 669310 123530 669550
rect 123770 669310 123860 669550
rect 124100 669310 124190 669550
rect 124430 669310 124520 669550
rect 124760 669310 124870 669550
rect 125110 669310 125200 669550
rect 125440 669310 125530 669550
rect 125770 669310 125860 669550
rect 126100 669310 126210 669550
rect 126450 669310 126540 669550
rect 126780 669310 126870 669550
rect 127110 669310 127200 669550
rect 127440 669310 127550 669550
rect 127790 669310 127880 669550
rect 128120 669310 128210 669550
rect 128450 669310 128540 669550
rect 128780 669310 128890 669550
rect 129130 669310 129220 669550
rect 129460 669310 129550 669550
rect 129790 669310 129880 669550
rect 130120 669310 130230 669550
rect 130470 669310 130560 669550
rect 130800 669310 130890 669550
rect 131130 669310 131220 669550
rect 131460 669310 131570 669550
rect 131810 669310 131900 669550
rect 132140 669310 132230 669550
rect 132470 669310 132560 669550
rect 132800 669310 132910 669550
rect 133150 669310 133170 669550
rect 122170 669220 133170 669310
rect 122170 668980 122190 669220
rect 122430 668980 122520 669220
rect 122760 668980 122850 669220
rect 123090 668980 123180 669220
rect 123420 668980 123530 669220
rect 123770 668980 123860 669220
rect 124100 668980 124190 669220
rect 124430 668980 124520 669220
rect 124760 668980 124870 669220
rect 125110 668980 125200 669220
rect 125440 668980 125530 669220
rect 125770 668980 125860 669220
rect 126100 668980 126210 669220
rect 126450 668980 126540 669220
rect 126780 668980 126870 669220
rect 127110 668980 127200 669220
rect 127440 668980 127550 669220
rect 127790 668980 127880 669220
rect 128120 668980 128210 669220
rect 128450 668980 128540 669220
rect 128780 668980 128890 669220
rect 129130 668980 129220 669220
rect 129460 668980 129550 669220
rect 129790 668980 129880 669220
rect 130120 668980 130230 669220
rect 130470 668980 130560 669220
rect 130800 668980 130890 669220
rect 131130 668980 131220 669220
rect 131460 668980 131570 669220
rect 131810 668980 131900 669220
rect 132140 668980 132230 669220
rect 132470 668980 132560 669220
rect 132800 668980 132910 669220
rect 133150 668980 133170 669220
rect 122170 668870 133170 668980
rect 122170 668630 122190 668870
rect 122430 668630 122520 668870
rect 122760 668630 122850 668870
rect 123090 668630 123180 668870
rect 123420 668630 123530 668870
rect 123770 668630 123860 668870
rect 124100 668630 124190 668870
rect 124430 668630 124520 668870
rect 124760 668630 124870 668870
rect 125110 668630 125200 668870
rect 125440 668630 125530 668870
rect 125770 668630 125860 668870
rect 126100 668630 126210 668870
rect 126450 668630 126540 668870
rect 126780 668630 126870 668870
rect 127110 668630 127200 668870
rect 127440 668630 127550 668870
rect 127790 668630 127880 668870
rect 128120 668630 128210 668870
rect 128450 668630 128540 668870
rect 128780 668630 128890 668870
rect 129130 668630 129220 668870
rect 129460 668630 129550 668870
rect 129790 668630 129880 668870
rect 130120 668630 130230 668870
rect 130470 668630 130560 668870
rect 130800 668630 130890 668870
rect 131130 668630 131220 668870
rect 131460 668630 131570 668870
rect 131810 668630 131900 668870
rect 132140 668630 132230 668870
rect 132470 668630 132560 668870
rect 132800 668630 132910 668870
rect 133150 668630 133170 668870
rect 122170 668540 133170 668630
rect 122170 668300 122190 668540
rect 122430 668300 122520 668540
rect 122760 668300 122850 668540
rect 123090 668300 123180 668540
rect 123420 668300 123530 668540
rect 123770 668300 123860 668540
rect 124100 668300 124190 668540
rect 124430 668300 124520 668540
rect 124760 668300 124870 668540
rect 125110 668300 125200 668540
rect 125440 668300 125530 668540
rect 125770 668300 125860 668540
rect 126100 668300 126210 668540
rect 126450 668300 126540 668540
rect 126780 668300 126870 668540
rect 127110 668300 127200 668540
rect 127440 668300 127550 668540
rect 127790 668300 127880 668540
rect 128120 668300 128210 668540
rect 128450 668300 128540 668540
rect 128780 668300 128890 668540
rect 129130 668300 129220 668540
rect 129460 668300 129550 668540
rect 129790 668300 129880 668540
rect 130120 668300 130230 668540
rect 130470 668300 130560 668540
rect 130800 668300 130890 668540
rect 131130 668300 131220 668540
rect 131460 668300 131570 668540
rect 131810 668300 131900 668540
rect 132140 668300 132230 668540
rect 132470 668300 132560 668540
rect 132800 668300 132910 668540
rect 133150 668300 133170 668540
rect 122170 668210 133170 668300
rect 122170 667970 122190 668210
rect 122430 667970 122520 668210
rect 122760 667970 122850 668210
rect 123090 667970 123180 668210
rect 123420 667970 123530 668210
rect 123770 667970 123860 668210
rect 124100 667970 124190 668210
rect 124430 667970 124520 668210
rect 124760 667970 124870 668210
rect 125110 667970 125200 668210
rect 125440 667970 125530 668210
rect 125770 667970 125860 668210
rect 126100 667970 126210 668210
rect 126450 667970 126540 668210
rect 126780 667970 126870 668210
rect 127110 667970 127200 668210
rect 127440 667970 127550 668210
rect 127790 667970 127880 668210
rect 128120 667970 128210 668210
rect 128450 667970 128540 668210
rect 128780 667970 128890 668210
rect 129130 667970 129220 668210
rect 129460 667970 129550 668210
rect 129790 667970 129880 668210
rect 130120 667970 130230 668210
rect 130470 667970 130560 668210
rect 130800 667970 130890 668210
rect 131130 667970 131220 668210
rect 131460 667970 131570 668210
rect 131810 667970 131900 668210
rect 132140 667970 132230 668210
rect 132470 667970 132560 668210
rect 132800 667970 132910 668210
rect 133150 667970 133170 668210
rect 122170 667880 133170 667970
rect 122170 667640 122190 667880
rect 122430 667640 122520 667880
rect 122760 667640 122850 667880
rect 123090 667640 123180 667880
rect 123420 667640 123530 667880
rect 123770 667640 123860 667880
rect 124100 667640 124190 667880
rect 124430 667640 124520 667880
rect 124760 667640 124870 667880
rect 125110 667640 125200 667880
rect 125440 667640 125530 667880
rect 125770 667640 125860 667880
rect 126100 667640 126210 667880
rect 126450 667640 126540 667880
rect 126780 667640 126870 667880
rect 127110 667640 127200 667880
rect 127440 667640 127550 667880
rect 127790 667640 127880 667880
rect 128120 667640 128210 667880
rect 128450 667640 128540 667880
rect 128780 667640 128890 667880
rect 129130 667640 129220 667880
rect 129460 667640 129550 667880
rect 129790 667640 129880 667880
rect 130120 667640 130230 667880
rect 130470 667640 130560 667880
rect 130800 667640 130890 667880
rect 131130 667640 131220 667880
rect 131460 667640 131570 667880
rect 131810 667640 131900 667880
rect 132140 667640 132230 667880
rect 132470 667640 132560 667880
rect 132800 667640 132910 667880
rect 133150 667640 133170 667880
rect 122170 667530 133170 667640
rect 122170 667290 122190 667530
rect 122430 667290 122520 667530
rect 122760 667290 122850 667530
rect 123090 667290 123180 667530
rect 123420 667290 123530 667530
rect 123770 667290 123860 667530
rect 124100 667290 124190 667530
rect 124430 667290 124520 667530
rect 124760 667290 124870 667530
rect 125110 667290 125200 667530
rect 125440 667290 125530 667530
rect 125770 667290 125860 667530
rect 126100 667290 126210 667530
rect 126450 667290 126540 667530
rect 126780 667290 126870 667530
rect 127110 667290 127200 667530
rect 127440 667290 127550 667530
rect 127790 667290 127880 667530
rect 128120 667290 128210 667530
rect 128450 667290 128540 667530
rect 128780 667290 128890 667530
rect 129130 667290 129220 667530
rect 129460 667290 129550 667530
rect 129790 667290 129880 667530
rect 130120 667290 130230 667530
rect 130470 667290 130560 667530
rect 130800 667290 130890 667530
rect 131130 667290 131220 667530
rect 131460 667290 131570 667530
rect 131810 667290 131900 667530
rect 132140 667290 132230 667530
rect 132470 667290 132560 667530
rect 132800 667290 132910 667530
rect 133150 667290 133170 667530
rect 122170 667200 133170 667290
rect 122170 666960 122190 667200
rect 122430 666960 122520 667200
rect 122760 666960 122850 667200
rect 123090 666960 123180 667200
rect 123420 666960 123530 667200
rect 123770 666960 123860 667200
rect 124100 666960 124190 667200
rect 124430 666960 124520 667200
rect 124760 666960 124870 667200
rect 125110 666960 125200 667200
rect 125440 666960 125530 667200
rect 125770 666960 125860 667200
rect 126100 666960 126210 667200
rect 126450 666960 126540 667200
rect 126780 666960 126870 667200
rect 127110 666960 127200 667200
rect 127440 666960 127550 667200
rect 127790 666960 127880 667200
rect 128120 666960 128210 667200
rect 128450 666960 128540 667200
rect 128780 666960 128890 667200
rect 129130 666960 129220 667200
rect 129460 666960 129550 667200
rect 129790 666960 129880 667200
rect 130120 666960 130230 667200
rect 130470 666960 130560 667200
rect 130800 666960 130890 667200
rect 131130 666960 131220 667200
rect 131460 666960 131570 667200
rect 131810 666960 131900 667200
rect 132140 666960 132230 667200
rect 132470 666960 132560 667200
rect 132800 666960 132910 667200
rect 133150 666960 133170 667200
rect 122170 666870 133170 666960
rect 122170 666630 122190 666870
rect 122430 666630 122520 666870
rect 122760 666630 122850 666870
rect 123090 666630 123180 666870
rect 123420 666630 123530 666870
rect 123770 666630 123860 666870
rect 124100 666630 124190 666870
rect 124430 666630 124520 666870
rect 124760 666630 124870 666870
rect 125110 666630 125200 666870
rect 125440 666630 125530 666870
rect 125770 666630 125860 666870
rect 126100 666630 126210 666870
rect 126450 666630 126540 666870
rect 126780 666630 126870 666870
rect 127110 666630 127200 666870
rect 127440 666630 127550 666870
rect 127790 666630 127880 666870
rect 128120 666630 128210 666870
rect 128450 666630 128540 666870
rect 128780 666630 128890 666870
rect 129130 666630 129220 666870
rect 129460 666630 129550 666870
rect 129790 666630 129880 666870
rect 130120 666630 130230 666870
rect 130470 666630 130560 666870
rect 130800 666630 130890 666870
rect 131130 666630 131220 666870
rect 131460 666630 131570 666870
rect 131810 666630 131900 666870
rect 132140 666630 132230 666870
rect 132470 666630 132560 666870
rect 132800 666630 132910 666870
rect 133150 666630 133170 666870
rect 122170 666540 133170 666630
rect 122170 666300 122190 666540
rect 122430 666300 122520 666540
rect 122760 666300 122850 666540
rect 123090 666300 123180 666540
rect 123420 666300 123530 666540
rect 123770 666300 123860 666540
rect 124100 666300 124190 666540
rect 124430 666300 124520 666540
rect 124760 666300 124870 666540
rect 125110 666300 125200 666540
rect 125440 666300 125530 666540
rect 125770 666300 125860 666540
rect 126100 666300 126210 666540
rect 126450 666300 126540 666540
rect 126780 666300 126870 666540
rect 127110 666300 127200 666540
rect 127440 666300 127550 666540
rect 127790 666300 127880 666540
rect 128120 666300 128210 666540
rect 128450 666300 128540 666540
rect 128780 666300 128890 666540
rect 129130 666300 129220 666540
rect 129460 666300 129550 666540
rect 129790 666300 129880 666540
rect 130120 666300 130230 666540
rect 130470 666300 130560 666540
rect 130800 666300 130890 666540
rect 131130 666300 131220 666540
rect 131460 666300 131570 666540
rect 131810 666300 131900 666540
rect 132140 666300 132230 666540
rect 132470 666300 132560 666540
rect 132800 666300 132910 666540
rect 133150 666300 133170 666540
rect 122170 666190 133170 666300
rect 122170 665950 122190 666190
rect 122430 665950 122520 666190
rect 122760 665950 122850 666190
rect 123090 665950 123180 666190
rect 123420 665950 123530 666190
rect 123770 665950 123860 666190
rect 124100 665950 124190 666190
rect 124430 665950 124520 666190
rect 124760 665950 124870 666190
rect 125110 665950 125200 666190
rect 125440 665950 125530 666190
rect 125770 665950 125860 666190
rect 126100 665950 126210 666190
rect 126450 665950 126540 666190
rect 126780 665950 126870 666190
rect 127110 665950 127200 666190
rect 127440 665950 127550 666190
rect 127790 665950 127880 666190
rect 128120 665950 128210 666190
rect 128450 665950 128540 666190
rect 128780 665950 128890 666190
rect 129130 665950 129220 666190
rect 129460 665950 129550 666190
rect 129790 665950 129880 666190
rect 130120 665950 130230 666190
rect 130470 665950 130560 666190
rect 130800 665950 130890 666190
rect 131130 665950 131220 666190
rect 131460 665950 131570 666190
rect 131810 665950 131900 666190
rect 132140 665950 132230 666190
rect 132470 665950 132560 666190
rect 132800 665950 132910 666190
rect 133150 665950 133170 666190
rect 122170 665860 133170 665950
rect 122170 665620 122190 665860
rect 122430 665620 122520 665860
rect 122760 665620 122850 665860
rect 123090 665620 123180 665860
rect 123420 665620 123530 665860
rect 123770 665620 123860 665860
rect 124100 665620 124190 665860
rect 124430 665620 124520 665860
rect 124760 665620 124870 665860
rect 125110 665620 125200 665860
rect 125440 665620 125530 665860
rect 125770 665620 125860 665860
rect 126100 665620 126210 665860
rect 126450 665620 126540 665860
rect 126780 665620 126870 665860
rect 127110 665620 127200 665860
rect 127440 665620 127550 665860
rect 127790 665620 127880 665860
rect 128120 665620 128210 665860
rect 128450 665620 128540 665860
rect 128780 665620 128890 665860
rect 129130 665620 129220 665860
rect 129460 665620 129550 665860
rect 129790 665620 129880 665860
rect 130120 665620 130230 665860
rect 130470 665620 130560 665860
rect 130800 665620 130890 665860
rect 131130 665620 131220 665860
rect 131460 665620 131570 665860
rect 131810 665620 131900 665860
rect 132140 665620 132230 665860
rect 132470 665620 132560 665860
rect 132800 665620 132910 665860
rect 133150 665620 133170 665860
rect 122170 665530 133170 665620
rect 122170 665290 122190 665530
rect 122430 665290 122520 665530
rect 122760 665290 122850 665530
rect 123090 665290 123180 665530
rect 123420 665290 123530 665530
rect 123770 665290 123860 665530
rect 124100 665290 124190 665530
rect 124430 665290 124520 665530
rect 124760 665290 124870 665530
rect 125110 665290 125200 665530
rect 125440 665290 125530 665530
rect 125770 665290 125860 665530
rect 126100 665290 126210 665530
rect 126450 665290 126540 665530
rect 126780 665290 126870 665530
rect 127110 665290 127200 665530
rect 127440 665290 127550 665530
rect 127790 665290 127880 665530
rect 128120 665290 128210 665530
rect 128450 665290 128540 665530
rect 128780 665290 128890 665530
rect 129130 665290 129220 665530
rect 129460 665290 129550 665530
rect 129790 665290 129880 665530
rect 130120 665290 130230 665530
rect 130470 665290 130560 665530
rect 130800 665290 130890 665530
rect 131130 665290 131220 665530
rect 131460 665290 131570 665530
rect 131810 665290 131900 665530
rect 132140 665290 132230 665530
rect 132470 665290 132560 665530
rect 132800 665290 132910 665530
rect 133150 665290 133170 665530
rect 122170 665200 133170 665290
rect 122170 664960 122190 665200
rect 122430 664960 122520 665200
rect 122760 664960 122850 665200
rect 123090 664960 123180 665200
rect 123420 664960 123530 665200
rect 123770 664960 123860 665200
rect 124100 664960 124190 665200
rect 124430 664960 124520 665200
rect 124760 664960 124870 665200
rect 125110 664960 125200 665200
rect 125440 664960 125530 665200
rect 125770 664960 125860 665200
rect 126100 664960 126210 665200
rect 126450 664960 126540 665200
rect 126780 664960 126870 665200
rect 127110 664960 127200 665200
rect 127440 664960 127550 665200
rect 127790 664960 127880 665200
rect 128120 664960 128210 665200
rect 128450 664960 128540 665200
rect 128780 664960 128890 665200
rect 129130 664960 129220 665200
rect 129460 664960 129550 665200
rect 129790 664960 129880 665200
rect 130120 664960 130230 665200
rect 130470 664960 130560 665200
rect 130800 664960 130890 665200
rect 131130 664960 131220 665200
rect 131460 664960 131570 665200
rect 131810 664960 131900 665200
rect 132140 664960 132230 665200
rect 132470 664960 132560 665200
rect 132800 664960 132910 665200
rect 133150 664960 133170 665200
rect 122170 664850 133170 664960
rect 122170 664610 122190 664850
rect 122430 664610 122520 664850
rect 122760 664610 122850 664850
rect 123090 664610 123180 664850
rect 123420 664610 123530 664850
rect 123770 664610 123860 664850
rect 124100 664610 124190 664850
rect 124430 664610 124520 664850
rect 124760 664610 124870 664850
rect 125110 664610 125200 664850
rect 125440 664610 125530 664850
rect 125770 664610 125860 664850
rect 126100 664610 126210 664850
rect 126450 664610 126540 664850
rect 126780 664610 126870 664850
rect 127110 664610 127200 664850
rect 127440 664610 127550 664850
rect 127790 664610 127880 664850
rect 128120 664610 128210 664850
rect 128450 664610 128540 664850
rect 128780 664610 128890 664850
rect 129130 664610 129220 664850
rect 129460 664610 129550 664850
rect 129790 664610 129880 664850
rect 130120 664610 130230 664850
rect 130470 664610 130560 664850
rect 130800 664610 130890 664850
rect 131130 664610 131220 664850
rect 131460 664610 131570 664850
rect 131810 664610 131900 664850
rect 132140 664610 132230 664850
rect 132470 664610 132560 664850
rect 132800 664610 132910 664850
rect 133150 664610 133170 664850
rect 122170 664520 133170 664610
rect 122170 664280 122190 664520
rect 122430 664280 122520 664520
rect 122760 664280 122850 664520
rect 123090 664280 123180 664520
rect 123420 664280 123530 664520
rect 123770 664280 123860 664520
rect 124100 664280 124190 664520
rect 124430 664280 124520 664520
rect 124760 664280 124870 664520
rect 125110 664280 125200 664520
rect 125440 664280 125530 664520
rect 125770 664280 125860 664520
rect 126100 664280 126210 664520
rect 126450 664280 126540 664520
rect 126780 664280 126870 664520
rect 127110 664280 127200 664520
rect 127440 664280 127550 664520
rect 127790 664280 127880 664520
rect 128120 664280 128210 664520
rect 128450 664280 128540 664520
rect 128780 664280 128890 664520
rect 129130 664280 129220 664520
rect 129460 664280 129550 664520
rect 129790 664280 129880 664520
rect 130120 664280 130230 664520
rect 130470 664280 130560 664520
rect 130800 664280 130890 664520
rect 131130 664280 131220 664520
rect 131460 664280 131570 664520
rect 131810 664280 131900 664520
rect 132140 664280 132230 664520
rect 132470 664280 132560 664520
rect 132800 664280 132910 664520
rect 133150 664280 133170 664520
rect 122170 664190 133170 664280
rect 122170 663950 122190 664190
rect 122430 663950 122520 664190
rect 122760 663950 122850 664190
rect 123090 663950 123180 664190
rect 123420 663950 123530 664190
rect 123770 663950 123860 664190
rect 124100 663950 124190 664190
rect 124430 663950 124520 664190
rect 124760 663950 124870 664190
rect 125110 663950 125200 664190
rect 125440 663950 125530 664190
rect 125770 663950 125860 664190
rect 126100 663950 126210 664190
rect 126450 663950 126540 664190
rect 126780 663950 126870 664190
rect 127110 663950 127200 664190
rect 127440 663950 127550 664190
rect 127790 663950 127880 664190
rect 128120 663950 128210 664190
rect 128450 663950 128540 664190
rect 128780 663950 128890 664190
rect 129130 663950 129220 664190
rect 129460 663950 129550 664190
rect 129790 663950 129880 664190
rect 130120 663950 130230 664190
rect 130470 663950 130560 664190
rect 130800 663950 130890 664190
rect 131130 663950 131220 664190
rect 131460 663950 131570 664190
rect 131810 663950 131900 664190
rect 132140 663950 132230 664190
rect 132470 663950 132560 664190
rect 132800 663950 132910 664190
rect 133150 663950 133170 664190
rect 122170 663860 133170 663950
rect 122170 663620 122190 663860
rect 122430 663620 122520 663860
rect 122760 663620 122850 663860
rect 123090 663620 123180 663860
rect 123420 663620 123530 663860
rect 123770 663620 123860 663860
rect 124100 663620 124190 663860
rect 124430 663620 124520 663860
rect 124760 663620 124870 663860
rect 125110 663620 125200 663860
rect 125440 663620 125530 663860
rect 125770 663620 125860 663860
rect 126100 663620 126210 663860
rect 126450 663620 126540 663860
rect 126780 663620 126870 663860
rect 127110 663620 127200 663860
rect 127440 663620 127550 663860
rect 127790 663620 127880 663860
rect 128120 663620 128210 663860
rect 128450 663620 128540 663860
rect 128780 663620 128890 663860
rect 129130 663620 129220 663860
rect 129460 663620 129550 663860
rect 129790 663620 129880 663860
rect 130120 663620 130230 663860
rect 130470 663620 130560 663860
rect 130800 663620 130890 663860
rect 131130 663620 131220 663860
rect 131460 663620 131570 663860
rect 131810 663620 131900 663860
rect 132140 663620 132230 663860
rect 132470 663620 132560 663860
rect 132800 663620 132910 663860
rect 133150 663620 133170 663860
rect 122170 663510 133170 663620
rect 122170 663270 122190 663510
rect 122430 663270 122520 663510
rect 122760 663270 122850 663510
rect 123090 663270 123180 663510
rect 123420 663270 123530 663510
rect 123770 663270 123860 663510
rect 124100 663270 124190 663510
rect 124430 663270 124520 663510
rect 124760 663270 124870 663510
rect 125110 663270 125200 663510
rect 125440 663270 125530 663510
rect 125770 663270 125860 663510
rect 126100 663270 126210 663510
rect 126450 663270 126540 663510
rect 126780 663270 126870 663510
rect 127110 663270 127200 663510
rect 127440 663270 127550 663510
rect 127790 663270 127880 663510
rect 128120 663270 128210 663510
rect 128450 663270 128540 663510
rect 128780 663270 128890 663510
rect 129130 663270 129220 663510
rect 129460 663270 129550 663510
rect 129790 663270 129880 663510
rect 130120 663270 130230 663510
rect 130470 663270 130560 663510
rect 130800 663270 130890 663510
rect 131130 663270 131220 663510
rect 131460 663270 131570 663510
rect 131810 663270 131900 663510
rect 132140 663270 132230 663510
rect 132470 663270 132560 663510
rect 132800 663270 132910 663510
rect 133150 663270 133170 663510
rect 122170 663180 133170 663270
rect 122170 662940 122190 663180
rect 122430 662940 122520 663180
rect 122760 662940 122850 663180
rect 123090 662940 123180 663180
rect 123420 662940 123530 663180
rect 123770 662940 123860 663180
rect 124100 662940 124190 663180
rect 124430 662940 124520 663180
rect 124760 662940 124870 663180
rect 125110 662940 125200 663180
rect 125440 662940 125530 663180
rect 125770 662940 125860 663180
rect 126100 662940 126210 663180
rect 126450 662940 126540 663180
rect 126780 662940 126870 663180
rect 127110 662940 127200 663180
rect 127440 662940 127550 663180
rect 127790 662940 127880 663180
rect 128120 662940 128210 663180
rect 128450 662940 128540 663180
rect 128780 662940 128890 663180
rect 129130 662940 129220 663180
rect 129460 662940 129550 663180
rect 129790 662940 129880 663180
rect 130120 662940 130230 663180
rect 130470 662940 130560 663180
rect 130800 662940 130890 663180
rect 131130 662940 131220 663180
rect 131460 662940 131570 663180
rect 131810 662940 131900 663180
rect 132140 662940 132230 663180
rect 132470 662940 132560 663180
rect 132800 662940 132910 663180
rect 133150 662940 133170 663180
rect 122170 662850 133170 662940
rect 122170 662610 122190 662850
rect 122430 662610 122520 662850
rect 122760 662610 122850 662850
rect 123090 662610 123180 662850
rect 123420 662610 123530 662850
rect 123770 662610 123860 662850
rect 124100 662610 124190 662850
rect 124430 662610 124520 662850
rect 124760 662610 124870 662850
rect 125110 662610 125200 662850
rect 125440 662610 125530 662850
rect 125770 662610 125860 662850
rect 126100 662610 126210 662850
rect 126450 662610 126540 662850
rect 126780 662610 126870 662850
rect 127110 662610 127200 662850
rect 127440 662610 127550 662850
rect 127790 662610 127880 662850
rect 128120 662610 128210 662850
rect 128450 662610 128540 662850
rect 128780 662610 128890 662850
rect 129130 662610 129220 662850
rect 129460 662610 129550 662850
rect 129790 662610 129880 662850
rect 130120 662610 130230 662850
rect 130470 662610 130560 662850
rect 130800 662610 130890 662850
rect 131130 662610 131220 662850
rect 131460 662610 131570 662850
rect 131810 662610 131900 662850
rect 132140 662610 132230 662850
rect 132470 662610 132560 662850
rect 132800 662610 132910 662850
rect 133150 662610 133170 662850
rect 122170 662520 133170 662610
rect 122170 662280 122190 662520
rect 122430 662280 122520 662520
rect 122760 662280 122850 662520
rect 123090 662280 123180 662520
rect 123420 662280 123530 662520
rect 123770 662280 123860 662520
rect 124100 662280 124190 662520
rect 124430 662280 124520 662520
rect 124760 662280 124870 662520
rect 125110 662280 125200 662520
rect 125440 662280 125530 662520
rect 125770 662280 125860 662520
rect 126100 662280 126210 662520
rect 126450 662280 126540 662520
rect 126780 662280 126870 662520
rect 127110 662280 127200 662520
rect 127440 662280 127550 662520
rect 127790 662280 127880 662520
rect 128120 662280 128210 662520
rect 128450 662280 128540 662520
rect 128780 662280 128890 662520
rect 129130 662280 129220 662520
rect 129460 662280 129550 662520
rect 129790 662280 129880 662520
rect 130120 662280 130230 662520
rect 130470 662280 130560 662520
rect 130800 662280 130890 662520
rect 131130 662280 131220 662520
rect 131460 662280 131570 662520
rect 131810 662280 131900 662520
rect 132140 662280 132230 662520
rect 132470 662280 132560 662520
rect 132800 662280 132910 662520
rect 133150 662280 133170 662520
rect 122170 662170 133170 662280
rect 122170 661930 122190 662170
rect 122430 661930 122520 662170
rect 122760 661930 122850 662170
rect 123090 661930 123180 662170
rect 123420 661930 123530 662170
rect 123770 661930 123860 662170
rect 124100 661930 124190 662170
rect 124430 661930 124520 662170
rect 124760 661930 124870 662170
rect 125110 661930 125200 662170
rect 125440 661930 125530 662170
rect 125770 661930 125860 662170
rect 126100 661930 126210 662170
rect 126450 661930 126540 662170
rect 126780 661930 126870 662170
rect 127110 661930 127200 662170
rect 127440 661930 127550 662170
rect 127790 661930 127880 662170
rect 128120 661930 128210 662170
rect 128450 661930 128540 662170
rect 128780 661930 128890 662170
rect 129130 661930 129220 662170
rect 129460 661930 129550 662170
rect 129790 661930 129880 662170
rect 130120 661930 130230 662170
rect 130470 661930 130560 662170
rect 130800 661930 130890 662170
rect 131130 661930 131220 662170
rect 131460 661930 131570 662170
rect 131810 661930 131900 662170
rect 132140 661930 132230 662170
rect 132470 661930 132560 662170
rect 132800 661930 132910 662170
rect 133150 661930 133170 662170
rect 122170 661840 133170 661930
rect 122170 661600 122190 661840
rect 122430 661600 122520 661840
rect 122760 661600 122850 661840
rect 123090 661600 123180 661840
rect 123420 661600 123530 661840
rect 123770 661600 123860 661840
rect 124100 661600 124190 661840
rect 124430 661600 124520 661840
rect 124760 661600 124870 661840
rect 125110 661600 125200 661840
rect 125440 661600 125530 661840
rect 125770 661600 125860 661840
rect 126100 661600 126210 661840
rect 126450 661600 126540 661840
rect 126780 661600 126870 661840
rect 127110 661600 127200 661840
rect 127440 661600 127550 661840
rect 127790 661600 127880 661840
rect 128120 661600 128210 661840
rect 128450 661600 128540 661840
rect 128780 661600 128890 661840
rect 129130 661600 129220 661840
rect 129460 661600 129550 661840
rect 129790 661600 129880 661840
rect 130120 661600 130230 661840
rect 130470 661600 130560 661840
rect 130800 661600 130890 661840
rect 131130 661600 131220 661840
rect 131460 661600 131570 661840
rect 131810 661600 131900 661840
rect 132140 661600 132230 661840
rect 132470 661600 132560 661840
rect 132800 661600 132910 661840
rect 133150 661600 133170 661840
rect 122170 661510 133170 661600
rect 122170 661270 122190 661510
rect 122430 661270 122520 661510
rect 122760 661270 122850 661510
rect 123090 661270 123180 661510
rect 123420 661270 123530 661510
rect 123770 661270 123860 661510
rect 124100 661270 124190 661510
rect 124430 661270 124520 661510
rect 124760 661270 124870 661510
rect 125110 661270 125200 661510
rect 125440 661270 125530 661510
rect 125770 661270 125860 661510
rect 126100 661270 126210 661510
rect 126450 661270 126540 661510
rect 126780 661270 126870 661510
rect 127110 661270 127200 661510
rect 127440 661270 127550 661510
rect 127790 661270 127880 661510
rect 128120 661270 128210 661510
rect 128450 661270 128540 661510
rect 128780 661270 128890 661510
rect 129130 661270 129220 661510
rect 129460 661270 129550 661510
rect 129790 661270 129880 661510
rect 130120 661270 130230 661510
rect 130470 661270 130560 661510
rect 130800 661270 130890 661510
rect 131130 661270 131220 661510
rect 131460 661270 131570 661510
rect 131810 661270 131900 661510
rect 132140 661270 132230 661510
rect 132470 661270 132560 661510
rect 132800 661270 132910 661510
rect 133150 661270 133170 661510
rect 122170 661180 133170 661270
rect 122170 660940 122190 661180
rect 122430 660940 122520 661180
rect 122760 660940 122850 661180
rect 123090 660940 123180 661180
rect 123420 660940 123530 661180
rect 123770 660940 123860 661180
rect 124100 660940 124190 661180
rect 124430 660940 124520 661180
rect 124760 660940 124870 661180
rect 125110 660940 125200 661180
rect 125440 660940 125530 661180
rect 125770 660940 125860 661180
rect 126100 660940 126210 661180
rect 126450 660940 126540 661180
rect 126780 660940 126870 661180
rect 127110 660940 127200 661180
rect 127440 660940 127550 661180
rect 127790 660940 127880 661180
rect 128120 660940 128210 661180
rect 128450 660940 128540 661180
rect 128780 660940 128890 661180
rect 129130 660940 129220 661180
rect 129460 660940 129550 661180
rect 129790 660940 129880 661180
rect 130120 660940 130230 661180
rect 130470 660940 130560 661180
rect 130800 660940 130890 661180
rect 131130 660940 131220 661180
rect 131460 660940 131570 661180
rect 131810 660940 131900 661180
rect 132140 660940 132230 661180
rect 132470 660940 132560 661180
rect 132800 660940 132910 661180
rect 133150 660940 133170 661180
rect 122170 660920 133170 660940
rect 133550 671900 144550 671920
rect 133550 671660 133570 671900
rect 133810 671660 133900 671900
rect 134140 671660 134230 671900
rect 134470 671660 134560 671900
rect 134800 671660 134910 671900
rect 135150 671660 135240 671900
rect 135480 671660 135570 671900
rect 135810 671660 135900 671900
rect 136140 671660 136250 671900
rect 136490 671660 136580 671900
rect 136820 671660 136910 671900
rect 137150 671660 137240 671900
rect 137480 671660 137590 671900
rect 137830 671660 137920 671900
rect 138160 671660 138250 671900
rect 138490 671660 138580 671900
rect 138820 671660 138930 671900
rect 139170 671660 139260 671900
rect 139500 671660 139590 671900
rect 139830 671660 139920 671900
rect 140160 671660 140270 671900
rect 140510 671660 140600 671900
rect 140840 671660 140930 671900
rect 141170 671660 141260 671900
rect 141500 671660 141610 671900
rect 141850 671660 141940 671900
rect 142180 671660 142270 671900
rect 142510 671660 142600 671900
rect 142840 671660 142950 671900
rect 143190 671660 143280 671900
rect 143520 671660 143610 671900
rect 143850 671660 143940 671900
rect 144180 671660 144290 671900
rect 144530 671660 144550 671900
rect 133550 671550 144550 671660
rect 133550 671310 133570 671550
rect 133810 671310 133900 671550
rect 134140 671310 134230 671550
rect 134470 671310 134560 671550
rect 134800 671310 134910 671550
rect 135150 671310 135240 671550
rect 135480 671310 135570 671550
rect 135810 671310 135900 671550
rect 136140 671310 136250 671550
rect 136490 671310 136580 671550
rect 136820 671310 136910 671550
rect 137150 671310 137240 671550
rect 137480 671310 137590 671550
rect 137830 671310 137920 671550
rect 138160 671310 138250 671550
rect 138490 671310 138580 671550
rect 138820 671310 138930 671550
rect 139170 671310 139260 671550
rect 139500 671310 139590 671550
rect 139830 671310 139920 671550
rect 140160 671310 140270 671550
rect 140510 671310 140600 671550
rect 140840 671310 140930 671550
rect 141170 671310 141260 671550
rect 141500 671310 141610 671550
rect 141850 671310 141940 671550
rect 142180 671310 142270 671550
rect 142510 671310 142600 671550
rect 142840 671310 142950 671550
rect 143190 671310 143280 671550
rect 143520 671310 143610 671550
rect 143850 671310 143940 671550
rect 144180 671310 144290 671550
rect 144530 671310 144550 671550
rect 133550 671220 144550 671310
rect 133550 670980 133570 671220
rect 133810 670980 133900 671220
rect 134140 670980 134230 671220
rect 134470 670980 134560 671220
rect 134800 670980 134910 671220
rect 135150 670980 135240 671220
rect 135480 670980 135570 671220
rect 135810 670980 135900 671220
rect 136140 670980 136250 671220
rect 136490 670980 136580 671220
rect 136820 670980 136910 671220
rect 137150 670980 137240 671220
rect 137480 670980 137590 671220
rect 137830 670980 137920 671220
rect 138160 670980 138250 671220
rect 138490 670980 138580 671220
rect 138820 670980 138930 671220
rect 139170 670980 139260 671220
rect 139500 670980 139590 671220
rect 139830 670980 139920 671220
rect 140160 670980 140270 671220
rect 140510 670980 140600 671220
rect 140840 670980 140930 671220
rect 141170 670980 141260 671220
rect 141500 670980 141610 671220
rect 141850 670980 141940 671220
rect 142180 670980 142270 671220
rect 142510 670980 142600 671220
rect 142840 670980 142950 671220
rect 143190 670980 143280 671220
rect 143520 670980 143610 671220
rect 143850 670980 143940 671220
rect 144180 670980 144290 671220
rect 144530 670980 144550 671220
rect 133550 670890 144550 670980
rect 133550 670650 133570 670890
rect 133810 670650 133900 670890
rect 134140 670650 134230 670890
rect 134470 670650 134560 670890
rect 134800 670650 134910 670890
rect 135150 670650 135240 670890
rect 135480 670650 135570 670890
rect 135810 670650 135900 670890
rect 136140 670650 136250 670890
rect 136490 670650 136580 670890
rect 136820 670650 136910 670890
rect 137150 670650 137240 670890
rect 137480 670650 137590 670890
rect 137830 670650 137920 670890
rect 138160 670650 138250 670890
rect 138490 670650 138580 670890
rect 138820 670650 138930 670890
rect 139170 670650 139260 670890
rect 139500 670650 139590 670890
rect 139830 670650 139920 670890
rect 140160 670650 140270 670890
rect 140510 670650 140600 670890
rect 140840 670650 140930 670890
rect 141170 670650 141260 670890
rect 141500 670650 141610 670890
rect 141850 670650 141940 670890
rect 142180 670650 142270 670890
rect 142510 670650 142600 670890
rect 142840 670650 142950 670890
rect 143190 670650 143280 670890
rect 143520 670650 143610 670890
rect 143850 670650 143940 670890
rect 144180 670650 144290 670890
rect 144530 670650 144550 670890
rect 133550 670560 144550 670650
rect 133550 670320 133570 670560
rect 133810 670320 133900 670560
rect 134140 670320 134230 670560
rect 134470 670320 134560 670560
rect 134800 670320 134910 670560
rect 135150 670320 135240 670560
rect 135480 670320 135570 670560
rect 135810 670320 135900 670560
rect 136140 670320 136250 670560
rect 136490 670320 136580 670560
rect 136820 670320 136910 670560
rect 137150 670320 137240 670560
rect 137480 670320 137590 670560
rect 137830 670320 137920 670560
rect 138160 670320 138250 670560
rect 138490 670320 138580 670560
rect 138820 670320 138930 670560
rect 139170 670320 139260 670560
rect 139500 670320 139590 670560
rect 139830 670320 139920 670560
rect 140160 670320 140270 670560
rect 140510 670320 140600 670560
rect 140840 670320 140930 670560
rect 141170 670320 141260 670560
rect 141500 670320 141610 670560
rect 141850 670320 141940 670560
rect 142180 670320 142270 670560
rect 142510 670320 142600 670560
rect 142840 670320 142950 670560
rect 143190 670320 143280 670560
rect 143520 670320 143610 670560
rect 143850 670320 143940 670560
rect 144180 670320 144290 670560
rect 144530 670320 144550 670560
rect 133550 670210 144550 670320
rect 133550 669970 133570 670210
rect 133810 669970 133900 670210
rect 134140 669970 134230 670210
rect 134470 669970 134560 670210
rect 134800 669970 134910 670210
rect 135150 669970 135240 670210
rect 135480 669970 135570 670210
rect 135810 669970 135900 670210
rect 136140 669970 136250 670210
rect 136490 669970 136580 670210
rect 136820 669970 136910 670210
rect 137150 669970 137240 670210
rect 137480 669970 137590 670210
rect 137830 669970 137920 670210
rect 138160 669970 138250 670210
rect 138490 669970 138580 670210
rect 138820 669970 138930 670210
rect 139170 669970 139260 670210
rect 139500 669970 139590 670210
rect 139830 669970 139920 670210
rect 140160 669970 140270 670210
rect 140510 669970 140600 670210
rect 140840 669970 140930 670210
rect 141170 669970 141260 670210
rect 141500 669970 141610 670210
rect 141850 669970 141940 670210
rect 142180 669970 142270 670210
rect 142510 669970 142600 670210
rect 142840 669970 142950 670210
rect 143190 669970 143280 670210
rect 143520 669970 143610 670210
rect 143850 669970 143940 670210
rect 144180 669970 144290 670210
rect 144530 669970 144550 670210
rect 133550 669880 144550 669970
rect 133550 669640 133570 669880
rect 133810 669640 133900 669880
rect 134140 669640 134230 669880
rect 134470 669640 134560 669880
rect 134800 669640 134910 669880
rect 135150 669640 135240 669880
rect 135480 669640 135570 669880
rect 135810 669640 135900 669880
rect 136140 669640 136250 669880
rect 136490 669640 136580 669880
rect 136820 669640 136910 669880
rect 137150 669640 137240 669880
rect 137480 669640 137590 669880
rect 137830 669640 137920 669880
rect 138160 669640 138250 669880
rect 138490 669640 138580 669880
rect 138820 669640 138930 669880
rect 139170 669640 139260 669880
rect 139500 669640 139590 669880
rect 139830 669640 139920 669880
rect 140160 669640 140270 669880
rect 140510 669640 140600 669880
rect 140840 669640 140930 669880
rect 141170 669640 141260 669880
rect 141500 669640 141610 669880
rect 141850 669640 141940 669880
rect 142180 669640 142270 669880
rect 142510 669640 142600 669880
rect 142840 669640 142950 669880
rect 143190 669640 143280 669880
rect 143520 669640 143610 669880
rect 143850 669640 143940 669880
rect 144180 669640 144290 669880
rect 144530 669640 144550 669880
rect 133550 669550 144550 669640
rect 133550 669310 133570 669550
rect 133810 669310 133900 669550
rect 134140 669310 134230 669550
rect 134470 669310 134560 669550
rect 134800 669310 134910 669550
rect 135150 669310 135240 669550
rect 135480 669310 135570 669550
rect 135810 669310 135900 669550
rect 136140 669310 136250 669550
rect 136490 669310 136580 669550
rect 136820 669310 136910 669550
rect 137150 669310 137240 669550
rect 137480 669310 137590 669550
rect 137830 669310 137920 669550
rect 138160 669310 138250 669550
rect 138490 669310 138580 669550
rect 138820 669310 138930 669550
rect 139170 669310 139260 669550
rect 139500 669310 139590 669550
rect 139830 669310 139920 669550
rect 140160 669310 140270 669550
rect 140510 669310 140600 669550
rect 140840 669310 140930 669550
rect 141170 669310 141260 669550
rect 141500 669310 141610 669550
rect 141850 669310 141940 669550
rect 142180 669310 142270 669550
rect 142510 669310 142600 669550
rect 142840 669310 142950 669550
rect 143190 669310 143280 669550
rect 143520 669310 143610 669550
rect 143850 669310 143940 669550
rect 144180 669310 144290 669550
rect 144530 669310 144550 669550
rect 133550 669220 144550 669310
rect 133550 668980 133570 669220
rect 133810 668980 133900 669220
rect 134140 668980 134230 669220
rect 134470 668980 134560 669220
rect 134800 668980 134910 669220
rect 135150 668980 135240 669220
rect 135480 668980 135570 669220
rect 135810 668980 135900 669220
rect 136140 668980 136250 669220
rect 136490 668980 136580 669220
rect 136820 668980 136910 669220
rect 137150 668980 137240 669220
rect 137480 668980 137590 669220
rect 137830 668980 137920 669220
rect 138160 668980 138250 669220
rect 138490 668980 138580 669220
rect 138820 668980 138930 669220
rect 139170 668980 139260 669220
rect 139500 668980 139590 669220
rect 139830 668980 139920 669220
rect 140160 668980 140270 669220
rect 140510 668980 140600 669220
rect 140840 668980 140930 669220
rect 141170 668980 141260 669220
rect 141500 668980 141610 669220
rect 141850 668980 141940 669220
rect 142180 668980 142270 669220
rect 142510 668980 142600 669220
rect 142840 668980 142950 669220
rect 143190 668980 143280 669220
rect 143520 668980 143610 669220
rect 143850 668980 143940 669220
rect 144180 668980 144290 669220
rect 144530 668980 144550 669220
rect 133550 668870 144550 668980
rect 133550 668630 133570 668870
rect 133810 668630 133900 668870
rect 134140 668630 134230 668870
rect 134470 668630 134560 668870
rect 134800 668630 134910 668870
rect 135150 668630 135240 668870
rect 135480 668630 135570 668870
rect 135810 668630 135900 668870
rect 136140 668630 136250 668870
rect 136490 668630 136580 668870
rect 136820 668630 136910 668870
rect 137150 668630 137240 668870
rect 137480 668630 137590 668870
rect 137830 668630 137920 668870
rect 138160 668630 138250 668870
rect 138490 668630 138580 668870
rect 138820 668630 138930 668870
rect 139170 668630 139260 668870
rect 139500 668630 139590 668870
rect 139830 668630 139920 668870
rect 140160 668630 140270 668870
rect 140510 668630 140600 668870
rect 140840 668630 140930 668870
rect 141170 668630 141260 668870
rect 141500 668630 141610 668870
rect 141850 668630 141940 668870
rect 142180 668630 142270 668870
rect 142510 668630 142600 668870
rect 142840 668630 142950 668870
rect 143190 668630 143280 668870
rect 143520 668630 143610 668870
rect 143850 668630 143940 668870
rect 144180 668630 144290 668870
rect 144530 668630 144550 668870
rect 133550 668540 144550 668630
rect 133550 668300 133570 668540
rect 133810 668300 133900 668540
rect 134140 668300 134230 668540
rect 134470 668300 134560 668540
rect 134800 668300 134910 668540
rect 135150 668300 135240 668540
rect 135480 668300 135570 668540
rect 135810 668300 135900 668540
rect 136140 668300 136250 668540
rect 136490 668300 136580 668540
rect 136820 668300 136910 668540
rect 137150 668300 137240 668540
rect 137480 668300 137590 668540
rect 137830 668300 137920 668540
rect 138160 668300 138250 668540
rect 138490 668300 138580 668540
rect 138820 668300 138930 668540
rect 139170 668300 139260 668540
rect 139500 668300 139590 668540
rect 139830 668300 139920 668540
rect 140160 668300 140270 668540
rect 140510 668300 140600 668540
rect 140840 668300 140930 668540
rect 141170 668300 141260 668540
rect 141500 668300 141610 668540
rect 141850 668300 141940 668540
rect 142180 668300 142270 668540
rect 142510 668300 142600 668540
rect 142840 668300 142950 668540
rect 143190 668300 143280 668540
rect 143520 668300 143610 668540
rect 143850 668300 143940 668540
rect 144180 668300 144290 668540
rect 144530 668300 144550 668540
rect 133550 668210 144550 668300
rect 133550 667970 133570 668210
rect 133810 667970 133900 668210
rect 134140 667970 134230 668210
rect 134470 667970 134560 668210
rect 134800 667970 134910 668210
rect 135150 667970 135240 668210
rect 135480 667970 135570 668210
rect 135810 667970 135900 668210
rect 136140 667970 136250 668210
rect 136490 667970 136580 668210
rect 136820 667970 136910 668210
rect 137150 667970 137240 668210
rect 137480 667970 137590 668210
rect 137830 667970 137920 668210
rect 138160 667970 138250 668210
rect 138490 667970 138580 668210
rect 138820 667970 138930 668210
rect 139170 667970 139260 668210
rect 139500 667970 139590 668210
rect 139830 667970 139920 668210
rect 140160 667970 140270 668210
rect 140510 667970 140600 668210
rect 140840 667970 140930 668210
rect 141170 667970 141260 668210
rect 141500 667970 141610 668210
rect 141850 667970 141940 668210
rect 142180 667970 142270 668210
rect 142510 667970 142600 668210
rect 142840 667970 142950 668210
rect 143190 667970 143280 668210
rect 143520 667970 143610 668210
rect 143850 667970 143940 668210
rect 144180 667970 144290 668210
rect 144530 667970 144550 668210
rect 133550 667880 144550 667970
rect 133550 667640 133570 667880
rect 133810 667640 133900 667880
rect 134140 667640 134230 667880
rect 134470 667640 134560 667880
rect 134800 667640 134910 667880
rect 135150 667640 135240 667880
rect 135480 667640 135570 667880
rect 135810 667640 135900 667880
rect 136140 667640 136250 667880
rect 136490 667640 136580 667880
rect 136820 667640 136910 667880
rect 137150 667640 137240 667880
rect 137480 667640 137590 667880
rect 137830 667640 137920 667880
rect 138160 667640 138250 667880
rect 138490 667640 138580 667880
rect 138820 667640 138930 667880
rect 139170 667640 139260 667880
rect 139500 667640 139590 667880
rect 139830 667640 139920 667880
rect 140160 667640 140270 667880
rect 140510 667640 140600 667880
rect 140840 667640 140930 667880
rect 141170 667640 141260 667880
rect 141500 667640 141610 667880
rect 141850 667640 141940 667880
rect 142180 667640 142270 667880
rect 142510 667640 142600 667880
rect 142840 667640 142950 667880
rect 143190 667640 143280 667880
rect 143520 667640 143610 667880
rect 143850 667640 143940 667880
rect 144180 667640 144290 667880
rect 144530 667640 144550 667880
rect 133550 667530 144550 667640
rect 133550 667290 133570 667530
rect 133810 667290 133900 667530
rect 134140 667290 134230 667530
rect 134470 667290 134560 667530
rect 134800 667290 134910 667530
rect 135150 667290 135240 667530
rect 135480 667290 135570 667530
rect 135810 667290 135900 667530
rect 136140 667290 136250 667530
rect 136490 667290 136580 667530
rect 136820 667290 136910 667530
rect 137150 667290 137240 667530
rect 137480 667290 137590 667530
rect 137830 667290 137920 667530
rect 138160 667290 138250 667530
rect 138490 667290 138580 667530
rect 138820 667290 138930 667530
rect 139170 667290 139260 667530
rect 139500 667290 139590 667530
rect 139830 667290 139920 667530
rect 140160 667290 140270 667530
rect 140510 667290 140600 667530
rect 140840 667290 140930 667530
rect 141170 667290 141260 667530
rect 141500 667290 141610 667530
rect 141850 667290 141940 667530
rect 142180 667290 142270 667530
rect 142510 667290 142600 667530
rect 142840 667290 142950 667530
rect 143190 667290 143280 667530
rect 143520 667290 143610 667530
rect 143850 667290 143940 667530
rect 144180 667290 144290 667530
rect 144530 667290 144550 667530
rect 133550 667200 144550 667290
rect 133550 666960 133570 667200
rect 133810 666960 133900 667200
rect 134140 666960 134230 667200
rect 134470 666960 134560 667200
rect 134800 666960 134910 667200
rect 135150 666960 135240 667200
rect 135480 666960 135570 667200
rect 135810 666960 135900 667200
rect 136140 666960 136250 667200
rect 136490 666960 136580 667200
rect 136820 666960 136910 667200
rect 137150 666960 137240 667200
rect 137480 666960 137590 667200
rect 137830 666960 137920 667200
rect 138160 666960 138250 667200
rect 138490 666960 138580 667200
rect 138820 666960 138930 667200
rect 139170 666960 139260 667200
rect 139500 666960 139590 667200
rect 139830 666960 139920 667200
rect 140160 666960 140270 667200
rect 140510 666960 140600 667200
rect 140840 666960 140930 667200
rect 141170 666960 141260 667200
rect 141500 666960 141610 667200
rect 141850 666960 141940 667200
rect 142180 666960 142270 667200
rect 142510 666960 142600 667200
rect 142840 666960 142950 667200
rect 143190 666960 143280 667200
rect 143520 666960 143610 667200
rect 143850 666960 143940 667200
rect 144180 666960 144290 667200
rect 144530 666960 144550 667200
rect 133550 666870 144550 666960
rect 133550 666630 133570 666870
rect 133810 666630 133900 666870
rect 134140 666630 134230 666870
rect 134470 666630 134560 666870
rect 134800 666630 134910 666870
rect 135150 666630 135240 666870
rect 135480 666630 135570 666870
rect 135810 666630 135900 666870
rect 136140 666630 136250 666870
rect 136490 666630 136580 666870
rect 136820 666630 136910 666870
rect 137150 666630 137240 666870
rect 137480 666630 137590 666870
rect 137830 666630 137920 666870
rect 138160 666630 138250 666870
rect 138490 666630 138580 666870
rect 138820 666630 138930 666870
rect 139170 666630 139260 666870
rect 139500 666630 139590 666870
rect 139830 666630 139920 666870
rect 140160 666630 140270 666870
rect 140510 666630 140600 666870
rect 140840 666630 140930 666870
rect 141170 666630 141260 666870
rect 141500 666630 141610 666870
rect 141850 666630 141940 666870
rect 142180 666630 142270 666870
rect 142510 666630 142600 666870
rect 142840 666630 142950 666870
rect 143190 666630 143280 666870
rect 143520 666630 143610 666870
rect 143850 666630 143940 666870
rect 144180 666630 144290 666870
rect 144530 666630 144550 666870
rect 133550 666540 144550 666630
rect 133550 666300 133570 666540
rect 133810 666300 133900 666540
rect 134140 666300 134230 666540
rect 134470 666300 134560 666540
rect 134800 666300 134910 666540
rect 135150 666300 135240 666540
rect 135480 666300 135570 666540
rect 135810 666300 135900 666540
rect 136140 666300 136250 666540
rect 136490 666300 136580 666540
rect 136820 666300 136910 666540
rect 137150 666300 137240 666540
rect 137480 666300 137590 666540
rect 137830 666300 137920 666540
rect 138160 666300 138250 666540
rect 138490 666300 138580 666540
rect 138820 666300 138930 666540
rect 139170 666300 139260 666540
rect 139500 666300 139590 666540
rect 139830 666300 139920 666540
rect 140160 666300 140270 666540
rect 140510 666300 140600 666540
rect 140840 666300 140930 666540
rect 141170 666300 141260 666540
rect 141500 666300 141610 666540
rect 141850 666300 141940 666540
rect 142180 666300 142270 666540
rect 142510 666300 142600 666540
rect 142840 666300 142950 666540
rect 143190 666300 143280 666540
rect 143520 666300 143610 666540
rect 143850 666300 143940 666540
rect 144180 666300 144290 666540
rect 144530 666300 144550 666540
rect 133550 666190 144550 666300
rect 133550 665950 133570 666190
rect 133810 665950 133900 666190
rect 134140 665950 134230 666190
rect 134470 665950 134560 666190
rect 134800 665950 134910 666190
rect 135150 665950 135240 666190
rect 135480 665950 135570 666190
rect 135810 665950 135900 666190
rect 136140 665950 136250 666190
rect 136490 665950 136580 666190
rect 136820 665950 136910 666190
rect 137150 665950 137240 666190
rect 137480 665950 137590 666190
rect 137830 665950 137920 666190
rect 138160 665950 138250 666190
rect 138490 665950 138580 666190
rect 138820 665950 138930 666190
rect 139170 665950 139260 666190
rect 139500 665950 139590 666190
rect 139830 665950 139920 666190
rect 140160 665950 140270 666190
rect 140510 665950 140600 666190
rect 140840 665950 140930 666190
rect 141170 665950 141260 666190
rect 141500 665950 141610 666190
rect 141850 665950 141940 666190
rect 142180 665950 142270 666190
rect 142510 665950 142600 666190
rect 142840 665950 142950 666190
rect 143190 665950 143280 666190
rect 143520 665950 143610 666190
rect 143850 665950 143940 666190
rect 144180 665950 144290 666190
rect 144530 665950 144550 666190
rect 133550 665860 144550 665950
rect 133550 665620 133570 665860
rect 133810 665620 133900 665860
rect 134140 665620 134230 665860
rect 134470 665620 134560 665860
rect 134800 665620 134910 665860
rect 135150 665620 135240 665860
rect 135480 665620 135570 665860
rect 135810 665620 135900 665860
rect 136140 665620 136250 665860
rect 136490 665620 136580 665860
rect 136820 665620 136910 665860
rect 137150 665620 137240 665860
rect 137480 665620 137590 665860
rect 137830 665620 137920 665860
rect 138160 665620 138250 665860
rect 138490 665620 138580 665860
rect 138820 665620 138930 665860
rect 139170 665620 139260 665860
rect 139500 665620 139590 665860
rect 139830 665620 139920 665860
rect 140160 665620 140270 665860
rect 140510 665620 140600 665860
rect 140840 665620 140930 665860
rect 141170 665620 141260 665860
rect 141500 665620 141610 665860
rect 141850 665620 141940 665860
rect 142180 665620 142270 665860
rect 142510 665620 142600 665860
rect 142840 665620 142950 665860
rect 143190 665620 143280 665860
rect 143520 665620 143610 665860
rect 143850 665620 143940 665860
rect 144180 665620 144290 665860
rect 144530 665620 144550 665860
rect 133550 665530 144550 665620
rect 133550 665290 133570 665530
rect 133810 665290 133900 665530
rect 134140 665290 134230 665530
rect 134470 665290 134560 665530
rect 134800 665290 134910 665530
rect 135150 665290 135240 665530
rect 135480 665290 135570 665530
rect 135810 665290 135900 665530
rect 136140 665290 136250 665530
rect 136490 665290 136580 665530
rect 136820 665290 136910 665530
rect 137150 665290 137240 665530
rect 137480 665290 137590 665530
rect 137830 665290 137920 665530
rect 138160 665290 138250 665530
rect 138490 665290 138580 665530
rect 138820 665290 138930 665530
rect 139170 665290 139260 665530
rect 139500 665290 139590 665530
rect 139830 665290 139920 665530
rect 140160 665290 140270 665530
rect 140510 665290 140600 665530
rect 140840 665290 140930 665530
rect 141170 665290 141260 665530
rect 141500 665290 141610 665530
rect 141850 665290 141940 665530
rect 142180 665290 142270 665530
rect 142510 665290 142600 665530
rect 142840 665290 142950 665530
rect 143190 665290 143280 665530
rect 143520 665290 143610 665530
rect 143850 665290 143940 665530
rect 144180 665290 144290 665530
rect 144530 665290 144550 665530
rect 133550 665200 144550 665290
rect 133550 664960 133570 665200
rect 133810 664960 133900 665200
rect 134140 664960 134230 665200
rect 134470 664960 134560 665200
rect 134800 664960 134910 665200
rect 135150 664960 135240 665200
rect 135480 664960 135570 665200
rect 135810 664960 135900 665200
rect 136140 664960 136250 665200
rect 136490 664960 136580 665200
rect 136820 664960 136910 665200
rect 137150 664960 137240 665200
rect 137480 664960 137590 665200
rect 137830 664960 137920 665200
rect 138160 664960 138250 665200
rect 138490 664960 138580 665200
rect 138820 664960 138930 665200
rect 139170 664960 139260 665200
rect 139500 664960 139590 665200
rect 139830 664960 139920 665200
rect 140160 664960 140270 665200
rect 140510 664960 140600 665200
rect 140840 664960 140930 665200
rect 141170 664960 141260 665200
rect 141500 664960 141610 665200
rect 141850 664960 141940 665200
rect 142180 664960 142270 665200
rect 142510 664960 142600 665200
rect 142840 664960 142950 665200
rect 143190 664960 143280 665200
rect 143520 664960 143610 665200
rect 143850 664960 143940 665200
rect 144180 664960 144290 665200
rect 144530 664960 144550 665200
rect 133550 664850 144550 664960
rect 133550 664610 133570 664850
rect 133810 664610 133900 664850
rect 134140 664610 134230 664850
rect 134470 664610 134560 664850
rect 134800 664610 134910 664850
rect 135150 664610 135240 664850
rect 135480 664610 135570 664850
rect 135810 664610 135900 664850
rect 136140 664610 136250 664850
rect 136490 664610 136580 664850
rect 136820 664610 136910 664850
rect 137150 664610 137240 664850
rect 137480 664610 137590 664850
rect 137830 664610 137920 664850
rect 138160 664610 138250 664850
rect 138490 664610 138580 664850
rect 138820 664610 138930 664850
rect 139170 664610 139260 664850
rect 139500 664610 139590 664850
rect 139830 664610 139920 664850
rect 140160 664610 140270 664850
rect 140510 664610 140600 664850
rect 140840 664610 140930 664850
rect 141170 664610 141260 664850
rect 141500 664610 141610 664850
rect 141850 664610 141940 664850
rect 142180 664610 142270 664850
rect 142510 664610 142600 664850
rect 142840 664610 142950 664850
rect 143190 664610 143280 664850
rect 143520 664610 143610 664850
rect 143850 664610 143940 664850
rect 144180 664610 144290 664850
rect 144530 664610 144550 664850
rect 133550 664520 144550 664610
rect 133550 664280 133570 664520
rect 133810 664280 133900 664520
rect 134140 664280 134230 664520
rect 134470 664280 134560 664520
rect 134800 664280 134910 664520
rect 135150 664280 135240 664520
rect 135480 664280 135570 664520
rect 135810 664280 135900 664520
rect 136140 664280 136250 664520
rect 136490 664280 136580 664520
rect 136820 664280 136910 664520
rect 137150 664280 137240 664520
rect 137480 664280 137590 664520
rect 137830 664280 137920 664520
rect 138160 664280 138250 664520
rect 138490 664280 138580 664520
rect 138820 664280 138930 664520
rect 139170 664280 139260 664520
rect 139500 664280 139590 664520
rect 139830 664280 139920 664520
rect 140160 664280 140270 664520
rect 140510 664280 140600 664520
rect 140840 664280 140930 664520
rect 141170 664280 141260 664520
rect 141500 664280 141610 664520
rect 141850 664280 141940 664520
rect 142180 664280 142270 664520
rect 142510 664280 142600 664520
rect 142840 664280 142950 664520
rect 143190 664280 143280 664520
rect 143520 664280 143610 664520
rect 143850 664280 143940 664520
rect 144180 664280 144290 664520
rect 144530 664280 144550 664520
rect 133550 664190 144550 664280
rect 133550 663950 133570 664190
rect 133810 663950 133900 664190
rect 134140 663950 134230 664190
rect 134470 663950 134560 664190
rect 134800 663950 134910 664190
rect 135150 663950 135240 664190
rect 135480 663950 135570 664190
rect 135810 663950 135900 664190
rect 136140 663950 136250 664190
rect 136490 663950 136580 664190
rect 136820 663950 136910 664190
rect 137150 663950 137240 664190
rect 137480 663950 137590 664190
rect 137830 663950 137920 664190
rect 138160 663950 138250 664190
rect 138490 663950 138580 664190
rect 138820 663950 138930 664190
rect 139170 663950 139260 664190
rect 139500 663950 139590 664190
rect 139830 663950 139920 664190
rect 140160 663950 140270 664190
rect 140510 663950 140600 664190
rect 140840 663950 140930 664190
rect 141170 663950 141260 664190
rect 141500 663950 141610 664190
rect 141850 663950 141940 664190
rect 142180 663950 142270 664190
rect 142510 663950 142600 664190
rect 142840 663950 142950 664190
rect 143190 663950 143280 664190
rect 143520 663950 143610 664190
rect 143850 663950 143940 664190
rect 144180 663950 144290 664190
rect 144530 663950 144550 664190
rect 133550 663860 144550 663950
rect 133550 663620 133570 663860
rect 133810 663620 133900 663860
rect 134140 663620 134230 663860
rect 134470 663620 134560 663860
rect 134800 663620 134910 663860
rect 135150 663620 135240 663860
rect 135480 663620 135570 663860
rect 135810 663620 135900 663860
rect 136140 663620 136250 663860
rect 136490 663620 136580 663860
rect 136820 663620 136910 663860
rect 137150 663620 137240 663860
rect 137480 663620 137590 663860
rect 137830 663620 137920 663860
rect 138160 663620 138250 663860
rect 138490 663620 138580 663860
rect 138820 663620 138930 663860
rect 139170 663620 139260 663860
rect 139500 663620 139590 663860
rect 139830 663620 139920 663860
rect 140160 663620 140270 663860
rect 140510 663620 140600 663860
rect 140840 663620 140930 663860
rect 141170 663620 141260 663860
rect 141500 663620 141610 663860
rect 141850 663620 141940 663860
rect 142180 663620 142270 663860
rect 142510 663620 142600 663860
rect 142840 663620 142950 663860
rect 143190 663620 143280 663860
rect 143520 663620 143610 663860
rect 143850 663620 143940 663860
rect 144180 663620 144290 663860
rect 144530 663620 144550 663860
rect 133550 663510 144550 663620
rect 133550 663270 133570 663510
rect 133810 663270 133900 663510
rect 134140 663270 134230 663510
rect 134470 663270 134560 663510
rect 134800 663270 134910 663510
rect 135150 663270 135240 663510
rect 135480 663270 135570 663510
rect 135810 663270 135900 663510
rect 136140 663270 136250 663510
rect 136490 663270 136580 663510
rect 136820 663270 136910 663510
rect 137150 663270 137240 663510
rect 137480 663270 137590 663510
rect 137830 663270 137920 663510
rect 138160 663270 138250 663510
rect 138490 663270 138580 663510
rect 138820 663270 138930 663510
rect 139170 663270 139260 663510
rect 139500 663270 139590 663510
rect 139830 663270 139920 663510
rect 140160 663270 140270 663510
rect 140510 663270 140600 663510
rect 140840 663270 140930 663510
rect 141170 663270 141260 663510
rect 141500 663270 141610 663510
rect 141850 663270 141940 663510
rect 142180 663270 142270 663510
rect 142510 663270 142600 663510
rect 142840 663270 142950 663510
rect 143190 663270 143280 663510
rect 143520 663270 143610 663510
rect 143850 663270 143940 663510
rect 144180 663270 144290 663510
rect 144530 663270 144550 663510
rect 133550 663180 144550 663270
rect 133550 662940 133570 663180
rect 133810 662940 133900 663180
rect 134140 662940 134230 663180
rect 134470 662940 134560 663180
rect 134800 662940 134910 663180
rect 135150 662940 135240 663180
rect 135480 662940 135570 663180
rect 135810 662940 135900 663180
rect 136140 662940 136250 663180
rect 136490 662940 136580 663180
rect 136820 662940 136910 663180
rect 137150 662940 137240 663180
rect 137480 662940 137590 663180
rect 137830 662940 137920 663180
rect 138160 662940 138250 663180
rect 138490 662940 138580 663180
rect 138820 662940 138930 663180
rect 139170 662940 139260 663180
rect 139500 662940 139590 663180
rect 139830 662940 139920 663180
rect 140160 662940 140270 663180
rect 140510 662940 140600 663180
rect 140840 662940 140930 663180
rect 141170 662940 141260 663180
rect 141500 662940 141610 663180
rect 141850 662940 141940 663180
rect 142180 662940 142270 663180
rect 142510 662940 142600 663180
rect 142840 662940 142950 663180
rect 143190 662940 143280 663180
rect 143520 662940 143610 663180
rect 143850 662940 143940 663180
rect 144180 662940 144290 663180
rect 144530 662940 144550 663180
rect 133550 662850 144550 662940
rect 133550 662610 133570 662850
rect 133810 662610 133900 662850
rect 134140 662610 134230 662850
rect 134470 662610 134560 662850
rect 134800 662610 134910 662850
rect 135150 662610 135240 662850
rect 135480 662610 135570 662850
rect 135810 662610 135900 662850
rect 136140 662610 136250 662850
rect 136490 662610 136580 662850
rect 136820 662610 136910 662850
rect 137150 662610 137240 662850
rect 137480 662610 137590 662850
rect 137830 662610 137920 662850
rect 138160 662610 138250 662850
rect 138490 662610 138580 662850
rect 138820 662610 138930 662850
rect 139170 662610 139260 662850
rect 139500 662610 139590 662850
rect 139830 662610 139920 662850
rect 140160 662610 140270 662850
rect 140510 662610 140600 662850
rect 140840 662610 140930 662850
rect 141170 662610 141260 662850
rect 141500 662610 141610 662850
rect 141850 662610 141940 662850
rect 142180 662610 142270 662850
rect 142510 662610 142600 662850
rect 142840 662610 142950 662850
rect 143190 662610 143280 662850
rect 143520 662610 143610 662850
rect 143850 662610 143940 662850
rect 144180 662610 144290 662850
rect 144530 662610 144550 662850
rect 133550 662520 144550 662610
rect 133550 662280 133570 662520
rect 133810 662280 133900 662520
rect 134140 662280 134230 662520
rect 134470 662280 134560 662520
rect 134800 662280 134910 662520
rect 135150 662280 135240 662520
rect 135480 662280 135570 662520
rect 135810 662280 135900 662520
rect 136140 662280 136250 662520
rect 136490 662280 136580 662520
rect 136820 662280 136910 662520
rect 137150 662280 137240 662520
rect 137480 662280 137590 662520
rect 137830 662280 137920 662520
rect 138160 662280 138250 662520
rect 138490 662280 138580 662520
rect 138820 662280 138930 662520
rect 139170 662280 139260 662520
rect 139500 662280 139590 662520
rect 139830 662280 139920 662520
rect 140160 662280 140270 662520
rect 140510 662280 140600 662520
rect 140840 662280 140930 662520
rect 141170 662280 141260 662520
rect 141500 662280 141610 662520
rect 141850 662280 141940 662520
rect 142180 662280 142270 662520
rect 142510 662280 142600 662520
rect 142840 662280 142950 662520
rect 143190 662280 143280 662520
rect 143520 662280 143610 662520
rect 143850 662280 143940 662520
rect 144180 662280 144290 662520
rect 144530 662280 144550 662520
rect 133550 662170 144550 662280
rect 133550 661930 133570 662170
rect 133810 661930 133900 662170
rect 134140 661930 134230 662170
rect 134470 661930 134560 662170
rect 134800 661930 134910 662170
rect 135150 661930 135240 662170
rect 135480 661930 135570 662170
rect 135810 661930 135900 662170
rect 136140 661930 136250 662170
rect 136490 661930 136580 662170
rect 136820 661930 136910 662170
rect 137150 661930 137240 662170
rect 137480 661930 137590 662170
rect 137830 661930 137920 662170
rect 138160 661930 138250 662170
rect 138490 661930 138580 662170
rect 138820 661930 138930 662170
rect 139170 661930 139260 662170
rect 139500 661930 139590 662170
rect 139830 661930 139920 662170
rect 140160 661930 140270 662170
rect 140510 661930 140600 662170
rect 140840 661930 140930 662170
rect 141170 661930 141260 662170
rect 141500 661930 141610 662170
rect 141850 661930 141940 662170
rect 142180 661930 142270 662170
rect 142510 661930 142600 662170
rect 142840 661930 142950 662170
rect 143190 661930 143280 662170
rect 143520 661930 143610 662170
rect 143850 661930 143940 662170
rect 144180 661930 144290 662170
rect 144530 661930 144550 662170
rect 133550 661840 144550 661930
rect 133550 661600 133570 661840
rect 133810 661600 133900 661840
rect 134140 661600 134230 661840
rect 134470 661600 134560 661840
rect 134800 661600 134910 661840
rect 135150 661600 135240 661840
rect 135480 661600 135570 661840
rect 135810 661600 135900 661840
rect 136140 661600 136250 661840
rect 136490 661600 136580 661840
rect 136820 661600 136910 661840
rect 137150 661600 137240 661840
rect 137480 661600 137590 661840
rect 137830 661600 137920 661840
rect 138160 661600 138250 661840
rect 138490 661600 138580 661840
rect 138820 661600 138930 661840
rect 139170 661600 139260 661840
rect 139500 661600 139590 661840
rect 139830 661600 139920 661840
rect 140160 661600 140270 661840
rect 140510 661600 140600 661840
rect 140840 661600 140930 661840
rect 141170 661600 141260 661840
rect 141500 661600 141610 661840
rect 141850 661600 141940 661840
rect 142180 661600 142270 661840
rect 142510 661600 142600 661840
rect 142840 661600 142950 661840
rect 143190 661600 143280 661840
rect 143520 661600 143610 661840
rect 143850 661600 143940 661840
rect 144180 661600 144290 661840
rect 144530 661600 144550 661840
rect 133550 661510 144550 661600
rect 133550 661270 133570 661510
rect 133810 661270 133900 661510
rect 134140 661270 134230 661510
rect 134470 661270 134560 661510
rect 134800 661270 134910 661510
rect 135150 661270 135240 661510
rect 135480 661270 135570 661510
rect 135810 661270 135900 661510
rect 136140 661270 136250 661510
rect 136490 661270 136580 661510
rect 136820 661270 136910 661510
rect 137150 661270 137240 661510
rect 137480 661270 137590 661510
rect 137830 661270 137920 661510
rect 138160 661270 138250 661510
rect 138490 661270 138580 661510
rect 138820 661270 138930 661510
rect 139170 661270 139260 661510
rect 139500 661270 139590 661510
rect 139830 661270 139920 661510
rect 140160 661270 140270 661510
rect 140510 661270 140600 661510
rect 140840 661270 140930 661510
rect 141170 661270 141260 661510
rect 141500 661270 141610 661510
rect 141850 661270 141940 661510
rect 142180 661270 142270 661510
rect 142510 661270 142600 661510
rect 142840 661270 142950 661510
rect 143190 661270 143280 661510
rect 143520 661270 143610 661510
rect 143850 661270 143940 661510
rect 144180 661270 144290 661510
rect 144530 661270 144550 661510
rect 133550 661180 144550 661270
rect 133550 660940 133570 661180
rect 133810 660940 133900 661180
rect 134140 660940 134230 661180
rect 134470 660940 134560 661180
rect 134800 660940 134910 661180
rect 135150 660940 135240 661180
rect 135480 660940 135570 661180
rect 135810 660940 135900 661180
rect 136140 660940 136250 661180
rect 136490 660940 136580 661180
rect 136820 660940 136910 661180
rect 137150 660940 137240 661180
rect 137480 660940 137590 661180
rect 137830 660940 137920 661180
rect 138160 660940 138250 661180
rect 138490 660940 138580 661180
rect 138820 660940 138930 661180
rect 139170 660940 139260 661180
rect 139500 660940 139590 661180
rect 139830 660940 139920 661180
rect 140160 660940 140270 661180
rect 140510 660940 140600 661180
rect 140840 660940 140930 661180
rect 141170 660940 141260 661180
rect 141500 660940 141610 661180
rect 141850 660940 141940 661180
rect 142180 660940 142270 661180
rect 142510 660940 142600 661180
rect 142840 660940 142950 661180
rect 143190 660940 143280 661180
rect 143520 660940 143610 661180
rect 143850 660940 143940 661180
rect 144180 660940 144290 661180
rect 144530 660940 144550 661180
rect 133550 660920 144550 660940
rect 144930 671900 155930 671920
rect 144930 671660 144950 671900
rect 145190 671660 145280 671900
rect 145520 671660 145610 671900
rect 145850 671660 145940 671900
rect 146180 671660 146290 671900
rect 146530 671660 146620 671900
rect 146860 671660 146950 671900
rect 147190 671660 147280 671900
rect 147520 671660 147630 671900
rect 147870 671660 147960 671900
rect 148200 671660 148290 671900
rect 148530 671660 148620 671900
rect 148860 671660 148970 671900
rect 149210 671660 149300 671900
rect 149540 671660 149630 671900
rect 149870 671660 149960 671900
rect 150200 671660 150310 671900
rect 150550 671660 150640 671900
rect 150880 671660 150970 671900
rect 151210 671660 151300 671900
rect 151540 671660 151650 671900
rect 151890 671660 151980 671900
rect 152220 671660 152310 671900
rect 152550 671660 152640 671900
rect 152880 671660 152990 671900
rect 153230 671660 153320 671900
rect 153560 671660 153650 671900
rect 153890 671660 153980 671900
rect 154220 671660 154330 671900
rect 154570 671660 154660 671900
rect 154900 671660 154990 671900
rect 155230 671660 155320 671900
rect 155560 671660 155670 671900
rect 155910 671660 155930 671900
rect 144930 671550 155930 671660
rect 144930 671310 144950 671550
rect 145190 671310 145280 671550
rect 145520 671310 145610 671550
rect 145850 671310 145940 671550
rect 146180 671310 146290 671550
rect 146530 671310 146620 671550
rect 146860 671310 146950 671550
rect 147190 671310 147280 671550
rect 147520 671310 147630 671550
rect 147870 671310 147960 671550
rect 148200 671310 148290 671550
rect 148530 671310 148620 671550
rect 148860 671310 148970 671550
rect 149210 671310 149300 671550
rect 149540 671310 149630 671550
rect 149870 671310 149960 671550
rect 150200 671310 150310 671550
rect 150550 671310 150640 671550
rect 150880 671310 150970 671550
rect 151210 671310 151300 671550
rect 151540 671310 151650 671550
rect 151890 671310 151980 671550
rect 152220 671310 152310 671550
rect 152550 671310 152640 671550
rect 152880 671310 152990 671550
rect 153230 671310 153320 671550
rect 153560 671310 153650 671550
rect 153890 671310 153980 671550
rect 154220 671310 154330 671550
rect 154570 671310 154660 671550
rect 154900 671310 154990 671550
rect 155230 671310 155320 671550
rect 155560 671310 155670 671550
rect 155910 671310 155930 671550
rect 144930 671220 155930 671310
rect 144930 670980 144950 671220
rect 145190 670980 145280 671220
rect 145520 670980 145610 671220
rect 145850 670980 145940 671220
rect 146180 670980 146290 671220
rect 146530 670980 146620 671220
rect 146860 670980 146950 671220
rect 147190 670980 147280 671220
rect 147520 670980 147630 671220
rect 147870 670980 147960 671220
rect 148200 670980 148290 671220
rect 148530 670980 148620 671220
rect 148860 670980 148970 671220
rect 149210 670980 149300 671220
rect 149540 670980 149630 671220
rect 149870 670980 149960 671220
rect 150200 670980 150310 671220
rect 150550 670980 150640 671220
rect 150880 670980 150970 671220
rect 151210 670980 151300 671220
rect 151540 670980 151650 671220
rect 151890 670980 151980 671220
rect 152220 670980 152310 671220
rect 152550 670980 152640 671220
rect 152880 670980 152990 671220
rect 153230 670980 153320 671220
rect 153560 670980 153650 671220
rect 153890 670980 153980 671220
rect 154220 670980 154330 671220
rect 154570 670980 154660 671220
rect 154900 670980 154990 671220
rect 155230 670980 155320 671220
rect 155560 670980 155670 671220
rect 155910 670980 155930 671220
rect 144930 670890 155930 670980
rect 144930 670650 144950 670890
rect 145190 670650 145280 670890
rect 145520 670650 145610 670890
rect 145850 670650 145940 670890
rect 146180 670650 146290 670890
rect 146530 670650 146620 670890
rect 146860 670650 146950 670890
rect 147190 670650 147280 670890
rect 147520 670650 147630 670890
rect 147870 670650 147960 670890
rect 148200 670650 148290 670890
rect 148530 670650 148620 670890
rect 148860 670650 148970 670890
rect 149210 670650 149300 670890
rect 149540 670650 149630 670890
rect 149870 670650 149960 670890
rect 150200 670650 150310 670890
rect 150550 670650 150640 670890
rect 150880 670650 150970 670890
rect 151210 670650 151300 670890
rect 151540 670650 151650 670890
rect 151890 670650 151980 670890
rect 152220 670650 152310 670890
rect 152550 670650 152640 670890
rect 152880 670650 152990 670890
rect 153230 670650 153320 670890
rect 153560 670650 153650 670890
rect 153890 670650 153980 670890
rect 154220 670650 154330 670890
rect 154570 670650 154660 670890
rect 154900 670650 154990 670890
rect 155230 670650 155320 670890
rect 155560 670650 155670 670890
rect 155910 670650 155930 670890
rect 144930 670560 155930 670650
rect 144930 670320 144950 670560
rect 145190 670320 145280 670560
rect 145520 670320 145610 670560
rect 145850 670320 145940 670560
rect 146180 670320 146290 670560
rect 146530 670320 146620 670560
rect 146860 670320 146950 670560
rect 147190 670320 147280 670560
rect 147520 670320 147630 670560
rect 147870 670320 147960 670560
rect 148200 670320 148290 670560
rect 148530 670320 148620 670560
rect 148860 670320 148970 670560
rect 149210 670320 149300 670560
rect 149540 670320 149630 670560
rect 149870 670320 149960 670560
rect 150200 670320 150310 670560
rect 150550 670320 150640 670560
rect 150880 670320 150970 670560
rect 151210 670320 151300 670560
rect 151540 670320 151650 670560
rect 151890 670320 151980 670560
rect 152220 670320 152310 670560
rect 152550 670320 152640 670560
rect 152880 670320 152990 670560
rect 153230 670320 153320 670560
rect 153560 670320 153650 670560
rect 153890 670320 153980 670560
rect 154220 670320 154330 670560
rect 154570 670320 154660 670560
rect 154900 670320 154990 670560
rect 155230 670320 155320 670560
rect 155560 670320 155670 670560
rect 155910 670320 155930 670560
rect 144930 670210 155930 670320
rect 144930 669970 144950 670210
rect 145190 669970 145280 670210
rect 145520 669970 145610 670210
rect 145850 669970 145940 670210
rect 146180 669970 146290 670210
rect 146530 669970 146620 670210
rect 146860 669970 146950 670210
rect 147190 669970 147280 670210
rect 147520 669970 147630 670210
rect 147870 669970 147960 670210
rect 148200 669970 148290 670210
rect 148530 669970 148620 670210
rect 148860 669970 148970 670210
rect 149210 669970 149300 670210
rect 149540 669970 149630 670210
rect 149870 669970 149960 670210
rect 150200 669970 150310 670210
rect 150550 669970 150640 670210
rect 150880 669970 150970 670210
rect 151210 669970 151300 670210
rect 151540 669970 151650 670210
rect 151890 669970 151980 670210
rect 152220 669970 152310 670210
rect 152550 669970 152640 670210
rect 152880 669970 152990 670210
rect 153230 669970 153320 670210
rect 153560 669970 153650 670210
rect 153890 669970 153980 670210
rect 154220 669970 154330 670210
rect 154570 669970 154660 670210
rect 154900 669970 154990 670210
rect 155230 669970 155320 670210
rect 155560 669970 155670 670210
rect 155910 669970 155930 670210
rect 144930 669880 155930 669970
rect 144930 669640 144950 669880
rect 145190 669640 145280 669880
rect 145520 669640 145610 669880
rect 145850 669640 145940 669880
rect 146180 669640 146290 669880
rect 146530 669640 146620 669880
rect 146860 669640 146950 669880
rect 147190 669640 147280 669880
rect 147520 669640 147630 669880
rect 147870 669640 147960 669880
rect 148200 669640 148290 669880
rect 148530 669640 148620 669880
rect 148860 669640 148970 669880
rect 149210 669640 149300 669880
rect 149540 669640 149630 669880
rect 149870 669640 149960 669880
rect 150200 669640 150310 669880
rect 150550 669640 150640 669880
rect 150880 669640 150970 669880
rect 151210 669640 151300 669880
rect 151540 669640 151650 669880
rect 151890 669640 151980 669880
rect 152220 669640 152310 669880
rect 152550 669640 152640 669880
rect 152880 669640 152990 669880
rect 153230 669640 153320 669880
rect 153560 669640 153650 669880
rect 153890 669640 153980 669880
rect 154220 669640 154330 669880
rect 154570 669640 154660 669880
rect 154900 669640 154990 669880
rect 155230 669640 155320 669880
rect 155560 669640 155670 669880
rect 155910 669640 155930 669880
rect 144930 669550 155930 669640
rect 144930 669310 144950 669550
rect 145190 669310 145280 669550
rect 145520 669310 145610 669550
rect 145850 669310 145940 669550
rect 146180 669310 146290 669550
rect 146530 669310 146620 669550
rect 146860 669310 146950 669550
rect 147190 669310 147280 669550
rect 147520 669310 147630 669550
rect 147870 669310 147960 669550
rect 148200 669310 148290 669550
rect 148530 669310 148620 669550
rect 148860 669310 148970 669550
rect 149210 669310 149300 669550
rect 149540 669310 149630 669550
rect 149870 669310 149960 669550
rect 150200 669310 150310 669550
rect 150550 669310 150640 669550
rect 150880 669310 150970 669550
rect 151210 669310 151300 669550
rect 151540 669310 151650 669550
rect 151890 669310 151980 669550
rect 152220 669310 152310 669550
rect 152550 669310 152640 669550
rect 152880 669310 152990 669550
rect 153230 669310 153320 669550
rect 153560 669310 153650 669550
rect 153890 669310 153980 669550
rect 154220 669310 154330 669550
rect 154570 669310 154660 669550
rect 154900 669310 154990 669550
rect 155230 669310 155320 669550
rect 155560 669310 155670 669550
rect 155910 669310 155930 669550
rect 144930 669220 155930 669310
rect 144930 668980 144950 669220
rect 145190 668980 145280 669220
rect 145520 668980 145610 669220
rect 145850 668980 145940 669220
rect 146180 668980 146290 669220
rect 146530 668980 146620 669220
rect 146860 668980 146950 669220
rect 147190 668980 147280 669220
rect 147520 668980 147630 669220
rect 147870 668980 147960 669220
rect 148200 668980 148290 669220
rect 148530 668980 148620 669220
rect 148860 668980 148970 669220
rect 149210 668980 149300 669220
rect 149540 668980 149630 669220
rect 149870 668980 149960 669220
rect 150200 668980 150310 669220
rect 150550 668980 150640 669220
rect 150880 668980 150970 669220
rect 151210 668980 151300 669220
rect 151540 668980 151650 669220
rect 151890 668980 151980 669220
rect 152220 668980 152310 669220
rect 152550 668980 152640 669220
rect 152880 668980 152990 669220
rect 153230 668980 153320 669220
rect 153560 668980 153650 669220
rect 153890 668980 153980 669220
rect 154220 668980 154330 669220
rect 154570 668980 154660 669220
rect 154900 668980 154990 669220
rect 155230 668980 155320 669220
rect 155560 668980 155670 669220
rect 155910 668980 155930 669220
rect 144930 668870 155930 668980
rect 144930 668630 144950 668870
rect 145190 668630 145280 668870
rect 145520 668630 145610 668870
rect 145850 668630 145940 668870
rect 146180 668630 146290 668870
rect 146530 668630 146620 668870
rect 146860 668630 146950 668870
rect 147190 668630 147280 668870
rect 147520 668630 147630 668870
rect 147870 668630 147960 668870
rect 148200 668630 148290 668870
rect 148530 668630 148620 668870
rect 148860 668630 148970 668870
rect 149210 668630 149300 668870
rect 149540 668630 149630 668870
rect 149870 668630 149960 668870
rect 150200 668630 150310 668870
rect 150550 668630 150640 668870
rect 150880 668630 150970 668870
rect 151210 668630 151300 668870
rect 151540 668630 151650 668870
rect 151890 668630 151980 668870
rect 152220 668630 152310 668870
rect 152550 668630 152640 668870
rect 152880 668630 152990 668870
rect 153230 668630 153320 668870
rect 153560 668630 153650 668870
rect 153890 668630 153980 668870
rect 154220 668630 154330 668870
rect 154570 668630 154660 668870
rect 154900 668630 154990 668870
rect 155230 668630 155320 668870
rect 155560 668630 155670 668870
rect 155910 668630 155930 668870
rect 144930 668540 155930 668630
rect 144930 668300 144950 668540
rect 145190 668300 145280 668540
rect 145520 668300 145610 668540
rect 145850 668300 145940 668540
rect 146180 668300 146290 668540
rect 146530 668300 146620 668540
rect 146860 668300 146950 668540
rect 147190 668300 147280 668540
rect 147520 668300 147630 668540
rect 147870 668300 147960 668540
rect 148200 668300 148290 668540
rect 148530 668300 148620 668540
rect 148860 668300 148970 668540
rect 149210 668300 149300 668540
rect 149540 668300 149630 668540
rect 149870 668300 149960 668540
rect 150200 668300 150310 668540
rect 150550 668300 150640 668540
rect 150880 668300 150970 668540
rect 151210 668300 151300 668540
rect 151540 668300 151650 668540
rect 151890 668300 151980 668540
rect 152220 668300 152310 668540
rect 152550 668300 152640 668540
rect 152880 668300 152990 668540
rect 153230 668300 153320 668540
rect 153560 668300 153650 668540
rect 153890 668300 153980 668540
rect 154220 668300 154330 668540
rect 154570 668300 154660 668540
rect 154900 668300 154990 668540
rect 155230 668300 155320 668540
rect 155560 668300 155670 668540
rect 155910 668300 155930 668540
rect 144930 668210 155930 668300
rect 144930 667970 144950 668210
rect 145190 667970 145280 668210
rect 145520 667970 145610 668210
rect 145850 667970 145940 668210
rect 146180 667970 146290 668210
rect 146530 667970 146620 668210
rect 146860 667970 146950 668210
rect 147190 667970 147280 668210
rect 147520 667970 147630 668210
rect 147870 667970 147960 668210
rect 148200 667970 148290 668210
rect 148530 667970 148620 668210
rect 148860 667970 148970 668210
rect 149210 667970 149300 668210
rect 149540 667970 149630 668210
rect 149870 667970 149960 668210
rect 150200 667970 150310 668210
rect 150550 667970 150640 668210
rect 150880 667970 150970 668210
rect 151210 667970 151300 668210
rect 151540 667970 151650 668210
rect 151890 667970 151980 668210
rect 152220 667970 152310 668210
rect 152550 667970 152640 668210
rect 152880 667970 152990 668210
rect 153230 667970 153320 668210
rect 153560 667970 153650 668210
rect 153890 667970 153980 668210
rect 154220 667970 154330 668210
rect 154570 667970 154660 668210
rect 154900 667970 154990 668210
rect 155230 667970 155320 668210
rect 155560 667970 155670 668210
rect 155910 667970 155930 668210
rect 144930 667880 155930 667970
rect 144930 667640 144950 667880
rect 145190 667640 145280 667880
rect 145520 667640 145610 667880
rect 145850 667640 145940 667880
rect 146180 667640 146290 667880
rect 146530 667640 146620 667880
rect 146860 667640 146950 667880
rect 147190 667640 147280 667880
rect 147520 667640 147630 667880
rect 147870 667640 147960 667880
rect 148200 667640 148290 667880
rect 148530 667640 148620 667880
rect 148860 667640 148970 667880
rect 149210 667640 149300 667880
rect 149540 667640 149630 667880
rect 149870 667640 149960 667880
rect 150200 667640 150310 667880
rect 150550 667640 150640 667880
rect 150880 667640 150970 667880
rect 151210 667640 151300 667880
rect 151540 667640 151650 667880
rect 151890 667640 151980 667880
rect 152220 667640 152310 667880
rect 152550 667640 152640 667880
rect 152880 667640 152990 667880
rect 153230 667640 153320 667880
rect 153560 667640 153650 667880
rect 153890 667640 153980 667880
rect 154220 667640 154330 667880
rect 154570 667640 154660 667880
rect 154900 667640 154990 667880
rect 155230 667640 155320 667880
rect 155560 667640 155670 667880
rect 155910 667640 155930 667880
rect 144930 667530 155930 667640
rect 144930 667290 144950 667530
rect 145190 667290 145280 667530
rect 145520 667290 145610 667530
rect 145850 667290 145940 667530
rect 146180 667290 146290 667530
rect 146530 667290 146620 667530
rect 146860 667290 146950 667530
rect 147190 667290 147280 667530
rect 147520 667290 147630 667530
rect 147870 667290 147960 667530
rect 148200 667290 148290 667530
rect 148530 667290 148620 667530
rect 148860 667290 148970 667530
rect 149210 667290 149300 667530
rect 149540 667290 149630 667530
rect 149870 667290 149960 667530
rect 150200 667290 150310 667530
rect 150550 667290 150640 667530
rect 150880 667290 150970 667530
rect 151210 667290 151300 667530
rect 151540 667290 151650 667530
rect 151890 667290 151980 667530
rect 152220 667290 152310 667530
rect 152550 667290 152640 667530
rect 152880 667290 152990 667530
rect 153230 667290 153320 667530
rect 153560 667290 153650 667530
rect 153890 667290 153980 667530
rect 154220 667290 154330 667530
rect 154570 667290 154660 667530
rect 154900 667290 154990 667530
rect 155230 667290 155320 667530
rect 155560 667290 155670 667530
rect 155910 667290 155930 667530
rect 144930 667200 155930 667290
rect 144930 666960 144950 667200
rect 145190 666960 145280 667200
rect 145520 666960 145610 667200
rect 145850 666960 145940 667200
rect 146180 666960 146290 667200
rect 146530 666960 146620 667200
rect 146860 666960 146950 667200
rect 147190 666960 147280 667200
rect 147520 666960 147630 667200
rect 147870 666960 147960 667200
rect 148200 666960 148290 667200
rect 148530 666960 148620 667200
rect 148860 666960 148970 667200
rect 149210 666960 149300 667200
rect 149540 666960 149630 667200
rect 149870 666960 149960 667200
rect 150200 666960 150310 667200
rect 150550 666960 150640 667200
rect 150880 666960 150970 667200
rect 151210 666960 151300 667200
rect 151540 666960 151650 667200
rect 151890 666960 151980 667200
rect 152220 666960 152310 667200
rect 152550 666960 152640 667200
rect 152880 666960 152990 667200
rect 153230 666960 153320 667200
rect 153560 666960 153650 667200
rect 153890 666960 153980 667200
rect 154220 666960 154330 667200
rect 154570 666960 154660 667200
rect 154900 666960 154990 667200
rect 155230 666960 155320 667200
rect 155560 666960 155670 667200
rect 155910 666960 155930 667200
rect 144930 666870 155930 666960
rect 144930 666630 144950 666870
rect 145190 666630 145280 666870
rect 145520 666630 145610 666870
rect 145850 666630 145940 666870
rect 146180 666630 146290 666870
rect 146530 666630 146620 666870
rect 146860 666630 146950 666870
rect 147190 666630 147280 666870
rect 147520 666630 147630 666870
rect 147870 666630 147960 666870
rect 148200 666630 148290 666870
rect 148530 666630 148620 666870
rect 148860 666630 148970 666870
rect 149210 666630 149300 666870
rect 149540 666630 149630 666870
rect 149870 666630 149960 666870
rect 150200 666630 150310 666870
rect 150550 666630 150640 666870
rect 150880 666630 150970 666870
rect 151210 666630 151300 666870
rect 151540 666630 151650 666870
rect 151890 666630 151980 666870
rect 152220 666630 152310 666870
rect 152550 666630 152640 666870
rect 152880 666630 152990 666870
rect 153230 666630 153320 666870
rect 153560 666630 153650 666870
rect 153890 666630 153980 666870
rect 154220 666630 154330 666870
rect 154570 666630 154660 666870
rect 154900 666630 154990 666870
rect 155230 666630 155320 666870
rect 155560 666630 155670 666870
rect 155910 666630 155930 666870
rect 144930 666540 155930 666630
rect 144930 666300 144950 666540
rect 145190 666300 145280 666540
rect 145520 666300 145610 666540
rect 145850 666300 145940 666540
rect 146180 666300 146290 666540
rect 146530 666300 146620 666540
rect 146860 666300 146950 666540
rect 147190 666300 147280 666540
rect 147520 666300 147630 666540
rect 147870 666300 147960 666540
rect 148200 666300 148290 666540
rect 148530 666300 148620 666540
rect 148860 666300 148970 666540
rect 149210 666300 149300 666540
rect 149540 666300 149630 666540
rect 149870 666300 149960 666540
rect 150200 666300 150310 666540
rect 150550 666300 150640 666540
rect 150880 666300 150970 666540
rect 151210 666300 151300 666540
rect 151540 666300 151650 666540
rect 151890 666300 151980 666540
rect 152220 666300 152310 666540
rect 152550 666300 152640 666540
rect 152880 666300 152990 666540
rect 153230 666300 153320 666540
rect 153560 666300 153650 666540
rect 153890 666300 153980 666540
rect 154220 666300 154330 666540
rect 154570 666300 154660 666540
rect 154900 666300 154990 666540
rect 155230 666300 155320 666540
rect 155560 666300 155670 666540
rect 155910 666300 155930 666540
rect 144930 666190 155930 666300
rect 144930 665950 144950 666190
rect 145190 665950 145280 666190
rect 145520 665950 145610 666190
rect 145850 665950 145940 666190
rect 146180 665950 146290 666190
rect 146530 665950 146620 666190
rect 146860 665950 146950 666190
rect 147190 665950 147280 666190
rect 147520 665950 147630 666190
rect 147870 665950 147960 666190
rect 148200 665950 148290 666190
rect 148530 665950 148620 666190
rect 148860 665950 148970 666190
rect 149210 665950 149300 666190
rect 149540 665950 149630 666190
rect 149870 665950 149960 666190
rect 150200 665950 150310 666190
rect 150550 665950 150640 666190
rect 150880 665950 150970 666190
rect 151210 665950 151300 666190
rect 151540 665950 151650 666190
rect 151890 665950 151980 666190
rect 152220 665950 152310 666190
rect 152550 665950 152640 666190
rect 152880 665950 152990 666190
rect 153230 665950 153320 666190
rect 153560 665950 153650 666190
rect 153890 665950 153980 666190
rect 154220 665950 154330 666190
rect 154570 665950 154660 666190
rect 154900 665950 154990 666190
rect 155230 665950 155320 666190
rect 155560 665950 155670 666190
rect 155910 665950 155930 666190
rect 144930 665860 155930 665950
rect 144930 665620 144950 665860
rect 145190 665620 145280 665860
rect 145520 665620 145610 665860
rect 145850 665620 145940 665860
rect 146180 665620 146290 665860
rect 146530 665620 146620 665860
rect 146860 665620 146950 665860
rect 147190 665620 147280 665860
rect 147520 665620 147630 665860
rect 147870 665620 147960 665860
rect 148200 665620 148290 665860
rect 148530 665620 148620 665860
rect 148860 665620 148970 665860
rect 149210 665620 149300 665860
rect 149540 665620 149630 665860
rect 149870 665620 149960 665860
rect 150200 665620 150310 665860
rect 150550 665620 150640 665860
rect 150880 665620 150970 665860
rect 151210 665620 151300 665860
rect 151540 665620 151650 665860
rect 151890 665620 151980 665860
rect 152220 665620 152310 665860
rect 152550 665620 152640 665860
rect 152880 665620 152990 665860
rect 153230 665620 153320 665860
rect 153560 665620 153650 665860
rect 153890 665620 153980 665860
rect 154220 665620 154330 665860
rect 154570 665620 154660 665860
rect 154900 665620 154990 665860
rect 155230 665620 155320 665860
rect 155560 665620 155670 665860
rect 155910 665620 155930 665860
rect 144930 665530 155930 665620
rect 144930 665290 144950 665530
rect 145190 665290 145280 665530
rect 145520 665290 145610 665530
rect 145850 665290 145940 665530
rect 146180 665290 146290 665530
rect 146530 665290 146620 665530
rect 146860 665290 146950 665530
rect 147190 665290 147280 665530
rect 147520 665290 147630 665530
rect 147870 665290 147960 665530
rect 148200 665290 148290 665530
rect 148530 665290 148620 665530
rect 148860 665290 148970 665530
rect 149210 665290 149300 665530
rect 149540 665290 149630 665530
rect 149870 665290 149960 665530
rect 150200 665290 150310 665530
rect 150550 665290 150640 665530
rect 150880 665290 150970 665530
rect 151210 665290 151300 665530
rect 151540 665290 151650 665530
rect 151890 665290 151980 665530
rect 152220 665290 152310 665530
rect 152550 665290 152640 665530
rect 152880 665290 152990 665530
rect 153230 665290 153320 665530
rect 153560 665290 153650 665530
rect 153890 665290 153980 665530
rect 154220 665290 154330 665530
rect 154570 665290 154660 665530
rect 154900 665290 154990 665530
rect 155230 665290 155320 665530
rect 155560 665290 155670 665530
rect 155910 665290 155930 665530
rect 144930 665200 155930 665290
rect 144930 664960 144950 665200
rect 145190 664960 145280 665200
rect 145520 664960 145610 665200
rect 145850 664960 145940 665200
rect 146180 664960 146290 665200
rect 146530 664960 146620 665200
rect 146860 664960 146950 665200
rect 147190 664960 147280 665200
rect 147520 664960 147630 665200
rect 147870 664960 147960 665200
rect 148200 664960 148290 665200
rect 148530 664960 148620 665200
rect 148860 664960 148970 665200
rect 149210 664960 149300 665200
rect 149540 664960 149630 665200
rect 149870 664960 149960 665200
rect 150200 664960 150310 665200
rect 150550 664960 150640 665200
rect 150880 664960 150970 665200
rect 151210 664960 151300 665200
rect 151540 664960 151650 665200
rect 151890 664960 151980 665200
rect 152220 664960 152310 665200
rect 152550 664960 152640 665200
rect 152880 664960 152990 665200
rect 153230 664960 153320 665200
rect 153560 664960 153650 665200
rect 153890 664960 153980 665200
rect 154220 664960 154330 665200
rect 154570 664960 154660 665200
rect 154900 664960 154990 665200
rect 155230 664960 155320 665200
rect 155560 664960 155670 665200
rect 155910 664960 155930 665200
rect 144930 664850 155930 664960
rect 144930 664610 144950 664850
rect 145190 664610 145280 664850
rect 145520 664610 145610 664850
rect 145850 664610 145940 664850
rect 146180 664610 146290 664850
rect 146530 664610 146620 664850
rect 146860 664610 146950 664850
rect 147190 664610 147280 664850
rect 147520 664610 147630 664850
rect 147870 664610 147960 664850
rect 148200 664610 148290 664850
rect 148530 664610 148620 664850
rect 148860 664610 148970 664850
rect 149210 664610 149300 664850
rect 149540 664610 149630 664850
rect 149870 664610 149960 664850
rect 150200 664610 150310 664850
rect 150550 664610 150640 664850
rect 150880 664610 150970 664850
rect 151210 664610 151300 664850
rect 151540 664610 151650 664850
rect 151890 664610 151980 664850
rect 152220 664610 152310 664850
rect 152550 664610 152640 664850
rect 152880 664610 152990 664850
rect 153230 664610 153320 664850
rect 153560 664610 153650 664850
rect 153890 664610 153980 664850
rect 154220 664610 154330 664850
rect 154570 664610 154660 664850
rect 154900 664610 154990 664850
rect 155230 664610 155320 664850
rect 155560 664610 155670 664850
rect 155910 664610 155930 664850
rect 144930 664520 155930 664610
rect 144930 664280 144950 664520
rect 145190 664280 145280 664520
rect 145520 664280 145610 664520
rect 145850 664280 145940 664520
rect 146180 664280 146290 664520
rect 146530 664280 146620 664520
rect 146860 664280 146950 664520
rect 147190 664280 147280 664520
rect 147520 664280 147630 664520
rect 147870 664280 147960 664520
rect 148200 664280 148290 664520
rect 148530 664280 148620 664520
rect 148860 664280 148970 664520
rect 149210 664280 149300 664520
rect 149540 664280 149630 664520
rect 149870 664280 149960 664520
rect 150200 664280 150310 664520
rect 150550 664280 150640 664520
rect 150880 664280 150970 664520
rect 151210 664280 151300 664520
rect 151540 664280 151650 664520
rect 151890 664280 151980 664520
rect 152220 664280 152310 664520
rect 152550 664280 152640 664520
rect 152880 664280 152990 664520
rect 153230 664280 153320 664520
rect 153560 664280 153650 664520
rect 153890 664280 153980 664520
rect 154220 664280 154330 664520
rect 154570 664280 154660 664520
rect 154900 664280 154990 664520
rect 155230 664280 155320 664520
rect 155560 664280 155670 664520
rect 155910 664280 155930 664520
rect 144930 664190 155930 664280
rect 144930 663950 144950 664190
rect 145190 663950 145280 664190
rect 145520 663950 145610 664190
rect 145850 663950 145940 664190
rect 146180 663950 146290 664190
rect 146530 663950 146620 664190
rect 146860 663950 146950 664190
rect 147190 663950 147280 664190
rect 147520 663950 147630 664190
rect 147870 663950 147960 664190
rect 148200 663950 148290 664190
rect 148530 663950 148620 664190
rect 148860 663950 148970 664190
rect 149210 663950 149300 664190
rect 149540 663950 149630 664190
rect 149870 663950 149960 664190
rect 150200 663950 150310 664190
rect 150550 663950 150640 664190
rect 150880 663950 150970 664190
rect 151210 663950 151300 664190
rect 151540 663950 151650 664190
rect 151890 663950 151980 664190
rect 152220 663950 152310 664190
rect 152550 663950 152640 664190
rect 152880 663950 152990 664190
rect 153230 663950 153320 664190
rect 153560 663950 153650 664190
rect 153890 663950 153980 664190
rect 154220 663950 154330 664190
rect 154570 663950 154660 664190
rect 154900 663950 154990 664190
rect 155230 663950 155320 664190
rect 155560 663950 155670 664190
rect 155910 663950 155930 664190
rect 144930 663860 155930 663950
rect 144930 663620 144950 663860
rect 145190 663620 145280 663860
rect 145520 663620 145610 663860
rect 145850 663620 145940 663860
rect 146180 663620 146290 663860
rect 146530 663620 146620 663860
rect 146860 663620 146950 663860
rect 147190 663620 147280 663860
rect 147520 663620 147630 663860
rect 147870 663620 147960 663860
rect 148200 663620 148290 663860
rect 148530 663620 148620 663860
rect 148860 663620 148970 663860
rect 149210 663620 149300 663860
rect 149540 663620 149630 663860
rect 149870 663620 149960 663860
rect 150200 663620 150310 663860
rect 150550 663620 150640 663860
rect 150880 663620 150970 663860
rect 151210 663620 151300 663860
rect 151540 663620 151650 663860
rect 151890 663620 151980 663860
rect 152220 663620 152310 663860
rect 152550 663620 152640 663860
rect 152880 663620 152990 663860
rect 153230 663620 153320 663860
rect 153560 663620 153650 663860
rect 153890 663620 153980 663860
rect 154220 663620 154330 663860
rect 154570 663620 154660 663860
rect 154900 663620 154990 663860
rect 155230 663620 155320 663860
rect 155560 663620 155670 663860
rect 155910 663620 155930 663860
rect 144930 663510 155930 663620
rect 144930 663270 144950 663510
rect 145190 663270 145280 663510
rect 145520 663270 145610 663510
rect 145850 663270 145940 663510
rect 146180 663270 146290 663510
rect 146530 663270 146620 663510
rect 146860 663270 146950 663510
rect 147190 663270 147280 663510
rect 147520 663270 147630 663510
rect 147870 663270 147960 663510
rect 148200 663270 148290 663510
rect 148530 663270 148620 663510
rect 148860 663270 148970 663510
rect 149210 663270 149300 663510
rect 149540 663270 149630 663510
rect 149870 663270 149960 663510
rect 150200 663270 150310 663510
rect 150550 663270 150640 663510
rect 150880 663270 150970 663510
rect 151210 663270 151300 663510
rect 151540 663270 151650 663510
rect 151890 663270 151980 663510
rect 152220 663270 152310 663510
rect 152550 663270 152640 663510
rect 152880 663270 152990 663510
rect 153230 663270 153320 663510
rect 153560 663270 153650 663510
rect 153890 663270 153980 663510
rect 154220 663270 154330 663510
rect 154570 663270 154660 663510
rect 154900 663270 154990 663510
rect 155230 663270 155320 663510
rect 155560 663270 155670 663510
rect 155910 663270 155930 663510
rect 144930 663180 155930 663270
rect 144930 662940 144950 663180
rect 145190 662940 145280 663180
rect 145520 662940 145610 663180
rect 145850 662940 145940 663180
rect 146180 662940 146290 663180
rect 146530 662940 146620 663180
rect 146860 662940 146950 663180
rect 147190 662940 147280 663180
rect 147520 662940 147630 663180
rect 147870 662940 147960 663180
rect 148200 662940 148290 663180
rect 148530 662940 148620 663180
rect 148860 662940 148970 663180
rect 149210 662940 149300 663180
rect 149540 662940 149630 663180
rect 149870 662940 149960 663180
rect 150200 662940 150310 663180
rect 150550 662940 150640 663180
rect 150880 662940 150970 663180
rect 151210 662940 151300 663180
rect 151540 662940 151650 663180
rect 151890 662940 151980 663180
rect 152220 662940 152310 663180
rect 152550 662940 152640 663180
rect 152880 662940 152990 663180
rect 153230 662940 153320 663180
rect 153560 662940 153650 663180
rect 153890 662940 153980 663180
rect 154220 662940 154330 663180
rect 154570 662940 154660 663180
rect 154900 662940 154990 663180
rect 155230 662940 155320 663180
rect 155560 662940 155670 663180
rect 155910 662940 155930 663180
rect 144930 662850 155930 662940
rect 144930 662610 144950 662850
rect 145190 662610 145280 662850
rect 145520 662610 145610 662850
rect 145850 662610 145940 662850
rect 146180 662610 146290 662850
rect 146530 662610 146620 662850
rect 146860 662610 146950 662850
rect 147190 662610 147280 662850
rect 147520 662610 147630 662850
rect 147870 662610 147960 662850
rect 148200 662610 148290 662850
rect 148530 662610 148620 662850
rect 148860 662610 148970 662850
rect 149210 662610 149300 662850
rect 149540 662610 149630 662850
rect 149870 662610 149960 662850
rect 150200 662610 150310 662850
rect 150550 662610 150640 662850
rect 150880 662610 150970 662850
rect 151210 662610 151300 662850
rect 151540 662610 151650 662850
rect 151890 662610 151980 662850
rect 152220 662610 152310 662850
rect 152550 662610 152640 662850
rect 152880 662610 152990 662850
rect 153230 662610 153320 662850
rect 153560 662610 153650 662850
rect 153890 662610 153980 662850
rect 154220 662610 154330 662850
rect 154570 662610 154660 662850
rect 154900 662610 154990 662850
rect 155230 662610 155320 662850
rect 155560 662610 155670 662850
rect 155910 662610 155930 662850
rect 144930 662520 155930 662610
rect 144930 662280 144950 662520
rect 145190 662280 145280 662520
rect 145520 662280 145610 662520
rect 145850 662280 145940 662520
rect 146180 662280 146290 662520
rect 146530 662280 146620 662520
rect 146860 662280 146950 662520
rect 147190 662280 147280 662520
rect 147520 662280 147630 662520
rect 147870 662280 147960 662520
rect 148200 662280 148290 662520
rect 148530 662280 148620 662520
rect 148860 662280 148970 662520
rect 149210 662280 149300 662520
rect 149540 662280 149630 662520
rect 149870 662280 149960 662520
rect 150200 662280 150310 662520
rect 150550 662280 150640 662520
rect 150880 662280 150970 662520
rect 151210 662280 151300 662520
rect 151540 662280 151650 662520
rect 151890 662280 151980 662520
rect 152220 662280 152310 662520
rect 152550 662280 152640 662520
rect 152880 662280 152990 662520
rect 153230 662280 153320 662520
rect 153560 662280 153650 662520
rect 153890 662280 153980 662520
rect 154220 662280 154330 662520
rect 154570 662280 154660 662520
rect 154900 662280 154990 662520
rect 155230 662280 155320 662520
rect 155560 662280 155670 662520
rect 155910 662280 155930 662520
rect 144930 662170 155930 662280
rect 144930 661930 144950 662170
rect 145190 661930 145280 662170
rect 145520 661930 145610 662170
rect 145850 661930 145940 662170
rect 146180 661930 146290 662170
rect 146530 661930 146620 662170
rect 146860 661930 146950 662170
rect 147190 661930 147280 662170
rect 147520 661930 147630 662170
rect 147870 661930 147960 662170
rect 148200 661930 148290 662170
rect 148530 661930 148620 662170
rect 148860 661930 148970 662170
rect 149210 661930 149300 662170
rect 149540 661930 149630 662170
rect 149870 661930 149960 662170
rect 150200 661930 150310 662170
rect 150550 661930 150640 662170
rect 150880 661930 150970 662170
rect 151210 661930 151300 662170
rect 151540 661930 151650 662170
rect 151890 661930 151980 662170
rect 152220 661930 152310 662170
rect 152550 661930 152640 662170
rect 152880 661930 152990 662170
rect 153230 661930 153320 662170
rect 153560 661930 153650 662170
rect 153890 661930 153980 662170
rect 154220 661930 154330 662170
rect 154570 661930 154660 662170
rect 154900 661930 154990 662170
rect 155230 661930 155320 662170
rect 155560 661930 155670 662170
rect 155910 661930 155930 662170
rect 144930 661840 155930 661930
rect 144930 661600 144950 661840
rect 145190 661600 145280 661840
rect 145520 661600 145610 661840
rect 145850 661600 145940 661840
rect 146180 661600 146290 661840
rect 146530 661600 146620 661840
rect 146860 661600 146950 661840
rect 147190 661600 147280 661840
rect 147520 661600 147630 661840
rect 147870 661600 147960 661840
rect 148200 661600 148290 661840
rect 148530 661600 148620 661840
rect 148860 661600 148970 661840
rect 149210 661600 149300 661840
rect 149540 661600 149630 661840
rect 149870 661600 149960 661840
rect 150200 661600 150310 661840
rect 150550 661600 150640 661840
rect 150880 661600 150970 661840
rect 151210 661600 151300 661840
rect 151540 661600 151650 661840
rect 151890 661600 151980 661840
rect 152220 661600 152310 661840
rect 152550 661600 152640 661840
rect 152880 661600 152990 661840
rect 153230 661600 153320 661840
rect 153560 661600 153650 661840
rect 153890 661600 153980 661840
rect 154220 661600 154330 661840
rect 154570 661600 154660 661840
rect 154900 661600 154990 661840
rect 155230 661600 155320 661840
rect 155560 661600 155670 661840
rect 155910 661600 155930 661840
rect 144930 661510 155930 661600
rect 144930 661270 144950 661510
rect 145190 661270 145280 661510
rect 145520 661270 145610 661510
rect 145850 661270 145940 661510
rect 146180 661270 146290 661510
rect 146530 661270 146620 661510
rect 146860 661270 146950 661510
rect 147190 661270 147280 661510
rect 147520 661270 147630 661510
rect 147870 661270 147960 661510
rect 148200 661270 148290 661510
rect 148530 661270 148620 661510
rect 148860 661270 148970 661510
rect 149210 661270 149300 661510
rect 149540 661270 149630 661510
rect 149870 661270 149960 661510
rect 150200 661270 150310 661510
rect 150550 661270 150640 661510
rect 150880 661270 150970 661510
rect 151210 661270 151300 661510
rect 151540 661270 151650 661510
rect 151890 661270 151980 661510
rect 152220 661270 152310 661510
rect 152550 661270 152640 661510
rect 152880 661270 152990 661510
rect 153230 661270 153320 661510
rect 153560 661270 153650 661510
rect 153890 661270 153980 661510
rect 154220 661270 154330 661510
rect 154570 661270 154660 661510
rect 154900 661270 154990 661510
rect 155230 661270 155320 661510
rect 155560 661270 155670 661510
rect 155910 661270 155930 661510
rect 144930 661180 155930 661270
rect 144930 660940 144950 661180
rect 145190 660940 145280 661180
rect 145520 660940 145610 661180
rect 145850 660940 145940 661180
rect 146180 660940 146290 661180
rect 146530 660940 146620 661180
rect 146860 660940 146950 661180
rect 147190 660940 147280 661180
rect 147520 660940 147630 661180
rect 147870 660940 147960 661180
rect 148200 660940 148290 661180
rect 148530 660940 148620 661180
rect 148860 660940 148970 661180
rect 149210 660940 149300 661180
rect 149540 660940 149630 661180
rect 149870 660940 149960 661180
rect 150200 660940 150310 661180
rect 150550 660940 150640 661180
rect 150880 660940 150970 661180
rect 151210 660940 151300 661180
rect 151540 660940 151650 661180
rect 151890 660940 151980 661180
rect 152220 660940 152310 661180
rect 152550 660940 152640 661180
rect 152880 660940 152990 661180
rect 153230 660940 153320 661180
rect 153560 660940 153650 661180
rect 153890 660940 153980 661180
rect 154220 660940 154330 661180
rect 154570 660940 154660 661180
rect 154900 660940 154990 661180
rect 155230 660940 155320 661180
rect 155560 660940 155670 661180
rect 155910 660940 155930 661180
rect 144930 660920 155930 660940
rect 110790 660340 121790 660360
rect 110790 660100 110810 660340
rect 111050 660100 111160 660340
rect 111400 660100 111490 660340
rect 111730 660100 111820 660340
rect 112060 660100 112150 660340
rect 112390 660100 112500 660340
rect 112740 660100 112830 660340
rect 113070 660100 113160 660340
rect 113400 660100 113490 660340
rect 113730 660100 113840 660340
rect 114080 660100 114170 660340
rect 114410 660100 114500 660340
rect 114740 660100 114830 660340
rect 115070 660100 115180 660340
rect 115420 660100 115510 660340
rect 115750 660100 115840 660340
rect 116080 660100 116170 660340
rect 116410 660100 116520 660340
rect 116760 660100 116850 660340
rect 117090 660100 117180 660340
rect 117420 660100 117510 660340
rect 117750 660100 117860 660340
rect 118100 660100 118190 660340
rect 118430 660100 118520 660340
rect 118760 660100 118850 660340
rect 119090 660100 119200 660340
rect 119440 660100 119530 660340
rect 119770 660100 119860 660340
rect 120100 660100 120190 660340
rect 120430 660100 120540 660340
rect 120780 660100 120870 660340
rect 121110 660100 121200 660340
rect 121440 660100 121530 660340
rect 121770 660100 121790 660340
rect 110790 660010 121790 660100
rect 110790 659770 110810 660010
rect 111050 659770 111160 660010
rect 111400 659770 111490 660010
rect 111730 659770 111820 660010
rect 112060 659770 112150 660010
rect 112390 659770 112500 660010
rect 112740 659770 112830 660010
rect 113070 659770 113160 660010
rect 113400 659770 113490 660010
rect 113730 659770 113840 660010
rect 114080 659770 114170 660010
rect 114410 659770 114500 660010
rect 114740 659770 114830 660010
rect 115070 659770 115180 660010
rect 115420 659770 115510 660010
rect 115750 659770 115840 660010
rect 116080 659770 116170 660010
rect 116410 659770 116520 660010
rect 116760 659770 116850 660010
rect 117090 659770 117180 660010
rect 117420 659770 117510 660010
rect 117750 659770 117860 660010
rect 118100 659770 118190 660010
rect 118430 659770 118520 660010
rect 118760 659770 118850 660010
rect 119090 659770 119200 660010
rect 119440 659770 119530 660010
rect 119770 659770 119860 660010
rect 120100 659770 120190 660010
rect 120430 659770 120540 660010
rect 120780 659770 120870 660010
rect 121110 659770 121200 660010
rect 121440 659770 121530 660010
rect 121770 659770 121790 660010
rect 110790 659680 121790 659770
rect 110790 659440 110810 659680
rect 111050 659440 111160 659680
rect 111400 659440 111490 659680
rect 111730 659440 111820 659680
rect 112060 659440 112150 659680
rect 112390 659440 112500 659680
rect 112740 659440 112830 659680
rect 113070 659440 113160 659680
rect 113400 659440 113490 659680
rect 113730 659440 113840 659680
rect 114080 659440 114170 659680
rect 114410 659440 114500 659680
rect 114740 659440 114830 659680
rect 115070 659440 115180 659680
rect 115420 659440 115510 659680
rect 115750 659440 115840 659680
rect 116080 659440 116170 659680
rect 116410 659440 116520 659680
rect 116760 659440 116850 659680
rect 117090 659440 117180 659680
rect 117420 659440 117510 659680
rect 117750 659440 117860 659680
rect 118100 659440 118190 659680
rect 118430 659440 118520 659680
rect 118760 659440 118850 659680
rect 119090 659440 119200 659680
rect 119440 659440 119530 659680
rect 119770 659440 119860 659680
rect 120100 659440 120190 659680
rect 120430 659440 120540 659680
rect 120780 659440 120870 659680
rect 121110 659440 121200 659680
rect 121440 659440 121530 659680
rect 121770 659440 121790 659680
rect 110790 659350 121790 659440
rect 110790 659110 110810 659350
rect 111050 659110 111160 659350
rect 111400 659110 111490 659350
rect 111730 659110 111820 659350
rect 112060 659110 112150 659350
rect 112390 659110 112500 659350
rect 112740 659110 112830 659350
rect 113070 659110 113160 659350
rect 113400 659110 113490 659350
rect 113730 659110 113840 659350
rect 114080 659110 114170 659350
rect 114410 659110 114500 659350
rect 114740 659110 114830 659350
rect 115070 659110 115180 659350
rect 115420 659110 115510 659350
rect 115750 659110 115840 659350
rect 116080 659110 116170 659350
rect 116410 659110 116520 659350
rect 116760 659110 116850 659350
rect 117090 659110 117180 659350
rect 117420 659110 117510 659350
rect 117750 659110 117860 659350
rect 118100 659110 118190 659350
rect 118430 659110 118520 659350
rect 118760 659110 118850 659350
rect 119090 659110 119200 659350
rect 119440 659110 119530 659350
rect 119770 659110 119860 659350
rect 120100 659110 120190 659350
rect 120430 659110 120540 659350
rect 120780 659110 120870 659350
rect 121110 659110 121200 659350
rect 121440 659110 121530 659350
rect 121770 659110 121790 659350
rect 110790 659000 121790 659110
rect 110790 658760 110810 659000
rect 111050 658760 111160 659000
rect 111400 658760 111490 659000
rect 111730 658760 111820 659000
rect 112060 658760 112150 659000
rect 112390 658760 112500 659000
rect 112740 658760 112830 659000
rect 113070 658760 113160 659000
rect 113400 658760 113490 659000
rect 113730 658760 113840 659000
rect 114080 658760 114170 659000
rect 114410 658760 114500 659000
rect 114740 658760 114830 659000
rect 115070 658760 115180 659000
rect 115420 658760 115510 659000
rect 115750 658760 115840 659000
rect 116080 658760 116170 659000
rect 116410 658760 116520 659000
rect 116760 658760 116850 659000
rect 117090 658760 117180 659000
rect 117420 658760 117510 659000
rect 117750 658760 117860 659000
rect 118100 658760 118190 659000
rect 118430 658760 118520 659000
rect 118760 658760 118850 659000
rect 119090 658760 119200 659000
rect 119440 658760 119530 659000
rect 119770 658760 119860 659000
rect 120100 658760 120190 659000
rect 120430 658760 120540 659000
rect 120780 658760 120870 659000
rect 121110 658760 121200 659000
rect 121440 658760 121530 659000
rect 121770 658760 121790 659000
rect 110790 658670 121790 658760
rect 110790 658430 110810 658670
rect 111050 658430 111160 658670
rect 111400 658430 111490 658670
rect 111730 658430 111820 658670
rect 112060 658430 112150 658670
rect 112390 658430 112500 658670
rect 112740 658430 112830 658670
rect 113070 658430 113160 658670
rect 113400 658430 113490 658670
rect 113730 658430 113840 658670
rect 114080 658430 114170 658670
rect 114410 658430 114500 658670
rect 114740 658430 114830 658670
rect 115070 658430 115180 658670
rect 115420 658430 115510 658670
rect 115750 658430 115840 658670
rect 116080 658430 116170 658670
rect 116410 658430 116520 658670
rect 116760 658430 116850 658670
rect 117090 658430 117180 658670
rect 117420 658430 117510 658670
rect 117750 658430 117860 658670
rect 118100 658430 118190 658670
rect 118430 658430 118520 658670
rect 118760 658430 118850 658670
rect 119090 658430 119200 658670
rect 119440 658430 119530 658670
rect 119770 658430 119860 658670
rect 120100 658430 120190 658670
rect 120430 658430 120540 658670
rect 120780 658430 120870 658670
rect 121110 658430 121200 658670
rect 121440 658430 121530 658670
rect 121770 658430 121790 658670
rect 110790 658340 121790 658430
rect 110790 658100 110810 658340
rect 111050 658100 111160 658340
rect 111400 658100 111490 658340
rect 111730 658100 111820 658340
rect 112060 658100 112150 658340
rect 112390 658100 112500 658340
rect 112740 658100 112830 658340
rect 113070 658100 113160 658340
rect 113400 658100 113490 658340
rect 113730 658100 113840 658340
rect 114080 658100 114170 658340
rect 114410 658100 114500 658340
rect 114740 658100 114830 658340
rect 115070 658100 115180 658340
rect 115420 658100 115510 658340
rect 115750 658100 115840 658340
rect 116080 658100 116170 658340
rect 116410 658100 116520 658340
rect 116760 658100 116850 658340
rect 117090 658100 117180 658340
rect 117420 658100 117510 658340
rect 117750 658100 117860 658340
rect 118100 658100 118190 658340
rect 118430 658100 118520 658340
rect 118760 658100 118850 658340
rect 119090 658100 119200 658340
rect 119440 658100 119530 658340
rect 119770 658100 119860 658340
rect 120100 658100 120190 658340
rect 120430 658100 120540 658340
rect 120780 658100 120870 658340
rect 121110 658100 121200 658340
rect 121440 658100 121530 658340
rect 121770 658100 121790 658340
rect 110790 658010 121790 658100
rect 110790 657770 110810 658010
rect 111050 657770 111160 658010
rect 111400 657770 111490 658010
rect 111730 657770 111820 658010
rect 112060 657770 112150 658010
rect 112390 657770 112500 658010
rect 112740 657770 112830 658010
rect 113070 657770 113160 658010
rect 113400 657770 113490 658010
rect 113730 657770 113840 658010
rect 114080 657770 114170 658010
rect 114410 657770 114500 658010
rect 114740 657770 114830 658010
rect 115070 657770 115180 658010
rect 115420 657770 115510 658010
rect 115750 657770 115840 658010
rect 116080 657770 116170 658010
rect 116410 657770 116520 658010
rect 116760 657770 116850 658010
rect 117090 657770 117180 658010
rect 117420 657770 117510 658010
rect 117750 657770 117860 658010
rect 118100 657770 118190 658010
rect 118430 657770 118520 658010
rect 118760 657770 118850 658010
rect 119090 657770 119200 658010
rect 119440 657770 119530 658010
rect 119770 657770 119860 658010
rect 120100 657770 120190 658010
rect 120430 657770 120540 658010
rect 120780 657770 120870 658010
rect 121110 657770 121200 658010
rect 121440 657770 121530 658010
rect 121770 657770 121790 658010
rect 110790 657660 121790 657770
rect 110790 657420 110810 657660
rect 111050 657420 111160 657660
rect 111400 657420 111490 657660
rect 111730 657420 111820 657660
rect 112060 657420 112150 657660
rect 112390 657420 112500 657660
rect 112740 657420 112830 657660
rect 113070 657420 113160 657660
rect 113400 657420 113490 657660
rect 113730 657420 113840 657660
rect 114080 657420 114170 657660
rect 114410 657420 114500 657660
rect 114740 657420 114830 657660
rect 115070 657420 115180 657660
rect 115420 657420 115510 657660
rect 115750 657420 115840 657660
rect 116080 657420 116170 657660
rect 116410 657420 116520 657660
rect 116760 657420 116850 657660
rect 117090 657420 117180 657660
rect 117420 657420 117510 657660
rect 117750 657420 117860 657660
rect 118100 657420 118190 657660
rect 118430 657420 118520 657660
rect 118760 657420 118850 657660
rect 119090 657420 119200 657660
rect 119440 657420 119530 657660
rect 119770 657420 119860 657660
rect 120100 657420 120190 657660
rect 120430 657420 120540 657660
rect 120780 657420 120870 657660
rect 121110 657420 121200 657660
rect 121440 657420 121530 657660
rect 121770 657420 121790 657660
rect 110790 657330 121790 657420
rect 110790 657090 110810 657330
rect 111050 657090 111160 657330
rect 111400 657090 111490 657330
rect 111730 657090 111820 657330
rect 112060 657090 112150 657330
rect 112390 657090 112500 657330
rect 112740 657090 112830 657330
rect 113070 657090 113160 657330
rect 113400 657090 113490 657330
rect 113730 657090 113840 657330
rect 114080 657090 114170 657330
rect 114410 657090 114500 657330
rect 114740 657090 114830 657330
rect 115070 657090 115180 657330
rect 115420 657090 115510 657330
rect 115750 657090 115840 657330
rect 116080 657090 116170 657330
rect 116410 657090 116520 657330
rect 116760 657090 116850 657330
rect 117090 657090 117180 657330
rect 117420 657090 117510 657330
rect 117750 657090 117860 657330
rect 118100 657090 118190 657330
rect 118430 657090 118520 657330
rect 118760 657090 118850 657330
rect 119090 657090 119200 657330
rect 119440 657090 119530 657330
rect 119770 657090 119860 657330
rect 120100 657090 120190 657330
rect 120430 657090 120540 657330
rect 120780 657090 120870 657330
rect 121110 657090 121200 657330
rect 121440 657090 121530 657330
rect 121770 657090 121790 657330
rect 110790 657000 121790 657090
rect 110790 656760 110810 657000
rect 111050 656760 111160 657000
rect 111400 656760 111490 657000
rect 111730 656760 111820 657000
rect 112060 656760 112150 657000
rect 112390 656760 112500 657000
rect 112740 656760 112830 657000
rect 113070 656760 113160 657000
rect 113400 656760 113490 657000
rect 113730 656760 113840 657000
rect 114080 656760 114170 657000
rect 114410 656760 114500 657000
rect 114740 656760 114830 657000
rect 115070 656760 115180 657000
rect 115420 656760 115510 657000
rect 115750 656760 115840 657000
rect 116080 656760 116170 657000
rect 116410 656760 116520 657000
rect 116760 656760 116850 657000
rect 117090 656760 117180 657000
rect 117420 656760 117510 657000
rect 117750 656760 117860 657000
rect 118100 656760 118190 657000
rect 118430 656760 118520 657000
rect 118760 656760 118850 657000
rect 119090 656760 119200 657000
rect 119440 656760 119530 657000
rect 119770 656760 119860 657000
rect 120100 656760 120190 657000
rect 120430 656760 120540 657000
rect 120780 656760 120870 657000
rect 121110 656760 121200 657000
rect 121440 656760 121530 657000
rect 121770 656760 121790 657000
rect 110790 656670 121790 656760
rect 110790 656430 110810 656670
rect 111050 656430 111160 656670
rect 111400 656430 111490 656670
rect 111730 656430 111820 656670
rect 112060 656430 112150 656670
rect 112390 656430 112500 656670
rect 112740 656430 112830 656670
rect 113070 656430 113160 656670
rect 113400 656430 113490 656670
rect 113730 656430 113840 656670
rect 114080 656430 114170 656670
rect 114410 656430 114500 656670
rect 114740 656430 114830 656670
rect 115070 656430 115180 656670
rect 115420 656430 115510 656670
rect 115750 656430 115840 656670
rect 116080 656430 116170 656670
rect 116410 656430 116520 656670
rect 116760 656430 116850 656670
rect 117090 656430 117180 656670
rect 117420 656430 117510 656670
rect 117750 656430 117860 656670
rect 118100 656430 118190 656670
rect 118430 656430 118520 656670
rect 118760 656430 118850 656670
rect 119090 656430 119200 656670
rect 119440 656430 119530 656670
rect 119770 656430 119860 656670
rect 120100 656430 120190 656670
rect 120430 656430 120540 656670
rect 120780 656430 120870 656670
rect 121110 656430 121200 656670
rect 121440 656430 121530 656670
rect 121770 656430 121790 656670
rect 110790 656320 121790 656430
rect 110790 656080 110810 656320
rect 111050 656080 111160 656320
rect 111400 656080 111490 656320
rect 111730 656080 111820 656320
rect 112060 656080 112150 656320
rect 112390 656080 112500 656320
rect 112740 656080 112830 656320
rect 113070 656080 113160 656320
rect 113400 656080 113490 656320
rect 113730 656080 113840 656320
rect 114080 656080 114170 656320
rect 114410 656080 114500 656320
rect 114740 656080 114830 656320
rect 115070 656080 115180 656320
rect 115420 656080 115510 656320
rect 115750 656080 115840 656320
rect 116080 656080 116170 656320
rect 116410 656080 116520 656320
rect 116760 656080 116850 656320
rect 117090 656080 117180 656320
rect 117420 656080 117510 656320
rect 117750 656080 117860 656320
rect 118100 656080 118190 656320
rect 118430 656080 118520 656320
rect 118760 656080 118850 656320
rect 119090 656080 119200 656320
rect 119440 656080 119530 656320
rect 119770 656080 119860 656320
rect 120100 656080 120190 656320
rect 120430 656080 120540 656320
rect 120780 656080 120870 656320
rect 121110 656080 121200 656320
rect 121440 656080 121530 656320
rect 121770 656080 121790 656320
rect 110790 655990 121790 656080
rect 110790 655750 110810 655990
rect 111050 655750 111160 655990
rect 111400 655750 111490 655990
rect 111730 655750 111820 655990
rect 112060 655750 112150 655990
rect 112390 655750 112500 655990
rect 112740 655750 112830 655990
rect 113070 655750 113160 655990
rect 113400 655750 113490 655990
rect 113730 655750 113840 655990
rect 114080 655750 114170 655990
rect 114410 655750 114500 655990
rect 114740 655750 114830 655990
rect 115070 655750 115180 655990
rect 115420 655750 115510 655990
rect 115750 655750 115840 655990
rect 116080 655750 116170 655990
rect 116410 655750 116520 655990
rect 116760 655750 116850 655990
rect 117090 655750 117180 655990
rect 117420 655750 117510 655990
rect 117750 655750 117860 655990
rect 118100 655750 118190 655990
rect 118430 655750 118520 655990
rect 118760 655750 118850 655990
rect 119090 655750 119200 655990
rect 119440 655750 119530 655990
rect 119770 655750 119860 655990
rect 120100 655750 120190 655990
rect 120430 655750 120540 655990
rect 120780 655750 120870 655990
rect 121110 655750 121200 655990
rect 121440 655750 121530 655990
rect 121770 655750 121790 655990
rect 110790 655660 121790 655750
rect 110790 655420 110810 655660
rect 111050 655420 111160 655660
rect 111400 655420 111490 655660
rect 111730 655420 111820 655660
rect 112060 655420 112150 655660
rect 112390 655420 112500 655660
rect 112740 655420 112830 655660
rect 113070 655420 113160 655660
rect 113400 655420 113490 655660
rect 113730 655420 113840 655660
rect 114080 655420 114170 655660
rect 114410 655420 114500 655660
rect 114740 655420 114830 655660
rect 115070 655420 115180 655660
rect 115420 655420 115510 655660
rect 115750 655420 115840 655660
rect 116080 655420 116170 655660
rect 116410 655420 116520 655660
rect 116760 655420 116850 655660
rect 117090 655420 117180 655660
rect 117420 655420 117510 655660
rect 117750 655420 117860 655660
rect 118100 655420 118190 655660
rect 118430 655420 118520 655660
rect 118760 655420 118850 655660
rect 119090 655420 119200 655660
rect 119440 655420 119530 655660
rect 119770 655420 119860 655660
rect 120100 655420 120190 655660
rect 120430 655420 120540 655660
rect 120780 655420 120870 655660
rect 121110 655420 121200 655660
rect 121440 655420 121530 655660
rect 121770 655420 121790 655660
rect 110790 655330 121790 655420
rect 110790 655090 110810 655330
rect 111050 655090 111160 655330
rect 111400 655090 111490 655330
rect 111730 655090 111820 655330
rect 112060 655090 112150 655330
rect 112390 655090 112500 655330
rect 112740 655090 112830 655330
rect 113070 655090 113160 655330
rect 113400 655090 113490 655330
rect 113730 655090 113840 655330
rect 114080 655090 114170 655330
rect 114410 655090 114500 655330
rect 114740 655090 114830 655330
rect 115070 655090 115180 655330
rect 115420 655090 115510 655330
rect 115750 655090 115840 655330
rect 116080 655090 116170 655330
rect 116410 655090 116520 655330
rect 116760 655090 116850 655330
rect 117090 655090 117180 655330
rect 117420 655090 117510 655330
rect 117750 655090 117860 655330
rect 118100 655090 118190 655330
rect 118430 655090 118520 655330
rect 118760 655090 118850 655330
rect 119090 655090 119200 655330
rect 119440 655090 119530 655330
rect 119770 655090 119860 655330
rect 120100 655090 120190 655330
rect 120430 655090 120540 655330
rect 120780 655090 120870 655330
rect 121110 655090 121200 655330
rect 121440 655090 121530 655330
rect 121770 655090 121790 655330
rect 110790 654980 121790 655090
rect 110790 654740 110810 654980
rect 111050 654740 111160 654980
rect 111400 654740 111490 654980
rect 111730 654740 111820 654980
rect 112060 654740 112150 654980
rect 112390 654740 112500 654980
rect 112740 654740 112830 654980
rect 113070 654740 113160 654980
rect 113400 654740 113490 654980
rect 113730 654740 113840 654980
rect 114080 654740 114170 654980
rect 114410 654740 114500 654980
rect 114740 654740 114830 654980
rect 115070 654740 115180 654980
rect 115420 654740 115510 654980
rect 115750 654740 115840 654980
rect 116080 654740 116170 654980
rect 116410 654740 116520 654980
rect 116760 654740 116850 654980
rect 117090 654740 117180 654980
rect 117420 654740 117510 654980
rect 117750 654740 117860 654980
rect 118100 654740 118190 654980
rect 118430 654740 118520 654980
rect 118760 654740 118850 654980
rect 119090 654740 119200 654980
rect 119440 654740 119530 654980
rect 119770 654740 119860 654980
rect 120100 654740 120190 654980
rect 120430 654740 120540 654980
rect 120780 654740 120870 654980
rect 121110 654740 121200 654980
rect 121440 654740 121530 654980
rect 121770 654740 121790 654980
rect 110790 654650 121790 654740
rect 110790 654410 110810 654650
rect 111050 654410 111160 654650
rect 111400 654410 111490 654650
rect 111730 654410 111820 654650
rect 112060 654410 112150 654650
rect 112390 654410 112500 654650
rect 112740 654410 112830 654650
rect 113070 654410 113160 654650
rect 113400 654410 113490 654650
rect 113730 654410 113840 654650
rect 114080 654410 114170 654650
rect 114410 654410 114500 654650
rect 114740 654410 114830 654650
rect 115070 654410 115180 654650
rect 115420 654410 115510 654650
rect 115750 654410 115840 654650
rect 116080 654410 116170 654650
rect 116410 654410 116520 654650
rect 116760 654410 116850 654650
rect 117090 654410 117180 654650
rect 117420 654410 117510 654650
rect 117750 654410 117860 654650
rect 118100 654410 118190 654650
rect 118430 654410 118520 654650
rect 118760 654410 118850 654650
rect 119090 654410 119200 654650
rect 119440 654410 119530 654650
rect 119770 654410 119860 654650
rect 120100 654410 120190 654650
rect 120430 654410 120540 654650
rect 120780 654410 120870 654650
rect 121110 654410 121200 654650
rect 121440 654410 121530 654650
rect 121770 654410 121790 654650
rect 110790 654320 121790 654410
rect 110790 654080 110810 654320
rect 111050 654080 111160 654320
rect 111400 654080 111490 654320
rect 111730 654080 111820 654320
rect 112060 654080 112150 654320
rect 112390 654080 112500 654320
rect 112740 654080 112830 654320
rect 113070 654080 113160 654320
rect 113400 654080 113490 654320
rect 113730 654080 113840 654320
rect 114080 654080 114170 654320
rect 114410 654080 114500 654320
rect 114740 654080 114830 654320
rect 115070 654080 115180 654320
rect 115420 654080 115510 654320
rect 115750 654080 115840 654320
rect 116080 654080 116170 654320
rect 116410 654080 116520 654320
rect 116760 654080 116850 654320
rect 117090 654080 117180 654320
rect 117420 654080 117510 654320
rect 117750 654080 117860 654320
rect 118100 654080 118190 654320
rect 118430 654080 118520 654320
rect 118760 654080 118850 654320
rect 119090 654080 119200 654320
rect 119440 654080 119530 654320
rect 119770 654080 119860 654320
rect 120100 654080 120190 654320
rect 120430 654080 120540 654320
rect 120780 654080 120870 654320
rect 121110 654080 121200 654320
rect 121440 654080 121530 654320
rect 121770 654080 121790 654320
rect 110790 653990 121790 654080
rect 110790 653750 110810 653990
rect 111050 653750 111160 653990
rect 111400 653750 111490 653990
rect 111730 653750 111820 653990
rect 112060 653750 112150 653990
rect 112390 653750 112500 653990
rect 112740 653750 112830 653990
rect 113070 653750 113160 653990
rect 113400 653750 113490 653990
rect 113730 653750 113840 653990
rect 114080 653750 114170 653990
rect 114410 653750 114500 653990
rect 114740 653750 114830 653990
rect 115070 653750 115180 653990
rect 115420 653750 115510 653990
rect 115750 653750 115840 653990
rect 116080 653750 116170 653990
rect 116410 653750 116520 653990
rect 116760 653750 116850 653990
rect 117090 653750 117180 653990
rect 117420 653750 117510 653990
rect 117750 653750 117860 653990
rect 118100 653750 118190 653990
rect 118430 653750 118520 653990
rect 118760 653750 118850 653990
rect 119090 653750 119200 653990
rect 119440 653750 119530 653990
rect 119770 653750 119860 653990
rect 120100 653750 120190 653990
rect 120430 653750 120540 653990
rect 120780 653750 120870 653990
rect 121110 653750 121200 653990
rect 121440 653750 121530 653990
rect 121770 653750 121790 653990
rect 110790 653640 121790 653750
rect 110790 653400 110810 653640
rect 111050 653400 111160 653640
rect 111400 653400 111490 653640
rect 111730 653400 111820 653640
rect 112060 653400 112150 653640
rect 112390 653400 112500 653640
rect 112740 653400 112830 653640
rect 113070 653400 113160 653640
rect 113400 653400 113490 653640
rect 113730 653400 113840 653640
rect 114080 653400 114170 653640
rect 114410 653400 114500 653640
rect 114740 653400 114830 653640
rect 115070 653400 115180 653640
rect 115420 653400 115510 653640
rect 115750 653400 115840 653640
rect 116080 653400 116170 653640
rect 116410 653400 116520 653640
rect 116760 653400 116850 653640
rect 117090 653400 117180 653640
rect 117420 653400 117510 653640
rect 117750 653400 117860 653640
rect 118100 653400 118190 653640
rect 118430 653400 118520 653640
rect 118760 653400 118850 653640
rect 119090 653400 119200 653640
rect 119440 653400 119530 653640
rect 119770 653400 119860 653640
rect 120100 653400 120190 653640
rect 120430 653400 120540 653640
rect 120780 653400 120870 653640
rect 121110 653400 121200 653640
rect 121440 653400 121530 653640
rect 121770 653400 121790 653640
rect 110790 653310 121790 653400
rect 110790 653070 110810 653310
rect 111050 653070 111160 653310
rect 111400 653070 111490 653310
rect 111730 653070 111820 653310
rect 112060 653070 112150 653310
rect 112390 653070 112500 653310
rect 112740 653070 112830 653310
rect 113070 653070 113160 653310
rect 113400 653070 113490 653310
rect 113730 653070 113840 653310
rect 114080 653070 114170 653310
rect 114410 653070 114500 653310
rect 114740 653070 114830 653310
rect 115070 653070 115180 653310
rect 115420 653070 115510 653310
rect 115750 653070 115840 653310
rect 116080 653070 116170 653310
rect 116410 653070 116520 653310
rect 116760 653070 116850 653310
rect 117090 653070 117180 653310
rect 117420 653070 117510 653310
rect 117750 653070 117860 653310
rect 118100 653070 118190 653310
rect 118430 653070 118520 653310
rect 118760 653070 118850 653310
rect 119090 653070 119200 653310
rect 119440 653070 119530 653310
rect 119770 653070 119860 653310
rect 120100 653070 120190 653310
rect 120430 653070 120540 653310
rect 120780 653070 120870 653310
rect 121110 653070 121200 653310
rect 121440 653070 121530 653310
rect 121770 653070 121790 653310
rect 110790 652980 121790 653070
rect 110790 652740 110810 652980
rect 111050 652740 111160 652980
rect 111400 652740 111490 652980
rect 111730 652740 111820 652980
rect 112060 652740 112150 652980
rect 112390 652740 112500 652980
rect 112740 652740 112830 652980
rect 113070 652740 113160 652980
rect 113400 652740 113490 652980
rect 113730 652740 113840 652980
rect 114080 652740 114170 652980
rect 114410 652740 114500 652980
rect 114740 652740 114830 652980
rect 115070 652740 115180 652980
rect 115420 652740 115510 652980
rect 115750 652740 115840 652980
rect 116080 652740 116170 652980
rect 116410 652740 116520 652980
rect 116760 652740 116850 652980
rect 117090 652740 117180 652980
rect 117420 652740 117510 652980
rect 117750 652740 117860 652980
rect 118100 652740 118190 652980
rect 118430 652740 118520 652980
rect 118760 652740 118850 652980
rect 119090 652740 119200 652980
rect 119440 652740 119530 652980
rect 119770 652740 119860 652980
rect 120100 652740 120190 652980
rect 120430 652740 120540 652980
rect 120780 652740 120870 652980
rect 121110 652740 121200 652980
rect 121440 652740 121530 652980
rect 121770 652740 121790 652980
rect 110790 652650 121790 652740
rect 110790 652410 110810 652650
rect 111050 652410 111160 652650
rect 111400 652410 111490 652650
rect 111730 652410 111820 652650
rect 112060 652410 112150 652650
rect 112390 652410 112500 652650
rect 112740 652410 112830 652650
rect 113070 652410 113160 652650
rect 113400 652410 113490 652650
rect 113730 652410 113840 652650
rect 114080 652410 114170 652650
rect 114410 652410 114500 652650
rect 114740 652410 114830 652650
rect 115070 652410 115180 652650
rect 115420 652410 115510 652650
rect 115750 652410 115840 652650
rect 116080 652410 116170 652650
rect 116410 652410 116520 652650
rect 116760 652410 116850 652650
rect 117090 652410 117180 652650
rect 117420 652410 117510 652650
rect 117750 652410 117860 652650
rect 118100 652410 118190 652650
rect 118430 652410 118520 652650
rect 118760 652410 118850 652650
rect 119090 652410 119200 652650
rect 119440 652410 119530 652650
rect 119770 652410 119860 652650
rect 120100 652410 120190 652650
rect 120430 652410 120540 652650
rect 120780 652410 120870 652650
rect 121110 652410 121200 652650
rect 121440 652410 121530 652650
rect 121770 652410 121790 652650
rect 110790 652300 121790 652410
rect 110790 652060 110810 652300
rect 111050 652060 111160 652300
rect 111400 652060 111490 652300
rect 111730 652060 111820 652300
rect 112060 652060 112150 652300
rect 112390 652060 112500 652300
rect 112740 652060 112830 652300
rect 113070 652060 113160 652300
rect 113400 652060 113490 652300
rect 113730 652060 113840 652300
rect 114080 652060 114170 652300
rect 114410 652060 114500 652300
rect 114740 652060 114830 652300
rect 115070 652060 115180 652300
rect 115420 652060 115510 652300
rect 115750 652060 115840 652300
rect 116080 652060 116170 652300
rect 116410 652060 116520 652300
rect 116760 652060 116850 652300
rect 117090 652060 117180 652300
rect 117420 652060 117510 652300
rect 117750 652060 117860 652300
rect 118100 652060 118190 652300
rect 118430 652060 118520 652300
rect 118760 652060 118850 652300
rect 119090 652060 119200 652300
rect 119440 652060 119530 652300
rect 119770 652060 119860 652300
rect 120100 652060 120190 652300
rect 120430 652060 120540 652300
rect 120780 652060 120870 652300
rect 121110 652060 121200 652300
rect 121440 652060 121530 652300
rect 121770 652060 121790 652300
rect 110790 651970 121790 652060
rect 110790 651730 110810 651970
rect 111050 651730 111160 651970
rect 111400 651730 111490 651970
rect 111730 651730 111820 651970
rect 112060 651730 112150 651970
rect 112390 651730 112500 651970
rect 112740 651730 112830 651970
rect 113070 651730 113160 651970
rect 113400 651730 113490 651970
rect 113730 651730 113840 651970
rect 114080 651730 114170 651970
rect 114410 651730 114500 651970
rect 114740 651730 114830 651970
rect 115070 651730 115180 651970
rect 115420 651730 115510 651970
rect 115750 651730 115840 651970
rect 116080 651730 116170 651970
rect 116410 651730 116520 651970
rect 116760 651730 116850 651970
rect 117090 651730 117180 651970
rect 117420 651730 117510 651970
rect 117750 651730 117860 651970
rect 118100 651730 118190 651970
rect 118430 651730 118520 651970
rect 118760 651730 118850 651970
rect 119090 651730 119200 651970
rect 119440 651730 119530 651970
rect 119770 651730 119860 651970
rect 120100 651730 120190 651970
rect 120430 651730 120540 651970
rect 120780 651730 120870 651970
rect 121110 651730 121200 651970
rect 121440 651730 121530 651970
rect 121770 651730 121790 651970
rect 110790 651640 121790 651730
rect 110790 651400 110810 651640
rect 111050 651400 111160 651640
rect 111400 651400 111490 651640
rect 111730 651400 111820 651640
rect 112060 651400 112150 651640
rect 112390 651400 112500 651640
rect 112740 651400 112830 651640
rect 113070 651400 113160 651640
rect 113400 651400 113490 651640
rect 113730 651400 113840 651640
rect 114080 651400 114170 651640
rect 114410 651400 114500 651640
rect 114740 651400 114830 651640
rect 115070 651400 115180 651640
rect 115420 651400 115510 651640
rect 115750 651400 115840 651640
rect 116080 651400 116170 651640
rect 116410 651400 116520 651640
rect 116760 651400 116850 651640
rect 117090 651400 117180 651640
rect 117420 651400 117510 651640
rect 117750 651400 117860 651640
rect 118100 651400 118190 651640
rect 118430 651400 118520 651640
rect 118760 651400 118850 651640
rect 119090 651400 119200 651640
rect 119440 651400 119530 651640
rect 119770 651400 119860 651640
rect 120100 651400 120190 651640
rect 120430 651400 120540 651640
rect 120780 651400 120870 651640
rect 121110 651400 121200 651640
rect 121440 651400 121530 651640
rect 121770 651400 121790 651640
rect 110790 651310 121790 651400
rect 110790 651070 110810 651310
rect 111050 651070 111160 651310
rect 111400 651070 111490 651310
rect 111730 651070 111820 651310
rect 112060 651070 112150 651310
rect 112390 651070 112500 651310
rect 112740 651070 112830 651310
rect 113070 651070 113160 651310
rect 113400 651070 113490 651310
rect 113730 651070 113840 651310
rect 114080 651070 114170 651310
rect 114410 651070 114500 651310
rect 114740 651070 114830 651310
rect 115070 651070 115180 651310
rect 115420 651070 115510 651310
rect 115750 651070 115840 651310
rect 116080 651070 116170 651310
rect 116410 651070 116520 651310
rect 116760 651070 116850 651310
rect 117090 651070 117180 651310
rect 117420 651070 117510 651310
rect 117750 651070 117860 651310
rect 118100 651070 118190 651310
rect 118430 651070 118520 651310
rect 118760 651070 118850 651310
rect 119090 651070 119200 651310
rect 119440 651070 119530 651310
rect 119770 651070 119860 651310
rect 120100 651070 120190 651310
rect 120430 651070 120540 651310
rect 120780 651070 120870 651310
rect 121110 651070 121200 651310
rect 121440 651070 121530 651310
rect 121770 651070 121790 651310
rect 110790 650960 121790 651070
rect 110790 650720 110810 650960
rect 111050 650720 111160 650960
rect 111400 650720 111490 650960
rect 111730 650720 111820 650960
rect 112060 650720 112150 650960
rect 112390 650720 112500 650960
rect 112740 650720 112830 650960
rect 113070 650720 113160 650960
rect 113400 650720 113490 650960
rect 113730 650720 113840 650960
rect 114080 650720 114170 650960
rect 114410 650720 114500 650960
rect 114740 650720 114830 650960
rect 115070 650720 115180 650960
rect 115420 650720 115510 650960
rect 115750 650720 115840 650960
rect 116080 650720 116170 650960
rect 116410 650720 116520 650960
rect 116760 650720 116850 650960
rect 117090 650720 117180 650960
rect 117420 650720 117510 650960
rect 117750 650720 117860 650960
rect 118100 650720 118190 650960
rect 118430 650720 118520 650960
rect 118760 650720 118850 650960
rect 119090 650720 119200 650960
rect 119440 650720 119530 650960
rect 119770 650720 119860 650960
rect 120100 650720 120190 650960
rect 120430 650720 120540 650960
rect 120780 650720 120870 650960
rect 121110 650720 121200 650960
rect 121440 650720 121530 650960
rect 121770 650720 121790 650960
rect 110790 650630 121790 650720
rect 110790 650390 110810 650630
rect 111050 650390 111160 650630
rect 111400 650390 111490 650630
rect 111730 650390 111820 650630
rect 112060 650390 112150 650630
rect 112390 650390 112500 650630
rect 112740 650390 112830 650630
rect 113070 650390 113160 650630
rect 113400 650390 113490 650630
rect 113730 650390 113840 650630
rect 114080 650390 114170 650630
rect 114410 650390 114500 650630
rect 114740 650390 114830 650630
rect 115070 650390 115180 650630
rect 115420 650390 115510 650630
rect 115750 650390 115840 650630
rect 116080 650390 116170 650630
rect 116410 650390 116520 650630
rect 116760 650390 116850 650630
rect 117090 650390 117180 650630
rect 117420 650390 117510 650630
rect 117750 650390 117860 650630
rect 118100 650390 118190 650630
rect 118430 650390 118520 650630
rect 118760 650390 118850 650630
rect 119090 650390 119200 650630
rect 119440 650390 119530 650630
rect 119770 650390 119860 650630
rect 120100 650390 120190 650630
rect 120430 650390 120540 650630
rect 120780 650390 120870 650630
rect 121110 650390 121200 650630
rect 121440 650390 121530 650630
rect 121770 650390 121790 650630
rect 110790 650300 121790 650390
rect 110790 650060 110810 650300
rect 111050 650060 111160 650300
rect 111400 650060 111490 650300
rect 111730 650060 111820 650300
rect 112060 650060 112150 650300
rect 112390 650060 112500 650300
rect 112740 650060 112830 650300
rect 113070 650060 113160 650300
rect 113400 650060 113490 650300
rect 113730 650060 113840 650300
rect 114080 650060 114170 650300
rect 114410 650060 114500 650300
rect 114740 650060 114830 650300
rect 115070 650060 115180 650300
rect 115420 650060 115510 650300
rect 115750 650060 115840 650300
rect 116080 650060 116170 650300
rect 116410 650060 116520 650300
rect 116760 650060 116850 650300
rect 117090 650060 117180 650300
rect 117420 650060 117510 650300
rect 117750 650060 117860 650300
rect 118100 650060 118190 650300
rect 118430 650060 118520 650300
rect 118760 650060 118850 650300
rect 119090 650060 119200 650300
rect 119440 650060 119530 650300
rect 119770 650060 119860 650300
rect 120100 650060 120190 650300
rect 120430 650060 120540 650300
rect 120780 650060 120870 650300
rect 121110 650060 121200 650300
rect 121440 650060 121530 650300
rect 121770 650060 121790 650300
rect 110790 649970 121790 650060
rect 110790 649730 110810 649970
rect 111050 649730 111160 649970
rect 111400 649730 111490 649970
rect 111730 649730 111820 649970
rect 112060 649730 112150 649970
rect 112390 649730 112500 649970
rect 112740 649730 112830 649970
rect 113070 649730 113160 649970
rect 113400 649730 113490 649970
rect 113730 649730 113840 649970
rect 114080 649730 114170 649970
rect 114410 649730 114500 649970
rect 114740 649730 114830 649970
rect 115070 649730 115180 649970
rect 115420 649730 115510 649970
rect 115750 649730 115840 649970
rect 116080 649730 116170 649970
rect 116410 649730 116520 649970
rect 116760 649730 116850 649970
rect 117090 649730 117180 649970
rect 117420 649730 117510 649970
rect 117750 649730 117860 649970
rect 118100 649730 118190 649970
rect 118430 649730 118520 649970
rect 118760 649730 118850 649970
rect 119090 649730 119200 649970
rect 119440 649730 119530 649970
rect 119770 649730 119860 649970
rect 120100 649730 120190 649970
rect 120430 649730 120540 649970
rect 120780 649730 120870 649970
rect 121110 649730 121200 649970
rect 121440 649730 121530 649970
rect 121770 649730 121790 649970
rect 110790 649620 121790 649730
rect 110790 649380 110810 649620
rect 111050 649380 111160 649620
rect 111400 649380 111490 649620
rect 111730 649380 111820 649620
rect 112060 649380 112150 649620
rect 112390 649380 112500 649620
rect 112740 649380 112830 649620
rect 113070 649380 113160 649620
rect 113400 649380 113490 649620
rect 113730 649380 113840 649620
rect 114080 649380 114170 649620
rect 114410 649380 114500 649620
rect 114740 649380 114830 649620
rect 115070 649380 115180 649620
rect 115420 649380 115510 649620
rect 115750 649380 115840 649620
rect 116080 649380 116170 649620
rect 116410 649380 116520 649620
rect 116760 649380 116850 649620
rect 117090 649380 117180 649620
rect 117420 649380 117510 649620
rect 117750 649380 117860 649620
rect 118100 649380 118190 649620
rect 118430 649380 118520 649620
rect 118760 649380 118850 649620
rect 119090 649380 119200 649620
rect 119440 649380 119530 649620
rect 119770 649380 119860 649620
rect 120100 649380 120190 649620
rect 120430 649380 120540 649620
rect 120780 649380 120870 649620
rect 121110 649380 121200 649620
rect 121440 649380 121530 649620
rect 121770 649380 121790 649620
rect 110790 649360 121790 649380
rect 122170 660340 133170 660360
rect 122170 660100 122190 660340
rect 122430 660100 122540 660340
rect 122780 660100 122870 660340
rect 123110 660100 123200 660340
rect 123440 660100 123530 660340
rect 123770 660100 123880 660340
rect 124120 660100 124210 660340
rect 124450 660100 124540 660340
rect 124780 660100 124870 660340
rect 125110 660100 125220 660340
rect 125460 660100 125550 660340
rect 125790 660100 125880 660340
rect 126120 660100 126210 660340
rect 126450 660100 126560 660340
rect 126800 660100 126890 660340
rect 127130 660100 127220 660340
rect 127460 660100 127550 660340
rect 127790 660100 127900 660340
rect 128140 660100 128230 660340
rect 128470 660100 128560 660340
rect 128800 660100 128890 660340
rect 129130 660100 129240 660340
rect 129480 660100 129570 660340
rect 129810 660100 129900 660340
rect 130140 660100 130230 660340
rect 130470 660100 130580 660340
rect 130820 660100 130910 660340
rect 131150 660100 131240 660340
rect 131480 660100 131570 660340
rect 131810 660100 131920 660340
rect 132160 660100 132250 660340
rect 132490 660100 132580 660340
rect 132820 660100 132910 660340
rect 133150 660100 133170 660340
rect 122170 660010 133170 660100
rect 122170 659770 122190 660010
rect 122430 659770 122540 660010
rect 122780 659770 122870 660010
rect 123110 659770 123200 660010
rect 123440 659770 123530 660010
rect 123770 659770 123880 660010
rect 124120 659770 124210 660010
rect 124450 659770 124540 660010
rect 124780 659770 124870 660010
rect 125110 659770 125220 660010
rect 125460 659770 125550 660010
rect 125790 659770 125880 660010
rect 126120 659770 126210 660010
rect 126450 659770 126560 660010
rect 126800 659770 126890 660010
rect 127130 659770 127220 660010
rect 127460 659770 127550 660010
rect 127790 659770 127900 660010
rect 128140 659770 128230 660010
rect 128470 659770 128560 660010
rect 128800 659770 128890 660010
rect 129130 659770 129240 660010
rect 129480 659770 129570 660010
rect 129810 659770 129900 660010
rect 130140 659770 130230 660010
rect 130470 659770 130580 660010
rect 130820 659770 130910 660010
rect 131150 659770 131240 660010
rect 131480 659770 131570 660010
rect 131810 659770 131920 660010
rect 132160 659770 132250 660010
rect 132490 659770 132580 660010
rect 132820 659770 132910 660010
rect 133150 659770 133170 660010
rect 122170 659680 133170 659770
rect 122170 659440 122190 659680
rect 122430 659440 122540 659680
rect 122780 659440 122870 659680
rect 123110 659440 123200 659680
rect 123440 659440 123530 659680
rect 123770 659440 123880 659680
rect 124120 659440 124210 659680
rect 124450 659440 124540 659680
rect 124780 659440 124870 659680
rect 125110 659440 125220 659680
rect 125460 659440 125550 659680
rect 125790 659440 125880 659680
rect 126120 659440 126210 659680
rect 126450 659440 126560 659680
rect 126800 659440 126890 659680
rect 127130 659440 127220 659680
rect 127460 659440 127550 659680
rect 127790 659440 127900 659680
rect 128140 659440 128230 659680
rect 128470 659440 128560 659680
rect 128800 659440 128890 659680
rect 129130 659440 129240 659680
rect 129480 659440 129570 659680
rect 129810 659440 129900 659680
rect 130140 659440 130230 659680
rect 130470 659440 130580 659680
rect 130820 659440 130910 659680
rect 131150 659440 131240 659680
rect 131480 659440 131570 659680
rect 131810 659440 131920 659680
rect 132160 659440 132250 659680
rect 132490 659440 132580 659680
rect 132820 659440 132910 659680
rect 133150 659440 133170 659680
rect 122170 659350 133170 659440
rect 122170 659110 122190 659350
rect 122430 659110 122540 659350
rect 122780 659110 122870 659350
rect 123110 659110 123200 659350
rect 123440 659110 123530 659350
rect 123770 659110 123880 659350
rect 124120 659110 124210 659350
rect 124450 659110 124540 659350
rect 124780 659110 124870 659350
rect 125110 659110 125220 659350
rect 125460 659110 125550 659350
rect 125790 659110 125880 659350
rect 126120 659110 126210 659350
rect 126450 659110 126560 659350
rect 126800 659110 126890 659350
rect 127130 659110 127220 659350
rect 127460 659110 127550 659350
rect 127790 659110 127900 659350
rect 128140 659110 128230 659350
rect 128470 659110 128560 659350
rect 128800 659110 128890 659350
rect 129130 659110 129240 659350
rect 129480 659110 129570 659350
rect 129810 659110 129900 659350
rect 130140 659110 130230 659350
rect 130470 659110 130580 659350
rect 130820 659110 130910 659350
rect 131150 659110 131240 659350
rect 131480 659110 131570 659350
rect 131810 659110 131920 659350
rect 132160 659110 132250 659350
rect 132490 659110 132580 659350
rect 132820 659110 132910 659350
rect 133150 659110 133170 659350
rect 122170 659000 133170 659110
rect 122170 658760 122190 659000
rect 122430 658760 122540 659000
rect 122780 658760 122870 659000
rect 123110 658760 123200 659000
rect 123440 658760 123530 659000
rect 123770 658760 123880 659000
rect 124120 658760 124210 659000
rect 124450 658760 124540 659000
rect 124780 658760 124870 659000
rect 125110 658760 125220 659000
rect 125460 658760 125550 659000
rect 125790 658760 125880 659000
rect 126120 658760 126210 659000
rect 126450 658760 126560 659000
rect 126800 658760 126890 659000
rect 127130 658760 127220 659000
rect 127460 658760 127550 659000
rect 127790 658760 127900 659000
rect 128140 658760 128230 659000
rect 128470 658760 128560 659000
rect 128800 658760 128890 659000
rect 129130 658760 129240 659000
rect 129480 658760 129570 659000
rect 129810 658760 129900 659000
rect 130140 658760 130230 659000
rect 130470 658760 130580 659000
rect 130820 658760 130910 659000
rect 131150 658760 131240 659000
rect 131480 658760 131570 659000
rect 131810 658760 131920 659000
rect 132160 658760 132250 659000
rect 132490 658760 132580 659000
rect 132820 658760 132910 659000
rect 133150 658760 133170 659000
rect 122170 658670 133170 658760
rect 122170 658430 122190 658670
rect 122430 658430 122540 658670
rect 122780 658430 122870 658670
rect 123110 658430 123200 658670
rect 123440 658430 123530 658670
rect 123770 658430 123880 658670
rect 124120 658430 124210 658670
rect 124450 658430 124540 658670
rect 124780 658430 124870 658670
rect 125110 658430 125220 658670
rect 125460 658430 125550 658670
rect 125790 658430 125880 658670
rect 126120 658430 126210 658670
rect 126450 658430 126560 658670
rect 126800 658430 126890 658670
rect 127130 658430 127220 658670
rect 127460 658430 127550 658670
rect 127790 658430 127900 658670
rect 128140 658430 128230 658670
rect 128470 658430 128560 658670
rect 128800 658430 128890 658670
rect 129130 658430 129240 658670
rect 129480 658430 129570 658670
rect 129810 658430 129900 658670
rect 130140 658430 130230 658670
rect 130470 658430 130580 658670
rect 130820 658430 130910 658670
rect 131150 658430 131240 658670
rect 131480 658430 131570 658670
rect 131810 658430 131920 658670
rect 132160 658430 132250 658670
rect 132490 658430 132580 658670
rect 132820 658430 132910 658670
rect 133150 658430 133170 658670
rect 122170 658340 133170 658430
rect 122170 658100 122190 658340
rect 122430 658100 122540 658340
rect 122780 658100 122870 658340
rect 123110 658100 123200 658340
rect 123440 658100 123530 658340
rect 123770 658100 123880 658340
rect 124120 658100 124210 658340
rect 124450 658100 124540 658340
rect 124780 658100 124870 658340
rect 125110 658100 125220 658340
rect 125460 658100 125550 658340
rect 125790 658100 125880 658340
rect 126120 658100 126210 658340
rect 126450 658100 126560 658340
rect 126800 658100 126890 658340
rect 127130 658100 127220 658340
rect 127460 658100 127550 658340
rect 127790 658100 127900 658340
rect 128140 658100 128230 658340
rect 128470 658100 128560 658340
rect 128800 658100 128890 658340
rect 129130 658100 129240 658340
rect 129480 658100 129570 658340
rect 129810 658100 129900 658340
rect 130140 658100 130230 658340
rect 130470 658100 130580 658340
rect 130820 658100 130910 658340
rect 131150 658100 131240 658340
rect 131480 658100 131570 658340
rect 131810 658100 131920 658340
rect 132160 658100 132250 658340
rect 132490 658100 132580 658340
rect 132820 658100 132910 658340
rect 133150 658100 133170 658340
rect 122170 658010 133170 658100
rect 122170 657770 122190 658010
rect 122430 657770 122540 658010
rect 122780 657770 122870 658010
rect 123110 657770 123200 658010
rect 123440 657770 123530 658010
rect 123770 657770 123880 658010
rect 124120 657770 124210 658010
rect 124450 657770 124540 658010
rect 124780 657770 124870 658010
rect 125110 657770 125220 658010
rect 125460 657770 125550 658010
rect 125790 657770 125880 658010
rect 126120 657770 126210 658010
rect 126450 657770 126560 658010
rect 126800 657770 126890 658010
rect 127130 657770 127220 658010
rect 127460 657770 127550 658010
rect 127790 657770 127900 658010
rect 128140 657770 128230 658010
rect 128470 657770 128560 658010
rect 128800 657770 128890 658010
rect 129130 657770 129240 658010
rect 129480 657770 129570 658010
rect 129810 657770 129900 658010
rect 130140 657770 130230 658010
rect 130470 657770 130580 658010
rect 130820 657770 130910 658010
rect 131150 657770 131240 658010
rect 131480 657770 131570 658010
rect 131810 657770 131920 658010
rect 132160 657770 132250 658010
rect 132490 657770 132580 658010
rect 132820 657770 132910 658010
rect 133150 657770 133170 658010
rect 122170 657660 133170 657770
rect 122170 657420 122190 657660
rect 122430 657420 122540 657660
rect 122780 657420 122870 657660
rect 123110 657420 123200 657660
rect 123440 657420 123530 657660
rect 123770 657420 123880 657660
rect 124120 657420 124210 657660
rect 124450 657420 124540 657660
rect 124780 657420 124870 657660
rect 125110 657420 125220 657660
rect 125460 657420 125550 657660
rect 125790 657420 125880 657660
rect 126120 657420 126210 657660
rect 126450 657420 126560 657660
rect 126800 657420 126890 657660
rect 127130 657420 127220 657660
rect 127460 657420 127550 657660
rect 127790 657420 127900 657660
rect 128140 657420 128230 657660
rect 128470 657420 128560 657660
rect 128800 657420 128890 657660
rect 129130 657420 129240 657660
rect 129480 657420 129570 657660
rect 129810 657420 129900 657660
rect 130140 657420 130230 657660
rect 130470 657420 130580 657660
rect 130820 657420 130910 657660
rect 131150 657420 131240 657660
rect 131480 657420 131570 657660
rect 131810 657420 131920 657660
rect 132160 657420 132250 657660
rect 132490 657420 132580 657660
rect 132820 657420 132910 657660
rect 133150 657420 133170 657660
rect 122170 657330 133170 657420
rect 122170 657090 122190 657330
rect 122430 657090 122540 657330
rect 122780 657090 122870 657330
rect 123110 657090 123200 657330
rect 123440 657090 123530 657330
rect 123770 657090 123880 657330
rect 124120 657090 124210 657330
rect 124450 657090 124540 657330
rect 124780 657090 124870 657330
rect 125110 657090 125220 657330
rect 125460 657090 125550 657330
rect 125790 657090 125880 657330
rect 126120 657090 126210 657330
rect 126450 657090 126560 657330
rect 126800 657090 126890 657330
rect 127130 657090 127220 657330
rect 127460 657090 127550 657330
rect 127790 657090 127900 657330
rect 128140 657090 128230 657330
rect 128470 657090 128560 657330
rect 128800 657090 128890 657330
rect 129130 657090 129240 657330
rect 129480 657090 129570 657330
rect 129810 657090 129900 657330
rect 130140 657090 130230 657330
rect 130470 657090 130580 657330
rect 130820 657090 130910 657330
rect 131150 657090 131240 657330
rect 131480 657090 131570 657330
rect 131810 657090 131920 657330
rect 132160 657090 132250 657330
rect 132490 657090 132580 657330
rect 132820 657090 132910 657330
rect 133150 657090 133170 657330
rect 122170 657000 133170 657090
rect 122170 656760 122190 657000
rect 122430 656760 122540 657000
rect 122780 656760 122870 657000
rect 123110 656760 123200 657000
rect 123440 656760 123530 657000
rect 123770 656760 123880 657000
rect 124120 656760 124210 657000
rect 124450 656760 124540 657000
rect 124780 656760 124870 657000
rect 125110 656760 125220 657000
rect 125460 656760 125550 657000
rect 125790 656760 125880 657000
rect 126120 656760 126210 657000
rect 126450 656760 126560 657000
rect 126800 656760 126890 657000
rect 127130 656760 127220 657000
rect 127460 656760 127550 657000
rect 127790 656760 127900 657000
rect 128140 656760 128230 657000
rect 128470 656760 128560 657000
rect 128800 656760 128890 657000
rect 129130 656760 129240 657000
rect 129480 656760 129570 657000
rect 129810 656760 129900 657000
rect 130140 656760 130230 657000
rect 130470 656760 130580 657000
rect 130820 656760 130910 657000
rect 131150 656760 131240 657000
rect 131480 656760 131570 657000
rect 131810 656760 131920 657000
rect 132160 656760 132250 657000
rect 132490 656760 132580 657000
rect 132820 656760 132910 657000
rect 133150 656760 133170 657000
rect 122170 656670 133170 656760
rect 122170 656430 122190 656670
rect 122430 656430 122540 656670
rect 122780 656430 122870 656670
rect 123110 656430 123200 656670
rect 123440 656430 123530 656670
rect 123770 656430 123880 656670
rect 124120 656430 124210 656670
rect 124450 656430 124540 656670
rect 124780 656430 124870 656670
rect 125110 656430 125220 656670
rect 125460 656430 125550 656670
rect 125790 656430 125880 656670
rect 126120 656430 126210 656670
rect 126450 656430 126560 656670
rect 126800 656430 126890 656670
rect 127130 656430 127220 656670
rect 127460 656430 127550 656670
rect 127790 656430 127900 656670
rect 128140 656430 128230 656670
rect 128470 656430 128560 656670
rect 128800 656430 128890 656670
rect 129130 656430 129240 656670
rect 129480 656430 129570 656670
rect 129810 656430 129900 656670
rect 130140 656430 130230 656670
rect 130470 656430 130580 656670
rect 130820 656430 130910 656670
rect 131150 656430 131240 656670
rect 131480 656430 131570 656670
rect 131810 656430 131920 656670
rect 132160 656430 132250 656670
rect 132490 656430 132580 656670
rect 132820 656430 132910 656670
rect 133150 656430 133170 656670
rect 122170 656320 133170 656430
rect 122170 656080 122190 656320
rect 122430 656080 122540 656320
rect 122780 656080 122870 656320
rect 123110 656080 123200 656320
rect 123440 656080 123530 656320
rect 123770 656080 123880 656320
rect 124120 656080 124210 656320
rect 124450 656080 124540 656320
rect 124780 656080 124870 656320
rect 125110 656080 125220 656320
rect 125460 656080 125550 656320
rect 125790 656080 125880 656320
rect 126120 656080 126210 656320
rect 126450 656080 126560 656320
rect 126800 656080 126890 656320
rect 127130 656080 127220 656320
rect 127460 656080 127550 656320
rect 127790 656080 127900 656320
rect 128140 656080 128230 656320
rect 128470 656080 128560 656320
rect 128800 656080 128890 656320
rect 129130 656080 129240 656320
rect 129480 656080 129570 656320
rect 129810 656080 129900 656320
rect 130140 656080 130230 656320
rect 130470 656080 130580 656320
rect 130820 656080 130910 656320
rect 131150 656080 131240 656320
rect 131480 656080 131570 656320
rect 131810 656080 131920 656320
rect 132160 656080 132250 656320
rect 132490 656080 132580 656320
rect 132820 656080 132910 656320
rect 133150 656080 133170 656320
rect 122170 655990 133170 656080
rect 122170 655750 122190 655990
rect 122430 655750 122540 655990
rect 122780 655750 122870 655990
rect 123110 655750 123200 655990
rect 123440 655750 123530 655990
rect 123770 655750 123880 655990
rect 124120 655750 124210 655990
rect 124450 655750 124540 655990
rect 124780 655750 124870 655990
rect 125110 655750 125220 655990
rect 125460 655750 125550 655990
rect 125790 655750 125880 655990
rect 126120 655750 126210 655990
rect 126450 655750 126560 655990
rect 126800 655750 126890 655990
rect 127130 655750 127220 655990
rect 127460 655750 127550 655990
rect 127790 655750 127900 655990
rect 128140 655750 128230 655990
rect 128470 655750 128560 655990
rect 128800 655750 128890 655990
rect 129130 655750 129240 655990
rect 129480 655750 129570 655990
rect 129810 655750 129900 655990
rect 130140 655750 130230 655990
rect 130470 655750 130580 655990
rect 130820 655750 130910 655990
rect 131150 655750 131240 655990
rect 131480 655750 131570 655990
rect 131810 655750 131920 655990
rect 132160 655750 132250 655990
rect 132490 655750 132580 655990
rect 132820 655750 132910 655990
rect 133150 655750 133170 655990
rect 122170 655660 133170 655750
rect 122170 655420 122190 655660
rect 122430 655420 122540 655660
rect 122780 655420 122870 655660
rect 123110 655420 123200 655660
rect 123440 655420 123530 655660
rect 123770 655420 123880 655660
rect 124120 655420 124210 655660
rect 124450 655420 124540 655660
rect 124780 655420 124870 655660
rect 125110 655420 125220 655660
rect 125460 655420 125550 655660
rect 125790 655420 125880 655660
rect 126120 655420 126210 655660
rect 126450 655420 126560 655660
rect 126800 655420 126890 655660
rect 127130 655420 127220 655660
rect 127460 655420 127550 655660
rect 127790 655420 127900 655660
rect 128140 655420 128230 655660
rect 128470 655420 128560 655660
rect 128800 655420 128890 655660
rect 129130 655420 129240 655660
rect 129480 655420 129570 655660
rect 129810 655420 129900 655660
rect 130140 655420 130230 655660
rect 130470 655420 130580 655660
rect 130820 655420 130910 655660
rect 131150 655420 131240 655660
rect 131480 655420 131570 655660
rect 131810 655420 131920 655660
rect 132160 655420 132250 655660
rect 132490 655420 132580 655660
rect 132820 655420 132910 655660
rect 133150 655420 133170 655660
rect 122170 655330 133170 655420
rect 122170 655090 122190 655330
rect 122430 655090 122540 655330
rect 122780 655090 122870 655330
rect 123110 655090 123200 655330
rect 123440 655090 123530 655330
rect 123770 655090 123880 655330
rect 124120 655090 124210 655330
rect 124450 655090 124540 655330
rect 124780 655090 124870 655330
rect 125110 655090 125220 655330
rect 125460 655090 125550 655330
rect 125790 655090 125880 655330
rect 126120 655090 126210 655330
rect 126450 655090 126560 655330
rect 126800 655090 126890 655330
rect 127130 655090 127220 655330
rect 127460 655090 127550 655330
rect 127790 655090 127900 655330
rect 128140 655090 128230 655330
rect 128470 655090 128560 655330
rect 128800 655090 128890 655330
rect 129130 655090 129240 655330
rect 129480 655090 129570 655330
rect 129810 655090 129900 655330
rect 130140 655090 130230 655330
rect 130470 655090 130580 655330
rect 130820 655090 130910 655330
rect 131150 655090 131240 655330
rect 131480 655090 131570 655330
rect 131810 655090 131920 655330
rect 132160 655090 132250 655330
rect 132490 655090 132580 655330
rect 132820 655090 132910 655330
rect 133150 655090 133170 655330
rect 122170 654980 133170 655090
rect 122170 654740 122190 654980
rect 122430 654740 122540 654980
rect 122780 654740 122870 654980
rect 123110 654740 123200 654980
rect 123440 654740 123530 654980
rect 123770 654740 123880 654980
rect 124120 654740 124210 654980
rect 124450 654740 124540 654980
rect 124780 654740 124870 654980
rect 125110 654740 125220 654980
rect 125460 654740 125550 654980
rect 125790 654740 125880 654980
rect 126120 654740 126210 654980
rect 126450 654740 126560 654980
rect 126800 654740 126890 654980
rect 127130 654740 127220 654980
rect 127460 654740 127550 654980
rect 127790 654740 127900 654980
rect 128140 654740 128230 654980
rect 128470 654740 128560 654980
rect 128800 654740 128890 654980
rect 129130 654740 129240 654980
rect 129480 654740 129570 654980
rect 129810 654740 129900 654980
rect 130140 654740 130230 654980
rect 130470 654740 130580 654980
rect 130820 654740 130910 654980
rect 131150 654740 131240 654980
rect 131480 654740 131570 654980
rect 131810 654740 131920 654980
rect 132160 654740 132250 654980
rect 132490 654740 132580 654980
rect 132820 654740 132910 654980
rect 133150 654740 133170 654980
rect 122170 654650 133170 654740
rect 122170 654410 122190 654650
rect 122430 654410 122540 654650
rect 122780 654410 122870 654650
rect 123110 654410 123200 654650
rect 123440 654410 123530 654650
rect 123770 654410 123880 654650
rect 124120 654410 124210 654650
rect 124450 654410 124540 654650
rect 124780 654410 124870 654650
rect 125110 654410 125220 654650
rect 125460 654410 125550 654650
rect 125790 654410 125880 654650
rect 126120 654410 126210 654650
rect 126450 654410 126560 654650
rect 126800 654410 126890 654650
rect 127130 654410 127220 654650
rect 127460 654410 127550 654650
rect 127790 654410 127900 654650
rect 128140 654410 128230 654650
rect 128470 654410 128560 654650
rect 128800 654410 128890 654650
rect 129130 654410 129240 654650
rect 129480 654410 129570 654650
rect 129810 654410 129900 654650
rect 130140 654410 130230 654650
rect 130470 654410 130580 654650
rect 130820 654410 130910 654650
rect 131150 654410 131240 654650
rect 131480 654410 131570 654650
rect 131810 654410 131920 654650
rect 132160 654410 132250 654650
rect 132490 654410 132580 654650
rect 132820 654410 132910 654650
rect 133150 654410 133170 654650
rect 122170 654320 133170 654410
rect 122170 654080 122190 654320
rect 122430 654080 122540 654320
rect 122780 654080 122870 654320
rect 123110 654080 123200 654320
rect 123440 654080 123530 654320
rect 123770 654080 123880 654320
rect 124120 654080 124210 654320
rect 124450 654080 124540 654320
rect 124780 654080 124870 654320
rect 125110 654080 125220 654320
rect 125460 654080 125550 654320
rect 125790 654080 125880 654320
rect 126120 654080 126210 654320
rect 126450 654080 126560 654320
rect 126800 654080 126890 654320
rect 127130 654080 127220 654320
rect 127460 654080 127550 654320
rect 127790 654080 127900 654320
rect 128140 654080 128230 654320
rect 128470 654080 128560 654320
rect 128800 654080 128890 654320
rect 129130 654080 129240 654320
rect 129480 654080 129570 654320
rect 129810 654080 129900 654320
rect 130140 654080 130230 654320
rect 130470 654080 130580 654320
rect 130820 654080 130910 654320
rect 131150 654080 131240 654320
rect 131480 654080 131570 654320
rect 131810 654080 131920 654320
rect 132160 654080 132250 654320
rect 132490 654080 132580 654320
rect 132820 654080 132910 654320
rect 133150 654080 133170 654320
rect 122170 653990 133170 654080
rect 122170 653750 122190 653990
rect 122430 653750 122540 653990
rect 122780 653750 122870 653990
rect 123110 653750 123200 653990
rect 123440 653750 123530 653990
rect 123770 653750 123880 653990
rect 124120 653750 124210 653990
rect 124450 653750 124540 653990
rect 124780 653750 124870 653990
rect 125110 653750 125220 653990
rect 125460 653750 125550 653990
rect 125790 653750 125880 653990
rect 126120 653750 126210 653990
rect 126450 653750 126560 653990
rect 126800 653750 126890 653990
rect 127130 653750 127220 653990
rect 127460 653750 127550 653990
rect 127790 653750 127900 653990
rect 128140 653750 128230 653990
rect 128470 653750 128560 653990
rect 128800 653750 128890 653990
rect 129130 653750 129240 653990
rect 129480 653750 129570 653990
rect 129810 653750 129900 653990
rect 130140 653750 130230 653990
rect 130470 653750 130580 653990
rect 130820 653750 130910 653990
rect 131150 653750 131240 653990
rect 131480 653750 131570 653990
rect 131810 653750 131920 653990
rect 132160 653750 132250 653990
rect 132490 653750 132580 653990
rect 132820 653750 132910 653990
rect 133150 653750 133170 653990
rect 122170 653640 133170 653750
rect 122170 653400 122190 653640
rect 122430 653400 122540 653640
rect 122780 653400 122870 653640
rect 123110 653400 123200 653640
rect 123440 653400 123530 653640
rect 123770 653400 123880 653640
rect 124120 653400 124210 653640
rect 124450 653400 124540 653640
rect 124780 653400 124870 653640
rect 125110 653400 125220 653640
rect 125460 653400 125550 653640
rect 125790 653400 125880 653640
rect 126120 653400 126210 653640
rect 126450 653400 126560 653640
rect 126800 653400 126890 653640
rect 127130 653400 127220 653640
rect 127460 653400 127550 653640
rect 127790 653400 127900 653640
rect 128140 653400 128230 653640
rect 128470 653400 128560 653640
rect 128800 653400 128890 653640
rect 129130 653400 129240 653640
rect 129480 653400 129570 653640
rect 129810 653400 129900 653640
rect 130140 653400 130230 653640
rect 130470 653400 130580 653640
rect 130820 653400 130910 653640
rect 131150 653400 131240 653640
rect 131480 653400 131570 653640
rect 131810 653400 131920 653640
rect 132160 653400 132250 653640
rect 132490 653400 132580 653640
rect 132820 653400 132910 653640
rect 133150 653400 133170 653640
rect 122170 653310 133170 653400
rect 122170 653070 122190 653310
rect 122430 653070 122540 653310
rect 122780 653070 122870 653310
rect 123110 653070 123200 653310
rect 123440 653070 123530 653310
rect 123770 653070 123880 653310
rect 124120 653070 124210 653310
rect 124450 653070 124540 653310
rect 124780 653070 124870 653310
rect 125110 653070 125220 653310
rect 125460 653070 125550 653310
rect 125790 653070 125880 653310
rect 126120 653070 126210 653310
rect 126450 653070 126560 653310
rect 126800 653070 126890 653310
rect 127130 653070 127220 653310
rect 127460 653070 127550 653310
rect 127790 653070 127900 653310
rect 128140 653070 128230 653310
rect 128470 653070 128560 653310
rect 128800 653070 128890 653310
rect 129130 653070 129240 653310
rect 129480 653070 129570 653310
rect 129810 653070 129900 653310
rect 130140 653070 130230 653310
rect 130470 653070 130580 653310
rect 130820 653070 130910 653310
rect 131150 653070 131240 653310
rect 131480 653070 131570 653310
rect 131810 653070 131920 653310
rect 132160 653070 132250 653310
rect 132490 653070 132580 653310
rect 132820 653070 132910 653310
rect 133150 653070 133170 653310
rect 122170 652980 133170 653070
rect 122170 652740 122190 652980
rect 122430 652740 122540 652980
rect 122780 652740 122870 652980
rect 123110 652740 123200 652980
rect 123440 652740 123530 652980
rect 123770 652740 123880 652980
rect 124120 652740 124210 652980
rect 124450 652740 124540 652980
rect 124780 652740 124870 652980
rect 125110 652740 125220 652980
rect 125460 652740 125550 652980
rect 125790 652740 125880 652980
rect 126120 652740 126210 652980
rect 126450 652740 126560 652980
rect 126800 652740 126890 652980
rect 127130 652740 127220 652980
rect 127460 652740 127550 652980
rect 127790 652740 127900 652980
rect 128140 652740 128230 652980
rect 128470 652740 128560 652980
rect 128800 652740 128890 652980
rect 129130 652740 129240 652980
rect 129480 652740 129570 652980
rect 129810 652740 129900 652980
rect 130140 652740 130230 652980
rect 130470 652740 130580 652980
rect 130820 652740 130910 652980
rect 131150 652740 131240 652980
rect 131480 652740 131570 652980
rect 131810 652740 131920 652980
rect 132160 652740 132250 652980
rect 132490 652740 132580 652980
rect 132820 652740 132910 652980
rect 133150 652740 133170 652980
rect 122170 652650 133170 652740
rect 122170 652410 122190 652650
rect 122430 652410 122540 652650
rect 122780 652410 122870 652650
rect 123110 652410 123200 652650
rect 123440 652410 123530 652650
rect 123770 652410 123880 652650
rect 124120 652410 124210 652650
rect 124450 652410 124540 652650
rect 124780 652410 124870 652650
rect 125110 652410 125220 652650
rect 125460 652410 125550 652650
rect 125790 652410 125880 652650
rect 126120 652410 126210 652650
rect 126450 652410 126560 652650
rect 126800 652410 126890 652650
rect 127130 652410 127220 652650
rect 127460 652410 127550 652650
rect 127790 652410 127900 652650
rect 128140 652410 128230 652650
rect 128470 652410 128560 652650
rect 128800 652410 128890 652650
rect 129130 652410 129240 652650
rect 129480 652410 129570 652650
rect 129810 652410 129900 652650
rect 130140 652410 130230 652650
rect 130470 652410 130580 652650
rect 130820 652410 130910 652650
rect 131150 652410 131240 652650
rect 131480 652410 131570 652650
rect 131810 652410 131920 652650
rect 132160 652410 132250 652650
rect 132490 652410 132580 652650
rect 132820 652410 132910 652650
rect 133150 652410 133170 652650
rect 122170 652300 133170 652410
rect 122170 652060 122190 652300
rect 122430 652060 122540 652300
rect 122780 652060 122870 652300
rect 123110 652060 123200 652300
rect 123440 652060 123530 652300
rect 123770 652060 123880 652300
rect 124120 652060 124210 652300
rect 124450 652060 124540 652300
rect 124780 652060 124870 652300
rect 125110 652060 125220 652300
rect 125460 652060 125550 652300
rect 125790 652060 125880 652300
rect 126120 652060 126210 652300
rect 126450 652060 126560 652300
rect 126800 652060 126890 652300
rect 127130 652060 127220 652300
rect 127460 652060 127550 652300
rect 127790 652060 127900 652300
rect 128140 652060 128230 652300
rect 128470 652060 128560 652300
rect 128800 652060 128890 652300
rect 129130 652060 129240 652300
rect 129480 652060 129570 652300
rect 129810 652060 129900 652300
rect 130140 652060 130230 652300
rect 130470 652060 130580 652300
rect 130820 652060 130910 652300
rect 131150 652060 131240 652300
rect 131480 652060 131570 652300
rect 131810 652060 131920 652300
rect 132160 652060 132250 652300
rect 132490 652060 132580 652300
rect 132820 652060 132910 652300
rect 133150 652060 133170 652300
rect 122170 651970 133170 652060
rect 122170 651730 122190 651970
rect 122430 651730 122540 651970
rect 122780 651730 122870 651970
rect 123110 651730 123200 651970
rect 123440 651730 123530 651970
rect 123770 651730 123880 651970
rect 124120 651730 124210 651970
rect 124450 651730 124540 651970
rect 124780 651730 124870 651970
rect 125110 651730 125220 651970
rect 125460 651730 125550 651970
rect 125790 651730 125880 651970
rect 126120 651730 126210 651970
rect 126450 651730 126560 651970
rect 126800 651730 126890 651970
rect 127130 651730 127220 651970
rect 127460 651730 127550 651970
rect 127790 651730 127900 651970
rect 128140 651730 128230 651970
rect 128470 651730 128560 651970
rect 128800 651730 128890 651970
rect 129130 651730 129240 651970
rect 129480 651730 129570 651970
rect 129810 651730 129900 651970
rect 130140 651730 130230 651970
rect 130470 651730 130580 651970
rect 130820 651730 130910 651970
rect 131150 651730 131240 651970
rect 131480 651730 131570 651970
rect 131810 651730 131920 651970
rect 132160 651730 132250 651970
rect 132490 651730 132580 651970
rect 132820 651730 132910 651970
rect 133150 651730 133170 651970
rect 122170 651640 133170 651730
rect 122170 651400 122190 651640
rect 122430 651400 122540 651640
rect 122780 651400 122870 651640
rect 123110 651400 123200 651640
rect 123440 651400 123530 651640
rect 123770 651400 123880 651640
rect 124120 651400 124210 651640
rect 124450 651400 124540 651640
rect 124780 651400 124870 651640
rect 125110 651400 125220 651640
rect 125460 651400 125550 651640
rect 125790 651400 125880 651640
rect 126120 651400 126210 651640
rect 126450 651400 126560 651640
rect 126800 651400 126890 651640
rect 127130 651400 127220 651640
rect 127460 651400 127550 651640
rect 127790 651400 127900 651640
rect 128140 651400 128230 651640
rect 128470 651400 128560 651640
rect 128800 651400 128890 651640
rect 129130 651400 129240 651640
rect 129480 651400 129570 651640
rect 129810 651400 129900 651640
rect 130140 651400 130230 651640
rect 130470 651400 130580 651640
rect 130820 651400 130910 651640
rect 131150 651400 131240 651640
rect 131480 651400 131570 651640
rect 131810 651400 131920 651640
rect 132160 651400 132250 651640
rect 132490 651400 132580 651640
rect 132820 651400 132910 651640
rect 133150 651400 133170 651640
rect 122170 651310 133170 651400
rect 122170 651070 122190 651310
rect 122430 651070 122540 651310
rect 122780 651070 122870 651310
rect 123110 651070 123200 651310
rect 123440 651070 123530 651310
rect 123770 651070 123880 651310
rect 124120 651070 124210 651310
rect 124450 651070 124540 651310
rect 124780 651070 124870 651310
rect 125110 651070 125220 651310
rect 125460 651070 125550 651310
rect 125790 651070 125880 651310
rect 126120 651070 126210 651310
rect 126450 651070 126560 651310
rect 126800 651070 126890 651310
rect 127130 651070 127220 651310
rect 127460 651070 127550 651310
rect 127790 651070 127900 651310
rect 128140 651070 128230 651310
rect 128470 651070 128560 651310
rect 128800 651070 128890 651310
rect 129130 651070 129240 651310
rect 129480 651070 129570 651310
rect 129810 651070 129900 651310
rect 130140 651070 130230 651310
rect 130470 651070 130580 651310
rect 130820 651070 130910 651310
rect 131150 651070 131240 651310
rect 131480 651070 131570 651310
rect 131810 651070 131920 651310
rect 132160 651070 132250 651310
rect 132490 651070 132580 651310
rect 132820 651070 132910 651310
rect 133150 651070 133170 651310
rect 122170 650960 133170 651070
rect 122170 650720 122190 650960
rect 122430 650720 122540 650960
rect 122780 650720 122870 650960
rect 123110 650720 123200 650960
rect 123440 650720 123530 650960
rect 123770 650720 123880 650960
rect 124120 650720 124210 650960
rect 124450 650720 124540 650960
rect 124780 650720 124870 650960
rect 125110 650720 125220 650960
rect 125460 650720 125550 650960
rect 125790 650720 125880 650960
rect 126120 650720 126210 650960
rect 126450 650720 126560 650960
rect 126800 650720 126890 650960
rect 127130 650720 127220 650960
rect 127460 650720 127550 650960
rect 127790 650720 127900 650960
rect 128140 650720 128230 650960
rect 128470 650720 128560 650960
rect 128800 650720 128890 650960
rect 129130 650720 129240 650960
rect 129480 650720 129570 650960
rect 129810 650720 129900 650960
rect 130140 650720 130230 650960
rect 130470 650720 130580 650960
rect 130820 650720 130910 650960
rect 131150 650720 131240 650960
rect 131480 650720 131570 650960
rect 131810 650720 131920 650960
rect 132160 650720 132250 650960
rect 132490 650720 132580 650960
rect 132820 650720 132910 650960
rect 133150 650720 133170 650960
rect 122170 650630 133170 650720
rect 122170 650390 122190 650630
rect 122430 650390 122540 650630
rect 122780 650390 122870 650630
rect 123110 650390 123200 650630
rect 123440 650390 123530 650630
rect 123770 650390 123880 650630
rect 124120 650390 124210 650630
rect 124450 650390 124540 650630
rect 124780 650390 124870 650630
rect 125110 650390 125220 650630
rect 125460 650390 125550 650630
rect 125790 650390 125880 650630
rect 126120 650390 126210 650630
rect 126450 650390 126560 650630
rect 126800 650390 126890 650630
rect 127130 650390 127220 650630
rect 127460 650390 127550 650630
rect 127790 650390 127900 650630
rect 128140 650390 128230 650630
rect 128470 650390 128560 650630
rect 128800 650390 128890 650630
rect 129130 650390 129240 650630
rect 129480 650390 129570 650630
rect 129810 650390 129900 650630
rect 130140 650390 130230 650630
rect 130470 650390 130580 650630
rect 130820 650390 130910 650630
rect 131150 650390 131240 650630
rect 131480 650390 131570 650630
rect 131810 650390 131920 650630
rect 132160 650390 132250 650630
rect 132490 650390 132580 650630
rect 132820 650390 132910 650630
rect 133150 650390 133170 650630
rect 122170 650300 133170 650390
rect 122170 650060 122190 650300
rect 122430 650060 122540 650300
rect 122780 650060 122870 650300
rect 123110 650060 123200 650300
rect 123440 650060 123530 650300
rect 123770 650060 123880 650300
rect 124120 650060 124210 650300
rect 124450 650060 124540 650300
rect 124780 650060 124870 650300
rect 125110 650060 125220 650300
rect 125460 650060 125550 650300
rect 125790 650060 125880 650300
rect 126120 650060 126210 650300
rect 126450 650060 126560 650300
rect 126800 650060 126890 650300
rect 127130 650060 127220 650300
rect 127460 650060 127550 650300
rect 127790 650060 127900 650300
rect 128140 650060 128230 650300
rect 128470 650060 128560 650300
rect 128800 650060 128890 650300
rect 129130 650060 129240 650300
rect 129480 650060 129570 650300
rect 129810 650060 129900 650300
rect 130140 650060 130230 650300
rect 130470 650060 130580 650300
rect 130820 650060 130910 650300
rect 131150 650060 131240 650300
rect 131480 650060 131570 650300
rect 131810 650060 131920 650300
rect 132160 650060 132250 650300
rect 132490 650060 132580 650300
rect 132820 650060 132910 650300
rect 133150 650060 133170 650300
rect 122170 649970 133170 650060
rect 122170 649730 122190 649970
rect 122430 649730 122540 649970
rect 122780 649730 122870 649970
rect 123110 649730 123200 649970
rect 123440 649730 123530 649970
rect 123770 649730 123880 649970
rect 124120 649730 124210 649970
rect 124450 649730 124540 649970
rect 124780 649730 124870 649970
rect 125110 649730 125220 649970
rect 125460 649730 125550 649970
rect 125790 649730 125880 649970
rect 126120 649730 126210 649970
rect 126450 649730 126560 649970
rect 126800 649730 126890 649970
rect 127130 649730 127220 649970
rect 127460 649730 127550 649970
rect 127790 649730 127900 649970
rect 128140 649730 128230 649970
rect 128470 649730 128560 649970
rect 128800 649730 128890 649970
rect 129130 649730 129240 649970
rect 129480 649730 129570 649970
rect 129810 649730 129900 649970
rect 130140 649730 130230 649970
rect 130470 649730 130580 649970
rect 130820 649730 130910 649970
rect 131150 649730 131240 649970
rect 131480 649730 131570 649970
rect 131810 649730 131920 649970
rect 132160 649730 132250 649970
rect 132490 649730 132580 649970
rect 132820 649730 132910 649970
rect 133150 649730 133170 649970
rect 122170 649620 133170 649730
rect 122170 649380 122190 649620
rect 122430 649380 122540 649620
rect 122780 649380 122870 649620
rect 123110 649380 123200 649620
rect 123440 649380 123530 649620
rect 123770 649380 123880 649620
rect 124120 649380 124210 649620
rect 124450 649380 124540 649620
rect 124780 649380 124870 649620
rect 125110 649380 125220 649620
rect 125460 649380 125550 649620
rect 125790 649380 125880 649620
rect 126120 649380 126210 649620
rect 126450 649380 126560 649620
rect 126800 649380 126890 649620
rect 127130 649380 127220 649620
rect 127460 649380 127550 649620
rect 127790 649380 127900 649620
rect 128140 649380 128230 649620
rect 128470 649380 128560 649620
rect 128800 649380 128890 649620
rect 129130 649380 129240 649620
rect 129480 649380 129570 649620
rect 129810 649380 129900 649620
rect 130140 649380 130230 649620
rect 130470 649380 130580 649620
rect 130820 649380 130910 649620
rect 131150 649380 131240 649620
rect 131480 649380 131570 649620
rect 131810 649380 131920 649620
rect 132160 649380 132250 649620
rect 132490 649380 132580 649620
rect 132820 649380 132910 649620
rect 133150 649380 133170 649620
rect 122170 649360 133170 649380
rect 133550 660340 144550 660360
rect 133550 660100 133570 660340
rect 133810 660100 133920 660340
rect 134160 660100 134250 660340
rect 134490 660100 134580 660340
rect 134820 660100 134910 660340
rect 135150 660100 135260 660340
rect 135500 660100 135590 660340
rect 135830 660100 135920 660340
rect 136160 660100 136250 660340
rect 136490 660100 136600 660340
rect 136840 660100 136930 660340
rect 137170 660100 137260 660340
rect 137500 660100 137590 660340
rect 137830 660100 137940 660340
rect 138180 660100 138270 660340
rect 138510 660100 138600 660340
rect 138840 660100 138930 660340
rect 139170 660100 139280 660340
rect 139520 660100 139610 660340
rect 139850 660100 139940 660340
rect 140180 660100 140270 660340
rect 140510 660100 140620 660340
rect 140860 660100 140950 660340
rect 141190 660100 141280 660340
rect 141520 660100 141610 660340
rect 141850 660100 141960 660340
rect 142200 660100 142290 660340
rect 142530 660100 142620 660340
rect 142860 660100 142950 660340
rect 143190 660100 143300 660340
rect 143540 660100 143630 660340
rect 143870 660100 143960 660340
rect 144200 660100 144290 660340
rect 144530 660100 144550 660340
rect 133550 660010 144550 660100
rect 133550 659770 133570 660010
rect 133810 659770 133920 660010
rect 134160 659770 134250 660010
rect 134490 659770 134580 660010
rect 134820 659770 134910 660010
rect 135150 659770 135260 660010
rect 135500 659770 135590 660010
rect 135830 659770 135920 660010
rect 136160 659770 136250 660010
rect 136490 659770 136600 660010
rect 136840 659770 136930 660010
rect 137170 659770 137260 660010
rect 137500 659770 137590 660010
rect 137830 659770 137940 660010
rect 138180 659770 138270 660010
rect 138510 659770 138600 660010
rect 138840 659770 138930 660010
rect 139170 659770 139280 660010
rect 139520 659770 139610 660010
rect 139850 659770 139940 660010
rect 140180 659770 140270 660010
rect 140510 659770 140620 660010
rect 140860 659770 140950 660010
rect 141190 659770 141280 660010
rect 141520 659770 141610 660010
rect 141850 659770 141960 660010
rect 142200 659770 142290 660010
rect 142530 659770 142620 660010
rect 142860 659770 142950 660010
rect 143190 659770 143300 660010
rect 143540 659770 143630 660010
rect 143870 659770 143960 660010
rect 144200 659770 144290 660010
rect 144530 659770 144550 660010
rect 133550 659680 144550 659770
rect 133550 659440 133570 659680
rect 133810 659440 133920 659680
rect 134160 659440 134250 659680
rect 134490 659440 134580 659680
rect 134820 659440 134910 659680
rect 135150 659440 135260 659680
rect 135500 659440 135590 659680
rect 135830 659440 135920 659680
rect 136160 659440 136250 659680
rect 136490 659440 136600 659680
rect 136840 659440 136930 659680
rect 137170 659440 137260 659680
rect 137500 659440 137590 659680
rect 137830 659440 137940 659680
rect 138180 659440 138270 659680
rect 138510 659440 138600 659680
rect 138840 659440 138930 659680
rect 139170 659440 139280 659680
rect 139520 659440 139610 659680
rect 139850 659440 139940 659680
rect 140180 659440 140270 659680
rect 140510 659440 140620 659680
rect 140860 659440 140950 659680
rect 141190 659440 141280 659680
rect 141520 659440 141610 659680
rect 141850 659440 141960 659680
rect 142200 659440 142290 659680
rect 142530 659440 142620 659680
rect 142860 659440 142950 659680
rect 143190 659440 143300 659680
rect 143540 659440 143630 659680
rect 143870 659440 143960 659680
rect 144200 659440 144290 659680
rect 144530 659440 144550 659680
rect 133550 659350 144550 659440
rect 133550 659110 133570 659350
rect 133810 659110 133920 659350
rect 134160 659110 134250 659350
rect 134490 659110 134580 659350
rect 134820 659110 134910 659350
rect 135150 659110 135260 659350
rect 135500 659110 135590 659350
rect 135830 659110 135920 659350
rect 136160 659110 136250 659350
rect 136490 659110 136600 659350
rect 136840 659110 136930 659350
rect 137170 659110 137260 659350
rect 137500 659110 137590 659350
rect 137830 659110 137940 659350
rect 138180 659110 138270 659350
rect 138510 659110 138600 659350
rect 138840 659110 138930 659350
rect 139170 659110 139280 659350
rect 139520 659110 139610 659350
rect 139850 659110 139940 659350
rect 140180 659110 140270 659350
rect 140510 659110 140620 659350
rect 140860 659110 140950 659350
rect 141190 659110 141280 659350
rect 141520 659110 141610 659350
rect 141850 659110 141960 659350
rect 142200 659110 142290 659350
rect 142530 659110 142620 659350
rect 142860 659110 142950 659350
rect 143190 659110 143300 659350
rect 143540 659110 143630 659350
rect 143870 659110 143960 659350
rect 144200 659110 144290 659350
rect 144530 659110 144550 659350
rect 133550 659000 144550 659110
rect 133550 658760 133570 659000
rect 133810 658760 133920 659000
rect 134160 658760 134250 659000
rect 134490 658760 134580 659000
rect 134820 658760 134910 659000
rect 135150 658760 135260 659000
rect 135500 658760 135590 659000
rect 135830 658760 135920 659000
rect 136160 658760 136250 659000
rect 136490 658760 136600 659000
rect 136840 658760 136930 659000
rect 137170 658760 137260 659000
rect 137500 658760 137590 659000
rect 137830 658760 137940 659000
rect 138180 658760 138270 659000
rect 138510 658760 138600 659000
rect 138840 658760 138930 659000
rect 139170 658760 139280 659000
rect 139520 658760 139610 659000
rect 139850 658760 139940 659000
rect 140180 658760 140270 659000
rect 140510 658760 140620 659000
rect 140860 658760 140950 659000
rect 141190 658760 141280 659000
rect 141520 658760 141610 659000
rect 141850 658760 141960 659000
rect 142200 658760 142290 659000
rect 142530 658760 142620 659000
rect 142860 658760 142950 659000
rect 143190 658760 143300 659000
rect 143540 658760 143630 659000
rect 143870 658760 143960 659000
rect 144200 658760 144290 659000
rect 144530 658760 144550 659000
rect 133550 658670 144550 658760
rect 133550 658430 133570 658670
rect 133810 658430 133920 658670
rect 134160 658430 134250 658670
rect 134490 658430 134580 658670
rect 134820 658430 134910 658670
rect 135150 658430 135260 658670
rect 135500 658430 135590 658670
rect 135830 658430 135920 658670
rect 136160 658430 136250 658670
rect 136490 658430 136600 658670
rect 136840 658430 136930 658670
rect 137170 658430 137260 658670
rect 137500 658430 137590 658670
rect 137830 658430 137940 658670
rect 138180 658430 138270 658670
rect 138510 658430 138600 658670
rect 138840 658430 138930 658670
rect 139170 658430 139280 658670
rect 139520 658430 139610 658670
rect 139850 658430 139940 658670
rect 140180 658430 140270 658670
rect 140510 658430 140620 658670
rect 140860 658430 140950 658670
rect 141190 658430 141280 658670
rect 141520 658430 141610 658670
rect 141850 658430 141960 658670
rect 142200 658430 142290 658670
rect 142530 658430 142620 658670
rect 142860 658430 142950 658670
rect 143190 658430 143300 658670
rect 143540 658430 143630 658670
rect 143870 658430 143960 658670
rect 144200 658430 144290 658670
rect 144530 658430 144550 658670
rect 133550 658340 144550 658430
rect 133550 658100 133570 658340
rect 133810 658100 133920 658340
rect 134160 658100 134250 658340
rect 134490 658100 134580 658340
rect 134820 658100 134910 658340
rect 135150 658100 135260 658340
rect 135500 658100 135590 658340
rect 135830 658100 135920 658340
rect 136160 658100 136250 658340
rect 136490 658100 136600 658340
rect 136840 658100 136930 658340
rect 137170 658100 137260 658340
rect 137500 658100 137590 658340
rect 137830 658100 137940 658340
rect 138180 658100 138270 658340
rect 138510 658100 138600 658340
rect 138840 658100 138930 658340
rect 139170 658100 139280 658340
rect 139520 658100 139610 658340
rect 139850 658100 139940 658340
rect 140180 658100 140270 658340
rect 140510 658100 140620 658340
rect 140860 658100 140950 658340
rect 141190 658100 141280 658340
rect 141520 658100 141610 658340
rect 141850 658100 141960 658340
rect 142200 658100 142290 658340
rect 142530 658100 142620 658340
rect 142860 658100 142950 658340
rect 143190 658100 143300 658340
rect 143540 658100 143630 658340
rect 143870 658100 143960 658340
rect 144200 658100 144290 658340
rect 144530 658100 144550 658340
rect 133550 658010 144550 658100
rect 133550 657770 133570 658010
rect 133810 657770 133920 658010
rect 134160 657770 134250 658010
rect 134490 657770 134580 658010
rect 134820 657770 134910 658010
rect 135150 657770 135260 658010
rect 135500 657770 135590 658010
rect 135830 657770 135920 658010
rect 136160 657770 136250 658010
rect 136490 657770 136600 658010
rect 136840 657770 136930 658010
rect 137170 657770 137260 658010
rect 137500 657770 137590 658010
rect 137830 657770 137940 658010
rect 138180 657770 138270 658010
rect 138510 657770 138600 658010
rect 138840 657770 138930 658010
rect 139170 657770 139280 658010
rect 139520 657770 139610 658010
rect 139850 657770 139940 658010
rect 140180 657770 140270 658010
rect 140510 657770 140620 658010
rect 140860 657770 140950 658010
rect 141190 657770 141280 658010
rect 141520 657770 141610 658010
rect 141850 657770 141960 658010
rect 142200 657770 142290 658010
rect 142530 657770 142620 658010
rect 142860 657770 142950 658010
rect 143190 657770 143300 658010
rect 143540 657770 143630 658010
rect 143870 657770 143960 658010
rect 144200 657770 144290 658010
rect 144530 657770 144550 658010
rect 133550 657660 144550 657770
rect 133550 657420 133570 657660
rect 133810 657420 133920 657660
rect 134160 657420 134250 657660
rect 134490 657420 134580 657660
rect 134820 657420 134910 657660
rect 135150 657420 135260 657660
rect 135500 657420 135590 657660
rect 135830 657420 135920 657660
rect 136160 657420 136250 657660
rect 136490 657420 136600 657660
rect 136840 657420 136930 657660
rect 137170 657420 137260 657660
rect 137500 657420 137590 657660
rect 137830 657420 137940 657660
rect 138180 657420 138270 657660
rect 138510 657420 138600 657660
rect 138840 657420 138930 657660
rect 139170 657420 139280 657660
rect 139520 657420 139610 657660
rect 139850 657420 139940 657660
rect 140180 657420 140270 657660
rect 140510 657420 140620 657660
rect 140860 657420 140950 657660
rect 141190 657420 141280 657660
rect 141520 657420 141610 657660
rect 141850 657420 141960 657660
rect 142200 657420 142290 657660
rect 142530 657420 142620 657660
rect 142860 657420 142950 657660
rect 143190 657420 143300 657660
rect 143540 657420 143630 657660
rect 143870 657420 143960 657660
rect 144200 657420 144290 657660
rect 144530 657420 144550 657660
rect 133550 657330 144550 657420
rect 133550 657090 133570 657330
rect 133810 657090 133920 657330
rect 134160 657090 134250 657330
rect 134490 657090 134580 657330
rect 134820 657090 134910 657330
rect 135150 657090 135260 657330
rect 135500 657090 135590 657330
rect 135830 657090 135920 657330
rect 136160 657090 136250 657330
rect 136490 657090 136600 657330
rect 136840 657090 136930 657330
rect 137170 657090 137260 657330
rect 137500 657090 137590 657330
rect 137830 657090 137940 657330
rect 138180 657090 138270 657330
rect 138510 657090 138600 657330
rect 138840 657090 138930 657330
rect 139170 657090 139280 657330
rect 139520 657090 139610 657330
rect 139850 657090 139940 657330
rect 140180 657090 140270 657330
rect 140510 657090 140620 657330
rect 140860 657090 140950 657330
rect 141190 657090 141280 657330
rect 141520 657090 141610 657330
rect 141850 657090 141960 657330
rect 142200 657090 142290 657330
rect 142530 657090 142620 657330
rect 142860 657090 142950 657330
rect 143190 657090 143300 657330
rect 143540 657090 143630 657330
rect 143870 657090 143960 657330
rect 144200 657090 144290 657330
rect 144530 657090 144550 657330
rect 133550 657000 144550 657090
rect 133550 656760 133570 657000
rect 133810 656760 133920 657000
rect 134160 656760 134250 657000
rect 134490 656760 134580 657000
rect 134820 656760 134910 657000
rect 135150 656760 135260 657000
rect 135500 656760 135590 657000
rect 135830 656760 135920 657000
rect 136160 656760 136250 657000
rect 136490 656760 136600 657000
rect 136840 656760 136930 657000
rect 137170 656760 137260 657000
rect 137500 656760 137590 657000
rect 137830 656760 137940 657000
rect 138180 656760 138270 657000
rect 138510 656760 138600 657000
rect 138840 656760 138930 657000
rect 139170 656760 139280 657000
rect 139520 656760 139610 657000
rect 139850 656760 139940 657000
rect 140180 656760 140270 657000
rect 140510 656760 140620 657000
rect 140860 656760 140950 657000
rect 141190 656760 141280 657000
rect 141520 656760 141610 657000
rect 141850 656760 141960 657000
rect 142200 656760 142290 657000
rect 142530 656760 142620 657000
rect 142860 656760 142950 657000
rect 143190 656760 143300 657000
rect 143540 656760 143630 657000
rect 143870 656760 143960 657000
rect 144200 656760 144290 657000
rect 144530 656760 144550 657000
rect 133550 656670 144550 656760
rect 133550 656430 133570 656670
rect 133810 656430 133920 656670
rect 134160 656430 134250 656670
rect 134490 656430 134580 656670
rect 134820 656430 134910 656670
rect 135150 656430 135260 656670
rect 135500 656430 135590 656670
rect 135830 656430 135920 656670
rect 136160 656430 136250 656670
rect 136490 656430 136600 656670
rect 136840 656430 136930 656670
rect 137170 656430 137260 656670
rect 137500 656430 137590 656670
rect 137830 656430 137940 656670
rect 138180 656430 138270 656670
rect 138510 656430 138600 656670
rect 138840 656430 138930 656670
rect 139170 656430 139280 656670
rect 139520 656430 139610 656670
rect 139850 656430 139940 656670
rect 140180 656430 140270 656670
rect 140510 656430 140620 656670
rect 140860 656430 140950 656670
rect 141190 656430 141280 656670
rect 141520 656430 141610 656670
rect 141850 656430 141960 656670
rect 142200 656430 142290 656670
rect 142530 656430 142620 656670
rect 142860 656430 142950 656670
rect 143190 656430 143300 656670
rect 143540 656430 143630 656670
rect 143870 656430 143960 656670
rect 144200 656430 144290 656670
rect 144530 656430 144550 656670
rect 133550 656320 144550 656430
rect 133550 656080 133570 656320
rect 133810 656080 133920 656320
rect 134160 656080 134250 656320
rect 134490 656080 134580 656320
rect 134820 656080 134910 656320
rect 135150 656080 135260 656320
rect 135500 656080 135590 656320
rect 135830 656080 135920 656320
rect 136160 656080 136250 656320
rect 136490 656080 136600 656320
rect 136840 656080 136930 656320
rect 137170 656080 137260 656320
rect 137500 656080 137590 656320
rect 137830 656080 137940 656320
rect 138180 656080 138270 656320
rect 138510 656080 138600 656320
rect 138840 656080 138930 656320
rect 139170 656080 139280 656320
rect 139520 656080 139610 656320
rect 139850 656080 139940 656320
rect 140180 656080 140270 656320
rect 140510 656080 140620 656320
rect 140860 656080 140950 656320
rect 141190 656080 141280 656320
rect 141520 656080 141610 656320
rect 141850 656080 141960 656320
rect 142200 656080 142290 656320
rect 142530 656080 142620 656320
rect 142860 656080 142950 656320
rect 143190 656080 143300 656320
rect 143540 656080 143630 656320
rect 143870 656080 143960 656320
rect 144200 656080 144290 656320
rect 144530 656080 144550 656320
rect 133550 655990 144550 656080
rect 133550 655750 133570 655990
rect 133810 655750 133920 655990
rect 134160 655750 134250 655990
rect 134490 655750 134580 655990
rect 134820 655750 134910 655990
rect 135150 655750 135260 655990
rect 135500 655750 135590 655990
rect 135830 655750 135920 655990
rect 136160 655750 136250 655990
rect 136490 655750 136600 655990
rect 136840 655750 136930 655990
rect 137170 655750 137260 655990
rect 137500 655750 137590 655990
rect 137830 655750 137940 655990
rect 138180 655750 138270 655990
rect 138510 655750 138600 655990
rect 138840 655750 138930 655990
rect 139170 655750 139280 655990
rect 139520 655750 139610 655990
rect 139850 655750 139940 655990
rect 140180 655750 140270 655990
rect 140510 655750 140620 655990
rect 140860 655750 140950 655990
rect 141190 655750 141280 655990
rect 141520 655750 141610 655990
rect 141850 655750 141960 655990
rect 142200 655750 142290 655990
rect 142530 655750 142620 655990
rect 142860 655750 142950 655990
rect 143190 655750 143300 655990
rect 143540 655750 143630 655990
rect 143870 655750 143960 655990
rect 144200 655750 144290 655990
rect 144530 655750 144550 655990
rect 133550 655660 144550 655750
rect 133550 655420 133570 655660
rect 133810 655420 133920 655660
rect 134160 655420 134250 655660
rect 134490 655420 134580 655660
rect 134820 655420 134910 655660
rect 135150 655420 135260 655660
rect 135500 655420 135590 655660
rect 135830 655420 135920 655660
rect 136160 655420 136250 655660
rect 136490 655420 136600 655660
rect 136840 655420 136930 655660
rect 137170 655420 137260 655660
rect 137500 655420 137590 655660
rect 137830 655420 137940 655660
rect 138180 655420 138270 655660
rect 138510 655420 138600 655660
rect 138840 655420 138930 655660
rect 139170 655420 139280 655660
rect 139520 655420 139610 655660
rect 139850 655420 139940 655660
rect 140180 655420 140270 655660
rect 140510 655420 140620 655660
rect 140860 655420 140950 655660
rect 141190 655420 141280 655660
rect 141520 655420 141610 655660
rect 141850 655420 141960 655660
rect 142200 655420 142290 655660
rect 142530 655420 142620 655660
rect 142860 655420 142950 655660
rect 143190 655420 143300 655660
rect 143540 655420 143630 655660
rect 143870 655420 143960 655660
rect 144200 655420 144290 655660
rect 144530 655420 144550 655660
rect 133550 655330 144550 655420
rect 133550 655090 133570 655330
rect 133810 655090 133920 655330
rect 134160 655090 134250 655330
rect 134490 655090 134580 655330
rect 134820 655090 134910 655330
rect 135150 655090 135260 655330
rect 135500 655090 135590 655330
rect 135830 655090 135920 655330
rect 136160 655090 136250 655330
rect 136490 655090 136600 655330
rect 136840 655090 136930 655330
rect 137170 655090 137260 655330
rect 137500 655090 137590 655330
rect 137830 655090 137940 655330
rect 138180 655090 138270 655330
rect 138510 655090 138600 655330
rect 138840 655090 138930 655330
rect 139170 655090 139280 655330
rect 139520 655090 139610 655330
rect 139850 655090 139940 655330
rect 140180 655090 140270 655330
rect 140510 655090 140620 655330
rect 140860 655090 140950 655330
rect 141190 655090 141280 655330
rect 141520 655090 141610 655330
rect 141850 655090 141960 655330
rect 142200 655090 142290 655330
rect 142530 655090 142620 655330
rect 142860 655090 142950 655330
rect 143190 655090 143300 655330
rect 143540 655090 143630 655330
rect 143870 655090 143960 655330
rect 144200 655090 144290 655330
rect 144530 655090 144550 655330
rect 133550 654980 144550 655090
rect 133550 654740 133570 654980
rect 133810 654740 133920 654980
rect 134160 654740 134250 654980
rect 134490 654740 134580 654980
rect 134820 654740 134910 654980
rect 135150 654740 135260 654980
rect 135500 654740 135590 654980
rect 135830 654740 135920 654980
rect 136160 654740 136250 654980
rect 136490 654740 136600 654980
rect 136840 654740 136930 654980
rect 137170 654740 137260 654980
rect 137500 654740 137590 654980
rect 137830 654740 137940 654980
rect 138180 654740 138270 654980
rect 138510 654740 138600 654980
rect 138840 654740 138930 654980
rect 139170 654740 139280 654980
rect 139520 654740 139610 654980
rect 139850 654740 139940 654980
rect 140180 654740 140270 654980
rect 140510 654740 140620 654980
rect 140860 654740 140950 654980
rect 141190 654740 141280 654980
rect 141520 654740 141610 654980
rect 141850 654740 141960 654980
rect 142200 654740 142290 654980
rect 142530 654740 142620 654980
rect 142860 654740 142950 654980
rect 143190 654740 143300 654980
rect 143540 654740 143630 654980
rect 143870 654740 143960 654980
rect 144200 654740 144290 654980
rect 144530 654740 144550 654980
rect 133550 654650 144550 654740
rect 133550 654410 133570 654650
rect 133810 654410 133920 654650
rect 134160 654410 134250 654650
rect 134490 654410 134580 654650
rect 134820 654410 134910 654650
rect 135150 654410 135260 654650
rect 135500 654410 135590 654650
rect 135830 654410 135920 654650
rect 136160 654410 136250 654650
rect 136490 654410 136600 654650
rect 136840 654410 136930 654650
rect 137170 654410 137260 654650
rect 137500 654410 137590 654650
rect 137830 654410 137940 654650
rect 138180 654410 138270 654650
rect 138510 654410 138600 654650
rect 138840 654410 138930 654650
rect 139170 654410 139280 654650
rect 139520 654410 139610 654650
rect 139850 654410 139940 654650
rect 140180 654410 140270 654650
rect 140510 654410 140620 654650
rect 140860 654410 140950 654650
rect 141190 654410 141280 654650
rect 141520 654410 141610 654650
rect 141850 654410 141960 654650
rect 142200 654410 142290 654650
rect 142530 654410 142620 654650
rect 142860 654410 142950 654650
rect 143190 654410 143300 654650
rect 143540 654410 143630 654650
rect 143870 654410 143960 654650
rect 144200 654410 144290 654650
rect 144530 654410 144550 654650
rect 133550 654320 144550 654410
rect 133550 654080 133570 654320
rect 133810 654080 133920 654320
rect 134160 654080 134250 654320
rect 134490 654080 134580 654320
rect 134820 654080 134910 654320
rect 135150 654080 135260 654320
rect 135500 654080 135590 654320
rect 135830 654080 135920 654320
rect 136160 654080 136250 654320
rect 136490 654080 136600 654320
rect 136840 654080 136930 654320
rect 137170 654080 137260 654320
rect 137500 654080 137590 654320
rect 137830 654080 137940 654320
rect 138180 654080 138270 654320
rect 138510 654080 138600 654320
rect 138840 654080 138930 654320
rect 139170 654080 139280 654320
rect 139520 654080 139610 654320
rect 139850 654080 139940 654320
rect 140180 654080 140270 654320
rect 140510 654080 140620 654320
rect 140860 654080 140950 654320
rect 141190 654080 141280 654320
rect 141520 654080 141610 654320
rect 141850 654080 141960 654320
rect 142200 654080 142290 654320
rect 142530 654080 142620 654320
rect 142860 654080 142950 654320
rect 143190 654080 143300 654320
rect 143540 654080 143630 654320
rect 143870 654080 143960 654320
rect 144200 654080 144290 654320
rect 144530 654080 144550 654320
rect 133550 653990 144550 654080
rect 133550 653750 133570 653990
rect 133810 653750 133920 653990
rect 134160 653750 134250 653990
rect 134490 653750 134580 653990
rect 134820 653750 134910 653990
rect 135150 653750 135260 653990
rect 135500 653750 135590 653990
rect 135830 653750 135920 653990
rect 136160 653750 136250 653990
rect 136490 653750 136600 653990
rect 136840 653750 136930 653990
rect 137170 653750 137260 653990
rect 137500 653750 137590 653990
rect 137830 653750 137940 653990
rect 138180 653750 138270 653990
rect 138510 653750 138600 653990
rect 138840 653750 138930 653990
rect 139170 653750 139280 653990
rect 139520 653750 139610 653990
rect 139850 653750 139940 653990
rect 140180 653750 140270 653990
rect 140510 653750 140620 653990
rect 140860 653750 140950 653990
rect 141190 653750 141280 653990
rect 141520 653750 141610 653990
rect 141850 653750 141960 653990
rect 142200 653750 142290 653990
rect 142530 653750 142620 653990
rect 142860 653750 142950 653990
rect 143190 653750 143300 653990
rect 143540 653750 143630 653990
rect 143870 653750 143960 653990
rect 144200 653750 144290 653990
rect 144530 653750 144550 653990
rect 133550 653640 144550 653750
rect 133550 653400 133570 653640
rect 133810 653400 133920 653640
rect 134160 653400 134250 653640
rect 134490 653400 134580 653640
rect 134820 653400 134910 653640
rect 135150 653400 135260 653640
rect 135500 653400 135590 653640
rect 135830 653400 135920 653640
rect 136160 653400 136250 653640
rect 136490 653400 136600 653640
rect 136840 653400 136930 653640
rect 137170 653400 137260 653640
rect 137500 653400 137590 653640
rect 137830 653400 137940 653640
rect 138180 653400 138270 653640
rect 138510 653400 138600 653640
rect 138840 653400 138930 653640
rect 139170 653400 139280 653640
rect 139520 653400 139610 653640
rect 139850 653400 139940 653640
rect 140180 653400 140270 653640
rect 140510 653400 140620 653640
rect 140860 653400 140950 653640
rect 141190 653400 141280 653640
rect 141520 653400 141610 653640
rect 141850 653400 141960 653640
rect 142200 653400 142290 653640
rect 142530 653400 142620 653640
rect 142860 653400 142950 653640
rect 143190 653400 143300 653640
rect 143540 653400 143630 653640
rect 143870 653400 143960 653640
rect 144200 653400 144290 653640
rect 144530 653400 144550 653640
rect 133550 653310 144550 653400
rect 133550 653070 133570 653310
rect 133810 653070 133920 653310
rect 134160 653070 134250 653310
rect 134490 653070 134580 653310
rect 134820 653070 134910 653310
rect 135150 653070 135260 653310
rect 135500 653070 135590 653310
rect 135830 653070 135920 653310
rect 136160 653070 136250 653310
rect 136490 653070 136600 653310
rect 136840 653070 136930 653310
rect 137170 653070 137260 653310
rect 137500 653070 137590 653310
rect 137830 653070 137940 653310
rect 138180 653070 138270 653310
rect 138510 653070 138600 653310
rect 138840 653070 138930 653310
rect 139170 653070 139280 653310
rect 139520 653070 139610 653310
rect 139850 653070 139940 653310
rect 140180 653070 140270 653310
rect 140510 653070 140620 653310
rect 140860 653070 140950 653310
rect 141190 653070 141280 653310
rect 141520 653070 141610 653310
rect 141850 653070 141960 653310
rect 142200 653070 142290 653310
rect 142530 653070 142620 653310
rect 142860 653070 142950 653310
rect 143190 653070 143300 653310
rect 143540 653070 143630 653310
rect 143870 653070 143960 653310
rect 144200 653070 144290 653310
rect 144530 653070 144550 653310
rect 133550 652980 144550 653070
rect 133550 652740 133570 652980
rect 133810 652740 133920 652980
rect 134160 652740 134250 652980
rect 134490 652740 134580 652980
rect 134820 652740 134910 652980
rect 135150 652740 135260 652980
rect 135500 652740 135590 652980
rect 135830 652740 135920 652980
rect 136160 652740 136250 652980
rect 136490 652740 136600 652980
rect 136840 652740 136930 652980
rect 137170 652740 137260 652980
rect 137500 652740 137590 652980
rect 137830 652740 137940 652980
rect 138180 652740 138270 652980
rect 138510 652740 138600 652980
rect 138840 652740 138930 652980
rect 139170 652740 139280 652980
rect 139520 652740 139610 652980
rect 139850 652740 139940 652980
rect 140180 652740 140270 652980
rect 140510 652740 140620 652980
rect 140860 652740 140950 652980
rect 141190 652740 141280 652980
rect 141520 652740 141610 652980
rect 141850 652740 141960 652980
rect 142200 652740 142290 652980
rect 142530 652740 142620 652980
rect 142860 652740 142950 652980
rect 143190 652740 143300 652980
rect 143540 652740 143630 652980
rect 143870 652740 143960 652980
rect 144200 652740 144290 652980
rect 144530 652740 144550 652980
rect 133550 652650 144550 652740
rect 133550 652410 133570 652650
rect 133810 652410 133920 652650
rect 134160 652410 134250 652650
rect 134490 652410 134580 652650
rect 134820 652410 134910 652650
rect 135150 652410 135260 652650
rect 135500 652410 135590 652650
rect 135830 652410 135920 652650
rect 136160 652410 136250 652650
rect 136490 652410 136600 652650
rect 136840 652410 136930 652650
rect 137170 652410 137260 652650
rect 137500 652410 137590 652650
rect 137830 652410 137940 652650
rect 138180 652410 138270 652650
rect 138510 652410 138600 652650
rect 138840 652410 138930 652650
rect 139170 652410 139280 652650
rect 139520 652410 139610 652650
rect 139850 652410 139940 652650
rect 140180 652410 140270 652650
rect 140510 652410 140620 652650
rect 140860 652410 140950 652650
rect 141190 652410 141280 652650
rect 141520 652410 141610 652650
rect 141850 652410 141960 652650
rect 142200 652410 142290 652650
rect 142530 652410 142620 652650
rect 142860 652410 142950 652650
rect 143190 652410 143300 652650
rect 143540 652410 143630 652650
rect 143870 652410 143960 652650
rect 144200 652410 144290 652650
rect 144530 652410 144550 652650
rect 133550 652300 144550 652410
rect 133550 652060 133570 652300
rect 133810 652060 133920 652300
rect 134160 652060 134250 652300
rect 134490 652060 134580 652300
rect 134820 652060 134910 652300
rect 135150 652060 135260 652300
rect 135500 652060 135590 652300
rect 135830 652060 135920 652300
rect 136160 652060 136250 652300
rect 136490 652060 136600 652300
rect 136840 652060 136930 652300
rect 137170 652060 137260 652300
rect 137500 652060 137590 652300
rect 137830 652060 137940 652300
rect 138180 652060 138270 652300
rect 138510 652060 138600 652300
rect 138840 652060 138930 652300
rect 139170 652060 139280 652300
rect 139520 652060 139610 652300
rect 139850 652060 139940 652300
rect 140180 652060 140270 652300
rect 140510 652060 140620 652300
rect 140860 652060 140950 652300
rect 141190 652060 141280 652300
rect 141520 652060 141610 652300
rect 141850 652060 141960 652300
rect 142200 652060 142290 652300
rect 142530 652060 142620 652300
rect 142860 652060 142950 652300
rect 143190 652060 143300 652300
rect 143540 652060 143630 652300
rect 143870 652060 143960 652300
rect 144200 652060 144290 652300
rect 144530 652060 144550 652300
rect 133550 651970 144550 652060
rect 133550 651730 133570 651970
rect 133810 651730 133920 651970
rect 134160 651730 134250 651970
rect 134490 651730 134580 651970
rect 134820 651730 134910 651970
rect 135150 651730 135260 651970
rect 135500 651730 135590 651970
rect 135830 651730 135920 651970
rect 136160 651730 136250 651970
rect 136490 651730 136600 651970
rect 136840 651730 136930 651970
rect 137170 651730 137260 651970
rect 137500 651730 137590 651970
rect 137830 651730 137940 651970
rect 138180 651730 138270 651970
rect 138510 651730 138600 651970
rect 138840 651730 138930 651970
rect 139170 651730 139280 651970
rect 139520 651730 139610 651970
rect 139850 651730 139940 651970
rect 140180 651730 140270 651970
rect 140510 651730 140620 651970
rect 140860 651730 140950 651970
rect 141190 651730 141280 651970
rect 141520 651730 141610 651970
rect 141850 651730 141960 651970
rect 142200 651730 142290 651970
rect 142530 651730 142620 651970
rect 142860 651730 142950 651970
rect 143190 651730 143300 651970
rect 143540 651730 143630 651970
rect 143870 651730 143960 651970
rect 144200 651730 144290 651970
rect 144530 651730 144550 651970
rect 133550 651640 144550 651730
rect 133550 651400 133570 651640
rect 133810 651400 133920 651640
rect 134160 651400 134250 651640
rect 134490 651400 134580 651640
rect 134820 651400 134910 651640
rect 135150 651400 135260 651640
rect 135500 651400 135590 651640
rect 135830 651400 135920 651640
rect 136160 651400 136250 651640
rect 136490 651400 136600 651640
rect 136840 651400 136930 651640
rect 137170 651400 137260 651640
rect 137500 651400 137590 651640
rect 137830 651400 137940 651640
rect 138180 651400 138270 651640
rect 138510 651400 138600 651640
rect 138840 651400 138930 651640
rect 139170 651400 139280 651640
rect 139520 651400 139610 651640
rect 139850 651400 139940 651640
rect 140180 651400 140270 651640
rect 140510 651400 140620 651640
rect 140860 651400 140950 651640
rect 141190 651400 141280 651640
rect 141520 651400 141610 651640
rect 141850 651400 141960 651640
rect 142200 651400 142290 651640
rect 142530 651400 142620 651640
rect 142860 651400 142950 651640
rect 143190 651400 143300 651640
rect 143540 651400 143630 651640
rect 143870 651400 143960 651640
rect 144200 651400 144290 651640
rect 144530 651400 144550 651640
rect 133550 651310 144550 651400
rect 133550 651070 133570 651310
rect 133810 651070 133920 651310
rect 134160 651070 134250 651310
rect 134490 651070 134580 651310
rect 134820 651070 134910 651310
rect 135150 651070 135260 651310
rect 135500 651070 135590 651310
rect 135830 651070 135920 651310
rect 136160 651070 136250 651310
rect 136490 651070 136600 651310
rect 136840 651070 136930 651310
rect 137170 651070 137260 651310
rect 137500 651070 137590 651310
rect 137830 651070 137940 651310
rect 138180 651070 138270 651310
rect 138510 651070 138600 651310
rect 138840 651070 138930 651310
rect 139170 651070 139280 651310
rect 139520 651070 139610 651310
rect 139850 651070 139940 651310
rect 140180 651070 140270 651310
rect 140510 651070 140620 651310
rect 140860 651070 140950 651310
rect 141190 651070 141280 651310
rect 141520 651070 141610 651310
rect 141850 651070 141960 651310
rect 142200 651070 142290 651310
rect 142530 651070 142620 651310
rect 142860 651070 142950 651310
rect 143190 651070 143300 651310
rect 143540 651070 143630 651310
rect 143870 651070 143960 651310
rect 144200 651070 144290 651310
rect 144530 651070 144550 651310
rect 133550 650960 144550 651070
rect 133550 650720 133570 650960
rect 133810 650720 133920 650960
rect 134160 650720 134250 650960
rect 134490 650720 134580 650960
rect 134820 650720 134910 650960
rect 135150 650720 135260 650960
rect 135500 650720 135590 650960
rect 135830 650720 135920 650960
rect 136160 650720 136250 650960
rect 136490 650720 136600 650960
rect 136840 650720 136930 650960
rect 137170 650720 137260 650960
rect 137500 650720 137590 650960
rect 137830 650720 137940 650960
rect 138180 650720 138270 650960
rect 138510 650720 138600 650960
rect 138840 650720 138930 650960
rect 139170 650720 139280 650960
rect 139520 650720 139610 650960
rect 139850 650720 139940 650960
rect 140180 650720 140270 650960
rect 140510 650720 140620 650960
rect 140860 650720 140950 650960
rect 141190 650720 141280 650960
rect 141520 650720 141610 650960
rect 141850 650720 141960 650960
rect 142200 650720 142290 650960
rect 142530 650720 142620 650960
rect 142860 650720 142950 650960
rect 143190 650720 143300 650960
rect 143540 650720 143630 650960
rect 143870 650720 143960 650960
rect 144200 650720 144290 650960
rect 144530 650720 144550 650960
rect 133550 650630 144550 650720
rect 133550 650390 133570 650630
rect 133810 650390 133920 650630
rect 134160 650390 134250 650630
rect 134490 650390 134580 650630
rect 134820 650390 134910 650630
rect 135150 650390 135260 650630
rect 135500 650390 135590 650630
rect 135830 650390 135920 650630
rect 136160 650390 136250 650630
rect 136490 650390 136600 650630
rect 136840 650390 136930 650630
rect 137170 650390 137260 650630
rect 137500 650390 137590 650630
rect 137830 650390 137940 650630
rect 138180 650390 138270 650630
rect 138510 650390 138600 650630
rect 138840 650390 138930 650630
rect 139170 650390 139280 650630
rect 139520 650390 139610 650630
rect 139850 650390 139940 650630
rect 140180 650390 140270 650630
rect 140510 650390 140620 650630
rect 140860 650390 140950 650630
rect 141190 650390 141280 650630
rect 141520 650390 141610 650630
rect 141850 650390 141960 650630
rect 142200 650390 142290 650630
rect 142530 650390 142620 650630
rect 142860 650390 142950 650630
rect 143190 650390 143300 650630
rect 143540 650390 143630 650630
rect 143870 650390 143960 650630
rect 144200 650390 144290 650630
rect 144530 650390 144550 650630
rect 133550 650300 144550 650390
rect 133550 650060 133570 650300
rect 133810 650060 133920 650300
rect 134160 650060 134250 650300
rect 134490 650060 134580 650300
rect 134820 650060 134910 650300
rect 135150 650060 135260 650300
rect 135500 650060 135590 650300
rect 135830 650060 135920 650300
rect 136160 650060 136250 650300
rect 136490 650060 136600 650300
rect 136840 650060 136930 650300
rect 137170 650060 137260 650300
rect 137500 650060 137590 650300
rect 137830 650060 137940 650300
rect 138180 650060 138270 650300
rect 138510 650060 138600 650300
rect 138840 650060 138930 650300
rect 139170 650060 139280 650300
rect 139520 650060 139610 650300
rect 139850 650060 139940 650300
rect 140180 650060 140270 650300
rect 140510 650060 140620 650300
rect 140860 650060 140950 650300
rect 141190 650060 141280 650300
rect 141520 650060 141610 650300
rect 141850 650060 141960 650300
rect 142200 650060 142290 650300
rect 142530 650060 142620 650300
rect 142860 650060 142950 650300
rect 143190 650060 143300 650300
rect 143540 650060 143630 650300
rect 143870 650060 143960 650300
rect 144200 650060 144290 650300
rect 144530 650060 144550 650300
rect 133550 649970 144550 650060
rect 133550 649730 133570 649970
rect 133810 649730 133920 649970
rect 134160 649730 134250 649970
rect 134490 649730 134580 649970
rect 134820 649730 134910 649970
rect 135150 649730 135260 649970
rect 135500 649730 135590 649970
rect 135830 649730 135920 649970
rect 136160 649730 136250 649970
rect 136490 649730 136600 649970
rect 136840 649730 136930 649970
rect 137170 649730 137260 649970
rect 137500 649730 137590 649970
rect 137830 649730 137940 649970
rect 138180 649730 138270 649970
rect 138510 649730 138600 649970
rect 138840 649730 138930 649970
rect 139170 649730 139280 649970
rect 139520 649730 139610 649970
rect 139850 649730 139940 649970
rect 140180 649730 140270 649970
rect 140510 649730 140620 649970
rect 140860 649730 140950 649970
rect 141190 649730 141280 649970
rect 141520 649730 141610 649970
rect 141850 649730 141960 649970
rect 142200 649730 142290 649970
rect 142530 649730 142620 649970
rect 142860 649730 142950 649970
rect 143190 649730 143300 649970
rect 143540 649730 143630 649970
rect 143870 649730 143960 649970
rect 144200 649730 144290 649970
rect 144530 649730 144550 649970
rect 133550 649620 144550 649730
rect 133550 649380 133570 649620
rect 133810 649380 133920 649620
rect 134160 649380 134250 649620
rect 134490 649380 134580 649620
rect 134820 649380 134910 649620
rect 135150 649380 135260 649620
rect 135500 649380 135590 649620
rect 135830 649380 135920 649620
rect 136160 649380 136250 649620
rect 136490 649380 136600 649620
rect 136840 649380 136930 649620
rect 137170 649380 137260 649620
rect 137500 649380 137590 649620
rect 137830 649380 137940 649620
rect 138180 649380 138270 649620
rect 138510 649380 138600 649620
rect 138840 649380 138930 649620
rect 139170 649380 139280 649620
rect 139520 649380 139610 649620
rect 139850 649380 139940 649620
rect 140180 649380 140270 649620
rect 140510 649380 140620 649620
rect 140860 649380 140950 649620
rect 141190 649380 141280 649620
rect 141520 649380 141610 649620
rect 141850 649380 141960 649620
rect 142200 649380 142290 649620
rect 142530 649380 142620 649620
rect 142860 649380 142950 649620
rect 143190 649380 143300 649620
rect 143540 649380 143630 649620
rect 143870 649380 143960 649620
rect 144200 649380 144290 649620
rect 144530 649380 144550 649620
rect 133550 649360 144550 649380
rect 144930 660340 155930 660360
rect 144930 660100 144950 660340
rect 145190 660100 145300 660340
rect 145540 660100 145630 660340
rect 145870 660100 145960 660340
rect 146200 660100 146290 660340
rect 146530 660100 146640 660340
rect 146880 660100 146970 660340
rect 147210 660100 147300 660340
rect 147540 660100 147630 660340
rect 147870 660100 147980 660340
rect 148220 660100 148310 660340
rect 148550 660100 148640 660340
rect 148880 660100 148970 660340
rect 149210 660100 149320 660340
rect 149560 660100 149650 660340
rect 149890 660100 149980 660340
rect 150220 660100 150310 660340
rect 150550 660100 150660 660340
rect 150900 660100 150990 660340
rect 151230 660100 151320 660340
rect 151560 660100 151650 660340
rect 151890 660100 152000 660340
rect 152240 660100 152330 660340
rect 152570 660100 152660 660340
rect 152900 660100 152990 660340
rect 153230 660100 153340 660340
rect 153580 660100 153670 660340
rect 153910 660100 154000 660340
rect 154240 660100 154330 660340
rect 154570 660100 154680 660340
rect 154920 660100 155010 660340
rect 155250 660100 155340 660340
rect 155580 660100 155670 660340
rect 155910 660100 155930 660340
rect 144930 660010 155930 660100
rect 144930 659770 144950 660010
rect 145190 659770 145300 660010
rect 145540 659770 145630 660010
rect 145870 659770 145960 660010
rect 146200 659770 146290 660010
rect 146530 659770 146640 660010
rect 146880 659770 146970 660010
rect 147210 659770 147300 660010
rect 147540 659770 147630 660010
rect 147870 659770 147980 660010
rect 148220 659770 148310 660010
rect 148550 659770 148640 660010
rect 148880 659770 148970 660010
rect 149210 659770 149320 660010
rect 149560 659770 149650 660010
rect 149890 659770 149980 660010
rect 150220 659770 150310 660010
rect 150550 659770 150660 660010
rect 150900 659770 150990 660010
rect 151230 659770 151320 660010
rect 151560 659770 151650 660010
rect 151890 659770 152000 660010
rect 152240 659770 152330 660010
rect 152570 659770 152660 660010
rect 152900 659770 152990 660010
rect 153230 659770 153340 660010
rect 153580 659770 153670 660010
rect 153910 659770 154000 660010
rect 154240 659770 154330 660010
rect 154570 659770 154680 660010
rect 154920 659770 155010 660010
rect 155250 659770 155340 660010
rect 155580 659770 155670 660010
rect 155910 659770 155930 660010
rect 144930 659680 155930 659770
rect 144930 659440 144950 659680
rect 145190 659440 145300 659680
rect 145540 659440 145630 659680
rect 145870 659440 145960 659680
rect 146200 659440 146290 659680
rect 146530 659440 146640 659680
rect 146880 659440 146970 659680
rect 147210 659440 147300 659680
rect 147540 659440 147630 659680
rect 147870 659440 147980 659680
rect 148220 659440 148310 659680
rect 148550 659440 148640 659680
rect 148880 659440 148970 659680
rect 149210 659440 149320 659680
rect 149560 659440 149650 659680
rect 149890 659440 149980 659680
rect 150220 659440 150310 659680
rect 150550 659440 150660 659680
rect 150900 659440 150990 659680
rect 151230 659440 151320 659680
rect 151560 659440 151650 659680
rect 151890 659440 152000 659680
rect 152240 659440 152330 659680
rect 152570 659440 152660 659680
rect 152900 659440 152990 659680
rect 153230 659440 153340 659680
rect 153580 659440 153670 659680
rect 153910 659440 154000 659680
rect 154240 659440 154330 659680
rect 154570 659440 154680 659680
rect 154920 659440 155010 659680
rect 155250 659440 155340 659680
rect 155580 659440 155670 659680
rect 155910 659440 155930 659680
rect 144930 659350 155930 659440
rect 144930 659110 144950 659350
rect 145190 659110 145300 659350
rect 145540 659110 145630 659350
rect 145870 659110 145960 659350
rect 146200 659110 146290 659350
rect 146530 659110 146640 659350
rect 146880 659110 146970 659350
rect 147210 659110 147300 659350
rect 147540 659110 147630 659350
rect 147870 659110 147980 659350
rect 148220 659110 148310 659350
rect 148550 659110 148640 659350
rect 148880 659110 148970 659350
rect 149210 659110 149320 659350
rect 149560 659110 149650 659350
rect 149890 659110 149980 659350
rect 150220 659110 150310 659350
rect 150550 659110 150660 659350
rect 150900 659110 150990 659350
rect 151230 659110 151320 659350
rect 151560 659110 151650 659350
rect 151890 659110 152000 659350
rect 152240 659110 152330 659350
rect 152570 659110 152660 659350
rect 152900 659110 152990 659350
rect 153230 659110 153340 659350
rect 153580 659110 153670 659350
rect 153910 659110 154000 659350
rect 154240 659110 154330 659350
rect 154570 659110 154680 659350
rect 154920 659110 155010 659350
rect 155250 659110 155340 659350
rect 155580 659110 155670 659350
rect 155910 659110 155930 659350
rect 144930 659000 155930 659110
rect 144930 658760 144950 659000
rect 145190 658760 145300 659000
rect 145540 658760 145630 659000
rect 145870 658760 145960 659000
rect 146200 658760 146290 659000
rect 146530 658760 146640 659000
rect 146880 658760 146970 659000
rect 147210 658760 147300 659000
rect 147540 658760 147630 659000
rect 147870 658760 147980 659000
rect 148220 658760 148310 659000
rect 148550 658760 148640 659000
rect 148880 658760 148970 659000
rect 149210 658760 149320 659000
rect 149560 658760 149650 659000
rect 149890 658760 149980 659000
rect 150220 658760 150310 659000
rect 150550 658760 150660 659000
rect 150900 658760 150990 659000
rect 151230 658760 151320 659000
rect 151560 658760 151650 659000
rect 151890 658760 152000 659000
rect 152240 658760 152330 659000
rect 152570 658760 152660 659000
rect 152900 658760 152990 659000
rect 153230 658760 153340 659000
rect 153580 658760 153670 659000
rect 153910 658760 154000 659000
rect 154240 658760 154330 659000
rect 154570 658760 154680 659000
rect 154920 658760 155010 659000
rect 155250 658760 155340 659000
rect 155580 658760 155670 659000
rect 155910 658760 155930 659000
rect 144930 658670 155930 658760
rect 144930 658430 144950 658670
rect 145190 658430 145300 658670
rect 145540 658430 145630 658670
rect 145870 658430 145960 658670
rect 146200 658430 146290 658670
rect 146530 658430 146640 658670
rect 146880 658430 146970 658670
rect 147210 658430 147300 658670
rect 147540 658430 147630 658670
rect 147870 658430 147980 658670
rect 148220 658430 148310 658670
rect 148550 658430 148640 658670
rect 148880 658430 148970 658670
rect 149210 658430 149320 658670
rect 149560 658430 149650 658670
rect 149890 658430 149980 658670
rect 150220 658430 150310 658670
rect 150550 658430 150660 658670
rect 150900 658430 150990 658670
rect 151230 658430 151320 658670
rect 151560 658430 151650 658670
rect 151890 658430 152000 658670
rect 152240 658430 152330 658670
rect 152570 658430 152660 658670
rect 152900 658430 152990 658670
rect 153230 658430 153340 658670
rect 153580 658430 153670 658670
rect 153910 658430 154000 658670
rect 154240 658430 154330 658670
rect 154570 658430 154680 658670
rect 154920 658430 155010 658670
rect 155250 658430 155340 658670
rect 155580 658430 155670 658670
rect 155910 658430 155930 658670
rect 144930 658340 155930 658430
rect 144930 658100 144950 658340
rect 145190 658100 145300 658340
rect 145540 658100 145630 658340
rect 145870 658100 145960 658340
rect 146200 658100 146290 658340
rect 146530 658100 146640 658340
rect 146880 658100 146970 658340
rect 147210 658100 147300 658340
rect 147540 658100 147630 658340
rect 147870 658100 147980 658340
rect 148220 658100 148310 658340
rect 148550 658100 148640 658340
rect 148880 658100 148970 658340
rect 149210 658100 149320 658340
rect 149560 658100 149650 658340
rect 149890 658100 149980 658340
rect 150220 658100 150310 658340
rect 150550 658100 150660 658340
rect 150900 658100 150990 658340
rect 151230 658100 151320 658340
rect 151560 658100 151650 658340
rect 151890 658100 152000 658340
rect 152240 658100 152330 658340
rect 152570 658100 152660 658340
rect 152900 658100 152990 658340
rect 153230 658100 153340 658340
rect 153580 658100 153670 658340
rect 153910 658100 154000 658340
rect 154240 658100 154330 658340
rect 154570 658100 154680 658340
rect 154920 658100 155010 658340
rect 155250 658100 155340 658340
rect 155580 658100 155670 658340
rect 155910 658100 155930 658340
rect 144930 658010 155930 658100
rect 144930 657770 144950 658010
rect 145190 657770 145300 658010
rect 145540 657770 145630 658010
rect 145870 657770 145960 658010
rect 146200 657770 146290 658010
rect 146530 657770 146640 658010
rect 146880 657770 146970 658010
rect 147210 657770 147300 658010
rect 147540 657770 147630 658010
rect 147870 657770 147980 658010
rect 148220 657770 148310 658010
rect 148550 657770 148640 658010
rect 148880 657770 148970 658010
rect 149210 657770 149320 658010
rect 149560 657770 149650 658010
rect 149890 657770 149980 658010
rect 150220 657770 150310 658010
rect 150550 657770 150660 658010
rect 150900 657770 150990 658010
rect 151230 657770 151320 658010
rect 151560 657770 151650 658010
rect 151890 657770 152000 658010
rect 152240 657770 152330 658010
rect 152570 657770 152660 658010
rect 152900 657770 152990 658010
rect 153230 657770 153340 658010
rect 153580 657770 153670 658010
rect 153910 657770 154000 658010
rect 154240 657770 154330 658010
rect 154570 657770 154680 658010
rect 154920 657770 155010 658010
rect 155250 657770 155340 658010
rect 155580 657770 155670 658010
rect 155910 657770 155930 658010
rect 144930 657660 155930 657770
rect 144930 657420 144950 657660
rect 145190 657420 145300 657660
rect 145540 657420 145630 657660
rect 145870 657420 145960 657660
rect 146200 657420 146290 657660
rect 146530 657420 146640 657660
rect 146880 657420 146970 657660
rect 147210 657420 147300 657660
rect 147540 657420 147630 657660
rect 147870 657420 147980 657660
rect 148220 657420 148310 657660
rect 148550 657420 148640 657660
rect 148880 657420 148970 657660
rect 149210 657420 149320 657660
rect 149560 657420 149650 657660
rect 149890 657420 149980 657660
rect 150220 657420 150310 657660
rect 150550 657420 150660 657660
rect 150900 657420 150990 657660
rect 151230 657420 151320 657660
rect 151560 657420 151650 657660
rect 151890 657420 152000 657660
rect 152240 657420 152330 657660
rect 152570 657420 152660 657660
rect 152900 657420 152990 657660
rect 153230 657420 153340 657660
rect 153580 657420 153670 657660
rect 153910 657420 154000 657660
rect 154240 657420 154330 657660
rect 154570 657420 154680 657660
rect 154920 657420 155010 657660
rect 155250 657420 155340 657660
rect 155580 657420 155670 657660
rect 155910 657420 155930 657660
rect 144930 657330 155930 657420
rect 144930 657090 144950 657330
rect 145190 657090 145300 657330
rect 145540 657090 145630 657330
rect 145870 657090 145960 657330
rect 146200 657090 146290 657330
rect 146530 657090 146640 657330
rect 146880 657090 146970 657330
rect 147210 657090 147300 657330
rect 147540 657090 147630 657330
rect 147870 657090 147980 657330
rect 148220 657090 148310 657330
rect 148550 657090 148640 657330
rect 148880 657090 148970 657330
rect 149210 657090 149320 657330
rect 149560 657090 149650 657330
rect 149890 657090 149980 657330
rect 150220 657090 150310 657330
rect 150550 657090 150660 657330
rect 150900 657090 150990 657330
rect 151230 657090 151320 657330
rect 151560 657090 151650 657330
rect 151890 657090 152000 657330
rect 152240 657090 152330 657330
rect 152570 657090 152660 657330
rect 152900 657090 152990 657330
rect 153230 657090 153340 657330
rect 153580 657090 153670 657330
rect 153910 657090 154000 657330
rect 154240 657090 154330 657330
rect 154570 657090 154680 657330
rect 154920 657090 155010 657330
rect 155250 657090 155340 657330
rect 155580 657090 155670 657330
rect 155910 657090 155930 657330
rect 144930 657000 155930 657090
rect 144930 656760 144950 657000
rect 145190 656760 145300 657000
rect 145540 656760 145630 657000
rect 145870 656760 145960 657000
rect 146200 656760 146290 657000
rect 146530 656760 146640 657000
rect 146880 656760 146970 657000
rect 147210 656760 147300 657000
rect 147540 656760 147630 657000
rect 147870 656760 147980 657000
rect 148220 656760 148310 657000
rect 148550 656760 148640 657000
rect 148880 656760 148970 657000
rect 149210 656760 149320 657000
rect 149560 656760 149650 657000
rect 149890 656760 149980 657000
rect 150220 656760 150310 657000
rect 150550 656760 150660 657000
rect 150900 656760 150990 657000
rect 151230 656760 151320 657000
rect 151560 656760 151650 657000
rect 151890 656760 152000 657000
rect 152240 656760 152330 657000
rect 152570 656760 152660 657000
rect 152900 656760 152990 657000
rect 153230 656760 153340 657000
rect 153580 656760 153670 657000
rect 153910 656760 154000 657000
rect 154240 656760 154330 657000
rect 154570 656760 154680 657000
rect 154920 656760 155010 657000
rect 155250 656760 155340 657000
rect 155580 656760 155670 657000
rect 155910 656760 155930 657000
rect 144930 656670 155930 656760
rect 144930 656430 144950 656670
rect 145190 656430 145300 656670
rect 145540 656430 145630 656670
rect 145870 656430 145960 656670
rect 146200 656430 146290 656670
rect 146530 656430 146640 656670
rect 146880 656430 146970 656670
rect 147210 656430 147300 656670
rect 147540 656430 147630 656670
rect 147870 656430 147980 656670
rect 148220 656430 148310 656670
rect 148550 656430 148640 656670
rect 148880 656430 148970 656670
rect 149210 656430 149320 656670
rect 149560 656430 149650 656670
rect 149890 656430 149980 656670
rect 150220 656430 150310 656670
rect 150550 656430 150660 656670
rect 150900 656430 150990 656670
rect 151230 656430 151320 656670
rect 151560 656430 151650 656670
rect 151890 656430 152000 656670
rect 152240 656430 152330 656670
rect 152570 656430 152660 656670
rect 152900 656430 152990 656670
rect 153230 656430 153340 656670
rect 153580 656430 153670 656670
rect 153910 656430 154000 656670
rect 154240 656430 154330 656670
rect 154570 656430 154680 656670
rect 154920 656430 155010 656670
rect 155250 656430 155340 656670
rect 155580 656430 155670 656670
rect 155910 656430 155930 656670
rect 144930 656320 155930 656430
rect 144930 656080 144950 656320
rect 145190 656080 145300 656320
rect 145540 656080 145630 656320
rect 145870 656080 145960 656320
rect 146200 656080 146290 656320
rect 146530 656080 146640 656320
rect 146880 656080 146970 656320
rect 147210 656080 147300 656320
rect 147540 656080 147630 656320
rect 147870 656080 147980 656320
rect 148220 656080 148310 656320
rect 148550 656080 148640 656320
rect 148880 656080 148970 656320
rect 149210 656080 149320 656320
rect 149560 656080 149650 656320
rect 149890 656080 149980 656320
rect 150220 656080 150310 656320
rect 150550 656080 150660 656320
rect 150900 656080 150990 656320
rect 151230 656080 151320 656320
rect 151560 656080 151650 656320
rect 151890 656080 152000 656320
rect 152240 656080 152330 656320
rect 152570 656080 152660 656320
rect 152900 656080 152990 656320
rect 153230 656080 153340 656320
rect 153580 656080 153670 656320
rect 153910 656080 154000 656320
rect 154240 656080 154330 656320
rect 154570 656080 154680 656320
rect 154920 656080 155010 656320
rect 155250 656080 155340 656320
rect 155580 656080 155670 656320
rect 155910 656080 155930 656320
rect 144930 655990 155930 656080
rect 144930 655750 144950 655990
rect 145190 655750 145300 655990
rect 145540 655750 145630 655990
rect 145870 655750 145960 655990
rect 146200 655750 146290 655990
rect 146530 655750 146640 655990
rect 146880 655750 146970 655990
rect 147210 655750 147300 655990
rect 147540 655750 147630 655990
rect 147870 655750 147980 655990
rect 148220 655750 148310 655990
rect 148550 655750 148640 655990
rect 148880 655750 148970 655990
rect 149210 655750 149320 655990
rect 149560 655750 149650 655990
rect 149890 655750 149980 655990
rect 150220 655750 150310 655990
rect 150550 655750 150660 655990
rect 150900 655750 150990 655990
rect 151230 655750 151320 655990
rect 151560 655750 151650 655990
rect 151890 655750 152000 655990
rect 152240 655750 152330 655990
rect 152570 655750 152660 655990
rect 152900 655750 152990 655990
rect 153230 655750 153340 655990
rect 153580 655750 153670 655990
rect 153910 655750 154000 655990
rect 154240 655750 154330 655990
rect 154570 655750 154680 655990
rect 154920 655750 155010 655990
rect 155250 655750 155340 655990
rect 155580 655750 155670 655990
rect 155910 655750 155930 655990
rect 144930 655660 155930 655750
rect 144930 655420 144950 655660
rect 145190 655420 145300 655660
rect 145540 655420 145630 655660
rect 145870 655420 145960 655660
rect 146200 655420 146290 655660
rect 146530 655420 146640 655660
rect 146880 655420 146970 655660
rect 147210 655420 147300 655660
rect 147540 655420 147630 655660
rect 147870 655420 147980 655660
rect 148220 655420 148310 655660
rect 148550 655420 148640 655660
rect 148880 655420 148970 655660
rect 149210 655420 149320 655660
rect 149560 655420 149650 655660
rect 149890 655420 149980 655660
rect 150220 655420 150310 655660
rect 150550 655420 150660 655660
rect 150900 655420 150990 655660
rect 151230 655420 151320 655660
rect 151560 655420 151650 655660
rect 151890 655420 152000 655660
rect 152240 655420 152330 655660
rect 152570 655420 152660 655660
rect 152900 655420 152990 655660
rect 153230 655420 153340 655660
rect 153580 655420 153670 655660
rect 153910 655420 154000 655660
rect 154240 655420 154330 655660
rect 154570 655420 154680 655660
rect 154920 655420 155010 655660
rect 155250 655420 155340 655660
rect 155580 655420 155670 655660
rect 155910 655420 155930 655660
rect 144930 655330 155930 655420
rect 144930 655090 144950 655330
rect 145190 655090 145300 655330
rect 145540 655090 145630 655330
rect 145870 655090 145960 655330
rect 146200 655090 146290 655330
rect 146530 655090 146640 655330
rect 146880 655090 146970 655330
rect 147210 655090 147300 655330
rect 147540 655090 147630 655330
rect 147870 655090 147980 655330
rect 148220 655090 148310 655330
rect 148550 655090 148640 655330
rect 148880 655090 148970 655330
rect 149210 655090 149320 655330
rect 149560 655090 149650 655330
rect 149890 655090 149980 655330
rect 150220 655090 150310 655330
rect 150550 655090 150660 655330
rect 150900 655090 150990 655330
rect 151230 655090 151320 655330
rect 151560 655090 151650 655330
rect 151890 655090 152000 655330
rect 152240 655090 152330 655330
rect 152570 655090 152660 655330
rect 152900 655090 152990 655330
rect 153230 655090 153340 655330
rect 153580 655090 153670 655330
rect 153910 655090 154000 655330
rect 154240 655090 154330 655330
rect 154570 655090 154680 655330
rect 154920 655090 155010 655330
rect 155250 655090 155340 655330
rect 155580 655090 155670 655330
rect 155910 655090 155930 655330
rect 144930 654980 155930 655090
rect 144930 654740 144950 654980
rect 145190 654740 145300 654980
rect 145540 654740 145630 654980
rect 145870 654740 145960 654980
rect 146200 654740 146290 654980
rect 146530 654740 146640 654980
rect 146880 654740 146970 654980
rect 147210 654740 147300 654980
rect 147540 654740 147630 654980
rect 147870 654740 147980 654980
rect 148220 654740 148310 654980
rect 148550 654740 148640 654980
rect 148880 654740 148970 654980
rect 149210 654740 149320 654980
rect 149560 654740 149650 654980
rect 149890 654740 149980 654980
rect 150220 654740 150310 654980
rect 150550 654740 150660 654980
rect 150900 654740 150990 654980
rect 151230 654740 151320 654980
rect 151560 654740 151650 654980
rect 151890 654740 152000 654980
rect 152240 654740 152330 654980
rect 152570 654740 152660 654980
rect 152900 654740 152990 654980
rect 153230 654740 153340 654980
rect 153580 654740 153670 654980
rect 153910 654740 154000 654980
rect 154240 654740 154330 654980
rect 154570 654740 154680 654980
rect 154920 654740 155010 654980
rect 155250 654740 155340 654980
rect 155580 654740 155670 654980
rect 155910 654740 155930 654980
rect 144930 654650 155930 654740
rect 144930 654410 144950 654650
rect 145190 654410 145300 654650
rect 145540 654410 145630 654650
rect 145870 654410 145960 654650
rect 146200 654410 146290 654650
rect 146530 654410 146640 654650
rect 146880 654410 146970 654650
rect 147210 654410 147300 654650
rect 147540 654410 147630 654650
rect 147870 654410 147980 654650
rect 148220 654410 148310 654650
rect 148550 654410 148640 654650
rect 148880 654410 148970 654650
rect 149210 654410 149320 654650
rect 149560 654410 149650 654650
rect 149890 654410 149980 654650
rect 150220 654410 150310 654650
rect 150550 654410 150660 654650
rect 150900 654410 150990 654650
rect 151230 654410 151320 654650
rect 151560 654410 151650 654650
rect 151890 654410 152000 654650
rect 152240 654410 152330 654650
rect 152570 654410 152660 654650
rect 152900 654410 152990 654650
rect 153230 654410 153340 654650
rect 153580 654410 153670 654650
rect 153910 654410 154000 654650
rect 154240 654410 154330 654650
rect 154570 654410 154680 654650
rect 154920 654410 155010 654650
rect 155250 654410 155340 654650
rect 155580 654410 155670 654650
rect 155910 654410 155930 654650
rect 144930 654320 155930 654410
rect 144930 654080 144950 654320
rect 145190 654080 145300 654320
rect 145540 654080 145630 654320
rect 145870 654080 145960 654320
rect 146200 654080 146290 654320
rect 146530 654080 146640 654320
rect 146880 654080 146970 654320
rect 147210 654080 147300 654320
rect 147540 654080 147630 654320
rect 147870 654080 147980 654320
rect 148220 654080 148310 654320
rect 148550 654080 148640 654320
rect 148880 654080 148970 654320
rect 149210 654080 149320 654320
rect 149560 654080 149650 654320
rect 149890 654080 149980 654320
rect 150220 654080 150310 654320
rect 150550 654080 150660 654320
rect 150900 654080 150990 654320
rect 151230 654080 151320 654320
rect 151560 654080 151650 654320
rect 151890 654080 152000 654320
rect 152240 654080 152330 654320
rect 152570 654080 152660 654320
rect 152900 654080 152990 654320
rect 153230 654080 153340 654320
rect 153580 654080 153670 654320
rect 153910 654080 154000 654320
rect 154240 654080 154330 654320
rect 154570 654080 154680 654320
rect 154920 654080 155010 654320
rect 155250 654080 155340 654320
rect 155580 654080 155670 654320
rect 155910 654080 155930 654320
rect 144930 653990 155930 654080
rect 144930 653750 144950 653990
rect 145190 653750 145300 653990
rect 145540 653750 145630 653990
rect 145870 653750 145960 653990
rect 146200 653750 146290 653990
rect 146530 653750 146640 653990
rect 146880 653750 146970 653990
rect 147210 653750 147300 653990
rect 147540 653750 147630 653990
rect 147870 653750 147980 653990
rect 148220 653750 148310 653990
rect 148550 653750 148640 653990
rect 148880 653750 148970 653990
rect 149210 653750 149320 653990
rect 149560 653750 149650 653990
rect 149890 653750 149980 653990
rect 150220 653750 150310 653990
rect 150550 653750 150660 653990
rect 150900 653750 150990 653990
rect 151230 653750 151320 653990
rect 151560 653750 151650 653990
rect 151890 653750 152000 653990
rect 152240 653750 152330 653990
rect 152570 653750 152660 653990
rect 152900 653750 152990 653990
rect 153230 653750 153340 653990
rect 153580 653750 153670 653990
rect 153910 653750 154000 653990
rect 154240 653750 154330 653990
rect 154570 653750 154680 653990
rect 154920 653750 155010 653990
rect 155250 653750 155340 653990
rect 155580 653750 155670 653990
rect 155910 653750 155930 653990
rect 144930 653640 155930 653750
rect 144930 653400 144950 653640
rect 145190 653400 145300 653640
rect 145540 653400 145630 653640
rect 145870 653400 145960 653640
rect 146200 653400 146290 653640
rect 146530 653400 146640 653640
rect 146880 653400 146970 653640
rect 147210 653400 147300 653640
rect 147540 653400 147630 653640
rect 147870 653400 147980 653640
rect 148220 653400 148310 653640
rect 148550 653400 148640 653640
rect 148880 653400 148970 653640
rect 149210 653400 149320 653640
rect 149560 653400 149650 653640
rect 149890 653400 149980 653640
rect 150220 653400 150310 653640
rect 150550 653400 150660 653640
rect 150900 653400 150990 653640
rect 151230 653400 151320 653640
rect 151560 653400 151650 653640
rect 151890 653400 152000 653640
rect 152240 653400 152330 653640
rect 152570 653400 152660 653640
rect 152900 653400 152990 653640
rect 153230 653400 153340 653640
rect 153580 653400 153670 653640
rect 153910 653400 154000 653640
rect 154240 653400 154330 653640
rect 154570 653400 154680 653640
rect 154920 653400 155010 653640
rect 155250 653400 155340 653640
rect 155580 653400 155670 653640
rect 155910 653400 155930 653640
rect 144930 653310 155930 653400
rect 144930 653070 144950 653310
rect 145190 653070 145300 653310
rect 145540 653070 145630 653310
rect 145870 653070 145960 653310
rect 146200 653070 146290 653310
rect 146530 653070 146640 653310
rect 146880 653070 146970 653310
rect 147210 653070 147300 653310
rect 147540 653070 147630 653310
rect 147870 653070 147980 653310
rect 148220 653070 148310 653310
rect 148550 653070 148640 653310
rect 148880 653070 148970 653310
rect 149210 653070 149320 653310
rect 149560 653070 149650 653310
rect 149890 653070 149980 653310
rect 150220 653070 150310 653310
rect 150550 653070 150660 653310
rect 150900 653070 150990 653310
rect 151230 653070 151320 653310
rect 151560 653070 151650 653310
rect 151890 653070 152000 653310
rect 152240 653070 152330 653310
rect 152570 653070 152660 653310
rect 152900 653070 152990 653310
rect 153230 653070 153340 653310
rect 153580 653070 153670 653310
rect 153910 653070 154000 653310
rect 154240 653070 154330 653310
rect 154570 653070 154680 653310
rect 154920 653070 155010 653310
rect 155250 653070 155340 653310
rect 155580 653070 155670 653310
rect 155910 653070 155930 653310
rect 144930 652980 155930 653070
rect 144930 652740 144950 652980
rect 145190 652740 145300 652980
rect 145540 652740 145630 652980
rect 145870 652740 145960 652980
rect 146200 652740 146290 652980
rect 146530 652740 146640 652980
rect 146880 652740 146970 652980
rect 147210 652740 147300 652980
rect 147540 652740 147630 652980
rect 147870 652740 147980 652980
rect 148220 652740 148310 652980
rect 148550 652740 148640 652980
rect 148880 652740 148970 652980
rect 149210 652740 149320 652980
rect 149560 652740 149650 652980
rect 149890 652740 149980 652980
rect 150220 652740 150310 652980
rect 150550 652740 150660 652980
rect 150900 652740 150990 652980
rect 151230 652740 151320 652980
rect 151560 652740 151650 652980
rect 151890 652740 152000 652980
rect 152240 652740 152330 652980
rect 152570 652740 152660 652980
rect 152900 652740 152990 652980
rect 153230 652740 153340 652980
rect 153580 652740 153670 652980
rect 153910 652740 154000 652980
rect 154240 652740 154330 652980
rect 154570 652740 154680 652980
rect 154920 652740 155010 652980
rect 155250 652740 155340 652980
rect 155580 652740 155670 652980
rect 155910 652740 155930 652980
rect 144930 652650 155930 652740
rect 144930 652410 144950 652650
rect 145190 652410 145300 652650
rect 145540 652410 145630 652650
rect 145870 652410 145960 652650
rect 146200 652410 146290 652650
rect 146530 652410 146640 652650
rect 146880 652410 146970 652650
rect 147210 652410 147300 652650
rect 147540 652410 147630 652650
rect 147870 652410 147980 652650
rect 148220 652410 148310 652650
rect 148550 652410 148640 652650
rect 148880 652410 148970 652650
rect 149210 652410 149320 652650
rect 149560 652410 149650 652650
rect 149890 652410 149980 652650
rect 150220 652410 150310 652650
rect 150550 652410 150660 652650
rect 150900 652410 150990 652650
rect 151230 652410 151320 652650
rect 151560 652410 151650 652650
rect 151890 652410 152000 652650
rect 152240 652410 152330 652650
rect 152570 652410 152660 652650
rect 152900 652410 152990 652650
rect 153230 652410 153340 652650
rect 153580 652410 153670 652650
rect 153910 652410 154000 652650
rect 154240 652410 154330 652650
rect 154570 652410 154680 652650
rect 154920 652410 155010 652650
rect 155250 652410 155340 652650
rect 155580 652410 155670 652650
rect 155910 652410 155930 652650
rect 144930 652300 155930 652410
rect 144930 652060 144950 652300
rect 145190 652060 145300 652300
rect 145540 652060 145630 652300
rect 145870 652060 145960 652300
rect 146200 652060 146290 652300
rect 146530 652060 146640 652300
rect 146880 652060 146970 652300
rect 147210 652060 147300 652300
rect 147540 652060 147630 652300
rect 147870 652060 147980 652300
rect 148220 652060 148310 652300
rect 148550 652060 148640 652300
rect 148880 652060 148970 652300
rect 149210 652060 149320 652300
rect 149560 652060 149650 652300
rect 149890 652060 149980 652300
rect 150220 652060 150310 652300
rect 150550 652060 150660 652300
rect 150900 652060 150990 652300
rect 151230 652060 151320 652300
rect 151560 652060 151650 652300
rect 151890 652060 152000 652300
rect 152240 652060 152330 652300
rect 152570 652060 152660 652300
rect 152900 652060 152990 652300
rect 153230 652060 153340 652300
rect 153580 652060 153670 652300
rect 153910 652060 154000 652300
rect 154240 652060 154330 652300
rect 154570 652060 154680 652300
rect 154920 652060 155010 652300
rect 155250 652060 155340 652300
rect 155580 652060 155670 652300
rect 155910 652060 155930 652300
rect 144930 651970 155930 652060
rect 144930 651730 144950 651970
rect 145190 651730 145300 651970
rect 145540 651730 145630 651970
rect 145870 651730 145960 651970
rect 146200 651730 146290 651970
rect 146530 651730 146640 651970
rect 146880 651730 146970 651970
rect 147210 651730 147300 651970
rect 147540 651730 147630 651970
rect 147870 651730 147980 651970
rect 148220 651730 148310 651970
rect 148550 651730 148640 651970
rect 148880 651730 148970 651970
rect 149210 651730 149320 651970
rect 149560 651730 149650 651970
rect 149890 651730 149980 651970
rect 150220 651730 150310 651970
rect 150550 651730 150660 651970
rect 150900 651730 150990 651970
rect 151230 651730 151320 651970
rect 151560 651730 151650 651970
rect 151890 651730 152000 651970
rect 152240 651730 152330 651970
rect 152570 651730 152660 651970
rect 152900 651730 152990 651970
rect 153230 651730 153340 651970
rect 153580 651730 153670 651970
rect 153910 651730 154000 651970
rect 154240 651730 154330 651970
rect 154570 651730 154680 651970
rect 154920 651730 155010 651970
rect 155250 651730 155340 651970
rect 155580 651730 155670 651970
rect 155910 651730 155930 651970
rect 144930 651640 155930 651730
rect 144930 651400 144950 651640
rect 145190 651400 145300 651640
rect 145540 651400 145630 651640
rect 145870 651400 145960 651640
rect 146200 651400 146290 651640
rect 146530 651400 146640 651640
rect 146880 651400 146970 651640
rect 147210 651400 147300 651640
rect 147540 651400 147630 651640
rect 147870 651400 147980 651640
rect 148220 651400 148310 651640
rect 148550 651400 148640 651640
rect 148880 651400 148970 651640
rect 149210 651400 149320 651640
rect 149560 651400 149650 651640
rect 149890 651400 149980 651640
rect 150220 651400 150310 651640
rect 150550 651400 150660 651640
rect 150900 651400 150990 651640
rect 151230 651400 151320 651640
rect 151560 651400 151650 651640
rect 151890 651400 152000 651640
rect 152240 651400 152330 651640
rect 152570 651400 152660 651640
rect 152900 651400 152990 651640
rect 153230 651400 153340 651640
rect 153580 651400 153670 651640
rect 153910 651400 154000 651640
rect 154240 651400 154330 651640
rect 154570 651400 154680 651640
rect 154920 651400 155010 651640
rect 155250 651400 155340 651640
rect 155580 651400 155670 651640
rect 155910 651400 155930 651640
rect 144930 651310 155930 651400
rect 144930 651070 144950 651310
rect 145190 651070 145300 651310
rect 145540 651070 145630 651310
rect 145870 651070 145960 651310
rect 146200 651070 146290 651310
rect 146530 651070 146640 651310
rect 146880 651070 146970 651310
rect 147210 651070 147300 651310
rect 147540 651070 147630 651310
rect 147870 651070 147980 651310
rect 148220 651070 148310 651310
rect 148550 651070 148640 651310
rect 148880 651070 148970 651310
rect 149210 651070 149320 651310
rect 149560 651070 149650 651310
rect 149890 651070 149980 651310
rect 150220 651070 150310 651310
rect 150550 651070 150660 651310
rect 150900 651070 150990 651310
rect 151230 651070 151320 651310
rect 151560 651070 151650 651310
rect 151890 651070 152000 651310
rect 152240 651070 152330 651310
rect 152570 651070 152660 651310
rect 152900 651070 152990 651310
rect 153230 651070 153340 651310
rect 153580 651070 153670 651310
rect 153910 651070 154000 651310
rect 154240 651070 154330 651310
rect 154570 651070 154680 651310
rect 154920 651070 155010 651310
rect 155250 651070 155340 651310
rect 155580 651070 155670 651310
rect 155910 651070 155930 651310
rect 144930 650960 155930 651070
rect 144930 650720 144950 650960
rect 145190 650720 145300 650960
rect 145540 650720 145630 650960
rect 145870 650720 145960 650960
rect 146200 650720 146290 650960
rect 146530 650720 146640 650960
rect 146880 650720 146970 650960
rect 147210 650720 147300 650960
rect 147540 650720 147630 650960
rect 147870 650720 147980 650960
rect 148220 650720 148310 650960
rect 148550 650720 148640 650960
rect 148880 650720 148970 650960
rect 149210 650720 149320 650960
rect 149560 650720 149650 650960
rect 149890 650720 149980 650960
rect 150220 650720 150310 650960
rect 150550 650720 150660 650960
rect 150900 650720 150990 650960
rect 151230 650720 151320 650960
rect 151560 650720 151650 650960
rect 151890 650720 152000 650960
rect 152240 650720 152330 650960
rect 152570 650720 152660 650960
rect 152900 650720 152990 650960
rect 153230 650720 153340 650960
rect 153580 650720 153670 650960
rect 153910 650720 154000 650960
rect 154240 650720 154330 650960
rect 154570 650720 154680 650960
rect 154920 650720 155010 650960
rect 155250 650720 155340 650960
rect 155580 650720 155670 650960
rect 155910 650720 155930 650960
rect 144930 650630 155930 650720
rect 144930 650390 144950 650630
rect 145190 650390 145300 650630
rect 145540 650390 145630 650630
rect 145870 650390 145960 650630
rect 146200 650390 146290 650630
rect 146530 650390 146640 650630
rect 146880 650390 146970 650630
rect 147210 650390 147300 650630
rect 147540 650390 147630 650630
rect 147870 650390 147980 650630
rect 148220 650390 148310 650630
rect 148550 650390 148640 650630
rect 148880 650390 148970 650630
rect 149210 650390 149320 650630
rect 149560 650390 149650 650630
rect 149890 650390 149980 650630
rect 150220 650390 150310 650630
rect 150550 650390 150660 650630
rect 150900 650390 150990 650630
rect 151230 650390 151320 650630
rect 151560 650390 151650 650630
rect 151890 650390 152000 650630
rect 152240 650390 152330 650630
rect 152570 650390 152660 650630
rect 152900 650390 152990 650630
rect 153230 650390 153340 650630
rect 153580 650390 153670 650630
rect 153910 650390 154000 650630
rect 154240 650390 154330 650630
rect 154570 650390 154680 650630
rect 154920 650390 155010 650630
rect 155250 650390 155340 650630
rect 155580 650390 155670 650630
rect 155910 650390 155930 650630
rect 144930 650300 155930 650390
rect 144930 650060 144950 650300
rect 145190 650060 145300 650300
rect 145540 650060 145630 650300
rect 145870 650060 145960 650300
rect 146200 650060 146290 650300
rect 146530 650060 146640 650300
rect 146880 650060 146970 650300
rect 147210 650060 147300 650300
rect 147540 650060 147630 650300
rect 147870 650060 147980 650300
rect 148220 650060 148310 650300
rect 148550 650060 148640 650300
rect 148880 650060 148970 650300
rect 149210 650060 149320 650300
rect 149560 650060 149650 650300
rect 149890 650060 149980 650300
rect 150220 650060 150310 650300
rect 150550 650060 150660 650300
rect 150900 650060 150990 650300
rect 151230 650060 151320 650300
rect 151560 650060 151650 650300
rect 151890 650060 152000 650300
rect 152240 650060 152330 650300
rect 152570 650060 152660 650300
rect 152900 650060 152990 650300
rect 153230 650060 153340 650300
rect 153580 650060 153670 650300
rect 153910 650060 154000 650300
rect 154240 650060 154330 650300
rect 154570 650060 154680 650300
rect 154920 650060 155010 650300
rect 155250 650060 155340 650300
rect 155580 650060 155670 650300
rect 155910 650060 155930 650300
rect 144930 649970 155930 650060
rect 144930 649730 144950 649970
rect 145190 649730 145300 649970
rect 145540 649730 145630 649970
rect 145870 649730 145960 649970
rect 146200 649730 146290 649970
rect 146530 649730 146640 649970
rect 146880 649730 146970 649970
rect 147210 649730 147300 649970
rect 147540 649730 147630 649970
rect 147870 649730 147980 649970
rect 148220 649730 148310 649970
rect 148550 649730 148640 649970
rect 148880 649730 148970 649970
rect 149210 649730 149320 649970
rect 149560 649730 149650 649970
rect 149890 649730 149980 649970
rect 150220 649730 150310 649970
rect 150550 649730 150660 649970
rect 150900 649730 150990 649970
rect 151230 649730 151320 649970
rect 151560 649730 151650 649970
rect 151890 649730 152000 649970
rect 152240 649730 152330 649970
rect 152570 649730 152660 649970
rect 152900 649730 152990 649970
rect 153230 649730 153340 649970
rect 153580 649730 153670 649970
rect 153910 649730 154000 649970
rect 154240 649730 154330 649970
rect 154570 649730 154680 649970
rect 154920 649730 155010 649970
rect 155250 649730 155340 649970
rect 155580 649730 155670 649970
rect 155910 649730 155930 649970
rect 144930 649620 155930 649730
rect 144930 649380 144950 649620
rect 145190 649380 145300 649620
rect 145540 649380 145630 649620
rect 145870 649380 145960 649620
rect 146200 649380 146290 649620
rect 146530 649380 146640 649620
rect 146880 649380 146970 649620
rect 147210 649380 147300 649620
rect 147540 649380 147630 649620
rect 147870 649380 147980 649620
rect 148220 649380 148310 649620
rect 148550 649380 148640 649620
rect 148880 649380 148970 649620
rect 149210 649380 149320 649620
rect 149560 649380 149650 649620
rect 149890 649380 149980 649620
rect 150220 649380 150310 649620
rect 150550 649380 150660 649620
rect 150900 649380 150990 649620
rect 151230 649380 151320 649620
rect 151560 649380 151650 649620
rect 151890 649380 152000 649620
rect 152240 649380 152330 649620
rect 152570 649380 152660 649620
rect 152900 649380 152990 649620
rect 153230 649380 153340 649620
rect 153580 649380 153670 649620
rect 153910 649380 154000 649620
rect 154240 649380 154330 649620
rect 154570 649380 154680 649620
rect 154920 649380 155010 649620
rect 155250 649380 155340 649620
rect 155580 649380 155670 649620
rect 155910 649380 155930 649620
rect 144930 649360 155930 649380
<< mimcap2contact >>
rect 110810 694600 111050 694840
rect 111140 694600 111380 694840
rect 111470 694600 111710 694840
rect 111800 694600 112040 694840
rect 112150 694600 112390 694840
rect 112480 694600 112720 694840
rect 112810 694600 113050 694840
rect 113140 694600 113380 694840
rect 113490 694600 113730 694840
rect 113820 694600 114060 694840
rect 114150 694600 114390 694840
rect 114480 694600 114720 694840
rect 114830 694600 115070 694840
rect 115160 694600 115400 694840
rect 115490 694600 115730 694840
rect 115820 694600 116060 694840
rect 116170 694600 116410 694840
rect 116500 694600 116740 694840
rect 116830 694600 117070 694840
rect 117160 694600 117400 694840
rect 117510 694600 117750 694840
rect 117840 694600 118080 694840
rect 118170 694600 118410 694840
rect 118500 694600 118740 694840
rect 118850 694600 119090 694840
rect 119180 694600 119420 694840
rect 119510 694600 119750 694840
rect 119840 694600 120080 694840
rect 120190 694600 120430 694840
rect 120520 694600 120760 694840
rect 120850 694600 121090 694840
rect 121180 694600 121420 694840
rect 121530 694600 121770 694840
rect 110810 694250 111050 694490
rect 111140 694250 111380 694490
rect 111470 694250 111710 694490
rect 111800 694250 112040 694490
rect 112150 694250 112390 694490
rect 112480 694250 112720 694490
rect 112810 694250 113050 694490
rect 113140 694250 113380 694490
rect 113490 694250 113730 694490
rect 113820 694250 114060 694490
rect 114150 694250 114390 694490
rect 114480 694250 114720 694490
rect 114830 694250 115070 694490
rect 115160 694250 115400 694490
rect 115490 694250 115730 694490
rect 115820 694250 116060 694490
rect 116170 694250 116410 694490
rect 116500 694250 116740 694490
rect 116830 694250 117070 694490
rect 117160 694250 117400 694490
rect 117510 694250 117750 694490
rect 117840 694250 118080 694490
rect 118170 694250 118410 694490
rect 118500 694250 118740 694490
rect 118850 694250 119090 694490
rect 119180 694250 119420 694490
rect 119510 694250 119750 694490
rect 119840 694250 120080 694490
rect 120190 694250 120430 694490
rect 120520 694250 120760 694490
rect 120850 694250 121090 694490
rect 121180 694250 121420 694490
rect 121530 694250 121770 694490
rect 110810 693920 111050 694160
rect 111140 693920 111380 694160
rect 111470 693920 111710 694160
rect 111800 693920 112040 694160
rect 112150 693920 112390 694160
rect 112480 693920 112720 694160
rect 112810 693920 113050 694160
rect 113140 693920 113380 694160
rect 113490 693920 113730 694160
rect 113820 693920 114060 694160
rect 114150 693920 114390 694160
rect 114480 693920 114720 694160
rect 114830 693920 115070 694160
rect 115160 693920 115400 694160
rect 115490 693920 115730 694160
rect 115820 693920 116060 694160
rect 116170 693920 116410 694160
rect 116500 693920 116740 694160
rect 116830 693920 117070 694160
rect 117160 693920 117400 694160
rect 117510 693920 117750 694160
rect 117840 693920 118080 694160
rect 118170 693920 118410 694160
rect 118500 693920 118740 694160
rect 118850 693920 119090 694160
rect 119180 693920 119420 694160
rect 119510 693920 119750 694160
rect 119840 693920 120080 694160
rect 120190 693920 120430 694160
rect 120520 693920 120760 694160
rect 120850 693920 121090 694160
rect 121180 693920 121420 694160
rect 121530 693920 121770 694160
rect 110810 693590 111050 693830
rect 111140 693590 111380 693830
rect 111470 693590 111710 693830
rect 111800 693590 112040 693830
rect 112150 693590 112390 693830
rect 112480 693590 112720 693830
rect 112810 693590 113050 693830
rect 113140 693590 113380 693830
rect 113490 693590 113730 693830
rect 113820 693590 114060 693830
rect 114150 693590 114390 693830
rect 114480 693590 114720 693830
rect 114830 693590 115070 693830
rect 115160 693590 115400 693830
rect 115490 693590 115730 693830
rect 115820 693590 116060 693830
rect 116170 693590 116410 693830
rect 116500 693590 116740 693830
rect 116830 693590 117070 693830
rect 117160 693590 117400 693830
rect 117510 693590 117750 693830
rect 117840 693590 118080 693830
rect 118170 693590 118410 693830
rect 118500 693590 118740 693830
rect 118850 693590 119090 693830
rect 119180 693590 119420 693830
rect 119510 693590 119750 693830
rect 119840 693590 120080 693830
rect 120190 693590 120430 693830
rect 120520 693590 120760 693830
rect 120850 693590 121090 693830
rect 121180 693590 121420 693830
rect 121530 693590 121770 693830
rect 110810 693260 111050 693500
rect 111140 693260 111380 693500
rect 111470 693260 111710 693500
rect 111800 693260 112040 693500
rect 112150 693260 112390 693500
rect 112480 693260 112720 693500
rect 112810 693260 113050 693500
rect 113140 693260 113380 693500
rect 113490 693260 113730 693500
rect 113820 693260 114060 693500
rect 114150 693260 114390 693500
rect 114480 693260 114720 693500
rect 114830 693260 115070 693500
rect 115160 693260 115400 693500
rect 115490 693260 115730 693500
rect 115820 693260 116060 693500
rect 116170 693260 116410 693500
rect 116500 693260 116740 693500
rect 116830 693260 117070 693500
rect 117160 693260 117400 693500
rect 117510 693260 117750 693500
rect 117840 693260 118080 693500
rect 118170 693260 118410 693500
rect 118500 693260 118740 693500
rect 118850 693260 119090 693500
rect 119180 693260 119420 693500
rect 119510 693260 119750 693500
rect 119840 693260 120080 693500
rect 120190 693260 120430 693500
rect 120520 693260 120760 693500
rect 120850 693260 121090 693500
rect 121180 693260 121420 693500
rect 121530 693260 121770 693500
rect 110810 692910 111050 693150
rect 111140 692910 111380 693150
rect 111470 692910 111710 693150
rect 111800 692910 112040 693150
rect 112150 692910 112390 693150
rect 112480 692910 112720 693150
rect 112810 692910 113050 693150
rect 113140 692910 113380 693150
rect 113490 692910 113730 693150
rect 113820 692910 114060 693150
rect 114150 692910 114390 693150
rect 114480 692910 114720 693150
rect 114830 692910 115070 693150
rect 115160 692910 115400 693150
rect 115490 692910 115730 693150
rect 115820 692910 116060 693150
rect 116170 692910 116410 693150
rect 116500 692910 116740 693150
rect 116830 692910 117070 693150
rect 117160 692910 117400 693150
rect 117510 692910 117750 693150
rect 117840 692910 118080 693150
rect 118170 692910 118410 693150
rect 118500 692910 118740 693150
rect 118850 692910 119090 693150
rect 119180 692910 119420 693150
rect 119510 692910 119750 693150
rect 119840 692910 120080 693150
rect 120190 692910 120430 693150
rect 120520 692910 120760 693150
rect 120850 692910 121090 693150
rect 121180 692910 121420 693150
rect 121530 692910 121770 693150
rect 110810 692580 111050 692820
rect 111140 692580 111380 692820
rect 111470 692580 111710 692820
rect 111800 692580 112040 692820
rect 112150 692580 112390 692820
rect 112480 692580 112720 692820
rect 112810 692580 113050 692820
rect 113140 692580 113380 692820
rect 113490 692580 113730 692820
rect 113820 692580 114060 692820
rect 114150 692580 114390 692820
rect 114480 692580 114720 692820
rect 114830 692580 115070 692820
rect 115160 692580 115400 692820
rect 115490 692580 115730 692820
rect 115820 692580 116060 692820
rect 116170 692580 116410 692820
rect 116500 692580 116740 692820
rect 116830 692580 117070 692820
rect 117160 692580 117400 692820
rect 117510 692580 117750 692820
rect 117840 692580 118080 692820
rect 118170 692580 118410 692820
rect 118500 692580 118740 692820
rect 118850 692580 119090 692820
rect 119180 692580 119420 692820
rect 119510 692580 119750 692820
rect 119840 692580 120080 692820
rect 120190 692580 120430 692820
rect 120520 692580 120760 692820
rect 120850 692580 121090 692820
rect 121180 692580 121420 692820
rect 121530 692580 121770 692820
rect 110810 692250 111050 692490
rect 111140 692250 111380 692490
rect 111470 692250 111710 692490
rect 111800 692250 112040 692490
rect 112150 692250 112390 692490
rect 112480 692250 112720 692490
rect 112810 692250 113050 692490
rect 113140 692250 113380 692490
rect 113490 692250 113730 692490
rect 113820 692250 114060 692490
rect 114150 692250 114390 692490
rect 114480 692250 114720 692490
rect 114830 692250 115070 692490
rect 115160 692250 115400 692490
rect 115490 692250 115730 692490
rect 115820 692250 116060 692490
rect 116170 692250 116410 692490
rect 116500 692250 116740 692490
rect 116830 692250 117070 692490
rect 117160 692250 117400 692490
rect 117510 692250 117750 692490
rect 117840 692250 118080 692490
rect 118170 692250 118410 692490
rect 118500 692250 118740 692490
rect 118850 692250 119090 692490
rect 119180 692250 119420 692490
rect 119510 692250 119750 692490
rect 119840 692250 120080 692490
rect 120190 692250 120430 692490
rect 120520 692250 120760 692490
rect 120850 692250 121090 692490
rect 121180 692250 121420 692490
rect 121530 692250 121770 692490
rect 110810 691920 111050 692160
rect 111140 691920 111380 692160
rect 111470 691920 111710 692160
rect 111800 691920 112040 692160
rect 112150 691920 112390 692160
rect 112480 691920 112720 692160
rect 112810 691920 113050 692160
rect 113140 691920 113380 692160
rect 113490 691920 113730 692160
rect 113820 691920 114060 692160
rect 114150 691920 114390 692160
rect 114480 691920 114720 692160
rect 114830 691920 115070 692160
rect 115160 691920 115400 692160
rect 115490 691920 115730 692160
rect 115820 691920 116060 692160
rect 116170 691920 116410 692160
rect 116500 691920 116740 692160
rect 116830 691920 117070 692160
rect 117160 691920 117400 692160
rect 117510 691920 117750 692160
rect 117840 691920 118080 692160
rect 118170 691920 118410 692160
rect 118500 691920 118740 692160
rect 118850 691920 119090 692160
rect 119180 691920 119420 692160
rect 119510 691920 119750 692160
rect 119840 691920 120080 692160
rect 120190 691920 120430 692160
rect 120520 691920 120760 692160
rect 120850 691920 121090 692160
rect 121180 691920 121420 692160
rect 121530 691920 121770 692160
rect 110810 691570 111050 691810
rect 111140 691570 111380 691810
rect 111470 691570 111710 691810
rect 111800 691570 112040 691810
rect 112150 691570 112390 691810
rect 112480 691570 112720 691810
rect 112810 691570 113050 691810
rect 113140 691570 113380 691810
rect 113490 691570 113730 691810
rect 113820 691570 114060 691810
rect 114150 691570 114390 691810
rect 114480 691570 114720 691810
rect 114830 691570 115070 691810
rect 115160 691570 115400 691810
rect 115490 691570 115730 691810
rect 115820 691570 116060 691810
rect 116170 691570 116410 691810
rect 116500 691570 116740 691810
rect 116830 691570 117070 691810
rect 117160 691570 117400 691810
rect 117510 691570 117750 691810
rect 117840 691570 118080 691810
rect 118170 691570 118410 691810
rect 118500 691570 118740 691810
rect 118850 691570 119090 691810
rect 119180 691570 119420 691810
rect 119510 691570 119750 691810
rect 119840 691570 120080 691810
rect 120190 691570 120430 691810
rect 120520 691570 120760 691810
rect 120850 691570 121090 691810
rect 121180 691570 121420 691810
rect 121530 691570 121770 691810
rect 110810 691240 111050 691480
rect 111140 691240 111380 691480
rect 111470 691240 111710 691480
rect 111800 691240 112040 691480
rect 112150 691240 112390 691480
rect 112480 691240 112720 691480
rect 112810 691240 113050 691480
rect 113140 691240 113380 691480
rect 113490 691240 113730 691480
rect 113820 691240 114060 691480
rect 114150 691240 114390 691480
rect 114480 691240 114720 691480
rect 114830 691240 115070 691480
rect 115160 691240 115400 691480
rect 115490 691240 115730 691480
rect 115820 691240 116060 691480
rect 116170 691240 116410 691480
rect 116500 691240 116740 691480
rect 116830 691240 117070 691480
rect 117160 691240 117400 691480
rect 117510 691240 117750 691480
rect 117840 691240 118080 691480
rect 118170 691240 118410 691480
rect 118500 691240 118740 691480
rect 118850 691240 119090 691480
rect 119180 691240 119420 691480
rect 119510 691240 119750 691480
rect 119840 691240 120080 691480
rect 120190 691240 120430 691480
rect 120520 691240 120760 691480
rect 120850 691240 121090 691480
rect 121180 691240 121420 691480
rect 121530 691240 121770 691480
rect 110810 690910 111050 691150
rect 111140 690910 111380 691150
rect 111470 690910 111710 691150
rect 111800 690910 112040 691150
rect 112150 690910 112390 691150
rect 112480 690910 112720 691150
rect 112810 690910 113050 691150
rect 113140 690910 113380 691150
rect 113490 690910 113730 691150
rect 113820 690910 114060 691150
rect 114150 690910 114390 691150
rect 114480 690910 114720 691150
rect 114830 690910 115070 691150
rect 115160 690910 115400 691150
rect 115490 690910 115730 691150
rect 115820 690910 116060 691150
rect 116170 690910 116410 691150
rect 116500 690910 116740 691150
rect 116830 690910 117070 691150
rect 117160 690910 117400 691150
rect 117510 690910 117750 691150
rect 117840 690910 118080 691150
rect 118170 690910 118410 691150
rect 118500 690910 118740 691150
rect 118850 690910 119090 691150
rect 119180 690910 119420 691150
rect 119510 690910 119750 691150
rect 119840 690910 120080 691150
rect 120190 690910 120430 691150
rect 120520 690910 120760 691150
rect 120850 690910 121090 691150
rect 121180 690910 121420 691150
rect 121530 690910 121770 691150
rect 110810 690580 111050 690820
rect 111140 690580 111380 690820
rect 111470 690580 111710 690820
rect 111800 690580 112040 690820
rect 112150 690580 112390 690820
rect 112480 690580 112720 690820
rect 112810 690580 113050 690820
rect 113140 690580 113380 690820
rect 113490 690580 113730 690820
rect 113820 690580 114060 690820
rect 114150 690580 114390 690820
rect 114480 690580 114720 690820
rect 114830 690580 115070 690820
rect 115160 690580 115400 690820
rect 115490 690580 115730 690820
rect 115820 690580 116060 690820
rect 116170 690580 116410 690820
rect 116500 690580 116740 690820
rect 116830 690580 117070 690820
rect 117160 690580 117400 690820
rect 117510 690580 117750 690820
rect 117840 690580 118080 690820
rect 118170 690580 118410 690820
rect 118500 690580 118740 690820
rect 118850 690580 119090 690820
rect 119180 690580 119420 690820
rect 119510 690580 119750 690820
rect 119840 690580 120080 690820
rect 120190 690580 120430 690820
rect 120520 690580 120760 690820
rect 120850 690580 121090 690820
rect 121180 690580 121420 690820
rect 121530 690580 121770 690820
rect 110810 690230 111050 690470
rect 111140 690230 111380 690470
rect 111470 690230 111710 690470
rect 111800 690230 112040 690470
rect 112150 690230 112390 690470
rect 112480 690230 112720 690470
rect 112810 690230 113050 690470
rect 113140 690230 113380 690470
rect 113490 690230 113730 690470
rect 113820 690230 114060 690470
rect 114150 690230 114390 690470
rect 114480 690230 114720 690470
rect 114830 690230 115070 690470
rect 115160 690230 115400 690470
rect 115490 690230 115730 690470
rect 115820 690230 116060 690470
rect 116170 690230 116410 690470
rect 116500 690230 116740 690470
rect 116830 690230 117070 690470
rect 117160 690230 117400 690470
rect 117510 690230 117750 690470
rect 117840 690230 118080 690470
rect 118170 690230 118410 690470
rect 118500 690230 118740 690470
rect 118850 690230 119090 690470
rect 119180 690230 119420 690470
rect 119510 690230 119750 690470
rect 119840 690230 120080 690470
rect 120190 690230 120430 690470
rect 120520 690230 120760 690470
rect 120850 690230 121090 690470
rect 121180 690230 121420 690470
rect 121530 690230 121770 690470
rect 110810 689900 111050 690140
rect 111140 689900 111380 690140
rect 111470 689900 111710 690140
rect 111800 689900 112040 690140
rect 112150 689900 112390 690140
rect 112480 689900 112720 690140
rect 112810 689900 113050 690140
rect 113140 689900 113380 690140
rect 113490 689900 113730 690140
rect 113820 689900 114060 690140
rect 114150 689900 114390 690140
rect 114480 689900 114720 690140
rect 114830 689900 115070 690140
rect 115160 689900 115400 690140
rect 115490 689900 115730 690140
rect 115820 689900 116060 690140
rect 116170 689900 116410 690140
rect 116500 689900 116740 690140
rect 116830 689900 117070 690140
rect 117160 689900 117400 690140
rect 117510 689900 117750 690140
rect 117840 689900 118080 690140
rect 118170 689900 118410 690140
rect 118500 689900 118740 690140
rect 118850 689900 119090 690140
rect 119180 689900 119420 690140
rect 119510 689900 119750 690140
rect 119840 689900 120080 690140
rect 120190 689900 120430 690140
rect 120520 689900 120760 690140
rect 120850 689900 121090 690140
rect 121180 689900 121420 690140
rect 121530 689900 121770 690140
rect 110810 689570 111050 689810
rect 111140 689570 111380 689810
rect 111470 689570 111710 689810
rect 111800 689570 112040 689810
rect 112150 689570 112390 689810
rect 112480 689570 112720 689810
rect 112810 689570 113050 689810
rect 113140 689570 113380 689810
rect 113490 689570 113730 689810
rect 113820 689570 114060 689810
rect 114150 689570 114390 689810
rect 114480 689570 114720 689810
rect 114830 689570 115070 689810
rect 115160 689570 115400 689810
rect 115490 689570 115730 689810
rect 115820 689570 116060 689810
rect 116170 689570 116410 689810
rect 116500 689570 116740 689810
rect 116830 689570 117070 689810
rect 117160 689570 117400 689810
rect 117510 689570 117750 689810
rect 117840 689570 118080 689810
rect 118170 689570 118410 689810
rect 118500 689570 118740 689810
rect 118850 689570 119090 689810
rect 119180 689570 119420 689810
rect 119510 689570 119750 689810
rect 119840 689570 120080 689810
rect 120190 689570 120430 689810
rect 120520 689570 120760 689810
rect 120850 689570 121090 689810
rect 121180 689570 121420 689810
rect 121530 689570 121770 689810
rect 110810 689240 111050 689480
rect 111140 689240 111380 689480
rect 111470 689240 111710 689480
rect 111800 689240 112040 689480
rect 112150 689240 112390 689480
rect 112480 689240 112720 689480
rect 112810 689240 113050 689480
rect 113140 689240 113380 689480
rect 113490 689240 113730 689480
rect 113820 689240 114060 689480
rect 114150 689240 114390 689480
rect 114480 689240 114720 689480
rect 114830 689240 115070 689480
rect 115160 689240 115400 689480
rect 115490 689240 115730 689480
rect 115820 689240 116060 689480
rect 116170 689240 116410 689480
rect 116500 689240 116740 689480
rect 116830 689240 117070 689480
rect 117160 689240 117400 689480
rect 117510 689240 117750 689480
rect 117840 689240 118080 689480
rect 118170 689240 118410 689480
rect 118500 689240 118740 689480
rect 118850 689240 119090 689480
rect 119180 689240 119420 689480
rect 119510 689240 119750 689480
rect 119840 689240 120080 689480
rect 120190 689240 120430 689480
rect 120520 689240 120760 689480
rect 120850 689240 121090 689480
rect 121180 689240 121420 689480
rect 121530 689240 121770 689480
rect 110810 688890 111050 689130
rect 111140 688890 111380 689130
rect 111470 688890 111710 689130
rect 111800 688890 112040 689130
rect 112150 688890 112390 689130
rect 112480 688890 112720 689130
rect 112810 688890 113050 689130
rect 113140 688890 113380 689130
rect 113490 688890 113730 689130
rect 113820 688890 114060 689130
rect 114150 688890 114390 689130
rect 114480 688890 114720 689130
rect 114830 688890 115070 689130
rect 115160 688890 115400 689130
rect 115490 688890 115730 689130
rect 115820 688890 116060 689130
rect 116170 688890 116410 689130
rect 116500 688890 116740 689130
rect 116830 688890 117070 689130
rect 117160 688890 117400 689130
rect 117510 688890 117750 689130
rect 117840 688890 118080 689130
rect 118170 688890 118410 689130
rect 118500 688890 118740 689130
rect 118850 688890 119090 689130
rect 119180 688890 119420 689130
rect 119510 688890 119750 689130
rect 119840 688890 120080 689130
rect 120190 688890 120430 689130
rect 120520 688890 120760 689130
rect 120850 688890 121090 689130
rect 121180 688890 121420 689130
rect 121530 688890 121770 689130
rect 110810 688560 111050 688800
rect 111140 688560 111380 688800
rect 111470 688560 111710 688800
rect 111800 688560 112040 688800
rect 112150 688560 112390 688800
rect 112480 688560 112720 688800
rect 112810 688560 113050 688800
rect 113140 688560 113380 688800
rect 113490 688560 113730 688800
rect 113820 688560 114060 688800
rect 114150 688560 114390 688800
rect 114480 688560 114720 688800
rect 114830 688560 115070 688800
rect 115160 688560 115400 688800
rect 115490 688560 115730 688800
rect 115820 688560 116060 688800
rect 116170 688560 116410 688800
rect 116500 688560 116740 688800
rect 116830 688560 117070 688800
rect 117160 688560 117400 688800
rect 117510 688560 117750 688800
rect 117840 688560 118080 688800
rect 118170 688560 118410 688800
rect 118500 688560 118740 688800
rect 118850 688560 119090 688800
rect 119180 688560 119420 688800
rect 119510 688560 119750 688800
rect 119840 688560 120080 688800
rect 120190 688560 120430 688800
rect 120520 688560 120760 688800
rect 120850 688560 121090 688800
rect 121180 688560 121420 688800
rect 121530 688560 121770 688800
rect 110810 688230 111050 688470
rect 111140 688230 111380 688470
rect 111470 688230 111710 688470
rect 111800 688230 112040 688470
rect 112150 688230 112390 688470
rect 112480 688230 112720 688470
rect 112810 688230 113050 688470
rect 113140 688230 113380 688470
rect 113490 688230 113730 688470
rect 113820 688230 114060 688470
rect 114150 688230 114390 688470
rect 114480 688230 114720 688470
rect 114830 688230 115070 688470
rect 115160 688230 115400 688470
rect 115490 688230 115730 688470
rect 115820 688230 116060 688470
rect 116170 688230 116410 688470
rect 116500 688230 116740 688470
rect 116830 688230 117070 688470
rect 117160 688230 117400 688470
rect 117510 688230 117750 688470
rect 117840 688230 118080 688470
rect 118170 688230 118410 688470
rect 118500 688230 118740 688470
rect 118850 688230 119090 688470
rect 119180 688230 119420 688470
rect 119510 688230 119750 688470
rect 119840 688230 120080 688470
rect 120190 688230 120430 688470
rect 120520 688230 120760 688470
rect 120850 688230 121090 688470
rect 121180 688230 121420 688470
rect 121530 688230 121770 688470
rect 110810 687900 111050 688140
rect 111140 687900 111380 688140
rect 111470 687900 111710 688140
rect 111800 687900 112040 688140
rect 112150 687900 112390 688140
rect 112480 687900 112720 688140
rect 112810 687900 113050 688140
rect 113140 687900 113380 688140
rect 113490 687900 113730 688140
rect 113820 687900 114060 688140
rect 114150 687900 114390 688140
rect 114480 687900 114720 688140
rect 114830 687900 115070 688140
rect 115160 687900 115400 688140
rect 115490 687900 115730 688140
rect 115820 687900 116060 688140
rect 116170 687900 116410 688140
rect 116500 687900 116740 688140
rect 116830 687900 117070 688140
rect 117160 687900 117400 688140
rect 117510 687900 117750 688140
rect 117840 687900 118080 688140
rect 118170 687900 118410 688140
rect 118500 687900 118740 688140
rect 118850 687900 119090 688140
rect 119180 687900 119420 688140
rect 119510 687900 119750 688140
rect 119840 687900 120080 688140
rect 120190 687900 120430 688140
rect 120520 687900 120760 688140
rect 120850 687900 121090 688140
rect 121180 687900 121420 688140
rect 121530 687900 121770 688140
rect 110810 687550 111050 687790
rect 111140 687550 111380 687790
rect 111470 687550 111710 687790
rect 111800 687550 112040 687790
rect 112150 687550 112390 687790
rect 112480 687550 112720 687790
rect 112810 687550 113050 687790
rect 113140 687550 113380 687790
rect 113490 687550 113730 687790
rect 113820 687550 114060 687790
rect 114150 687550 114390 687790
rect 114480 687550 114720 687790
rect 114830 687550 115070 687790
rect 115160 687550 115400 687790
rect 115490 687550 115730 687790
rect 115820 687550 116060 687790
rect 116170 687550 116410 687790
rect 116500 687550 116740 687790
rect 116830 687550 117070 687790
rect 117160 687550 117400 687790
rect 117510 687550 117750 687790
rect 117840 687550 118080 687790
rect 118170 687550 118410 687790
rect 118500 687550 118740 687790
rect 118850 687550 119090 687790
rect 119180 687550 119420 687790
rect 119510 687550 119750 687790
rect 119840 687550 120080 687790
rect 120190 687550 120430 687790
rect 120520 687550 120760 687790
rect 120850 687550 121090 687790
rect 121180 687550 121420 687790
rect 121530 687550 121770 687790
rect 110810 687220 111050 687460
rect 111140 687220 111380 687460
rect 111470 687220 111710 687460
rect 111800 687220 112040 687460
rect 112150 687220 112390 687460
rect 112480 687220 112720 687460
rect 112810 687220 113050 687460
rect 113140 687220 113380 687460
rect 113490 687220 113730 687460
rect 113820 687220 114060 687460
rect 114150 687220 114390 687460
rect 114480 687220 114720 687460
rect 114830 687220 115070 687460
rect 115160 687220 115400 687460
rect 115490 687220 115730 687460
rect 115820 687220 116060 687460
rect 116170 687220 116410 687460
rect 116500 687220 116740 687460
rect 116830 687220 117070 687460
rect 117160 687220 117400 687460
rect 117510 687220 117750 687460
rect 117840 687220 118080 687460
rect 118170 687220 118410 687460
rect 118500 687220 118740 687460
rect 118850 687220 119090 687460
rect 119180 687220 119420 687460
rect 119510 687220 119750 687460
rect 119840 687220 120080 687460
rect 120190 687220 120430 687460
rect 120520 687220 120760 687460
rect 120850 687220 121090 687460
rect 121180 687220 121420 687460
rect 121530 687220 121770 687460
rect 110810 686890 111050 687130
rect 111140 686890 111380 687130
rect 111470 686890 111710 687130
rect 111800 686890 112040 687130
rect 112150 686890 112390 687130
rect 112480 686890 112720 687130
rect 112810 686890 113050 687130
rect 113140 686890 113380 687130
rect 113490 686890 113730 687130
rect 113820 686890 114060 687130
rect 114150 686890 114390 687130
rect 114480 686890 114720 687130
rect 114830 686890 115070 687130
rect 115160 686890 115400 687130
rect 115490 686890 115730 687130
rect 115820 686890 116060 687130
rect 116170 686890 116410 687130
rect 116500 686890 116740 687130
rect 116830 686890 117070 687130
rect 117160 686890 117400 687130
rect 117510 686890 117750 687130
rect 117840 686890 118080 687130
rect 118170 686890 118410 687130
rect 118500 686890 118740 687130
rect 118850 686890 119090 687130
rect 119180 686890 119420 687130
rect 119510 686890 119750 687130
rect 119840 686890 120080 687130
rect 120190 686890 120430 687130
rect 120520 686890 120760 687130
rect 120850 686890 121090 687130
rect 121180 686890 121420 687130
rect 121530 686890 121770 687130
rect 110810 686560 111050 686800
rect 111140 686560 111380 686800
rect 111470 686560 111710 686800
rect 111800 686560 112040 686800
rect 112150 686560 112390 686800
rect 112480 686560 112720 686800
rect 112810 686560 113050 686800
rect 113140 686560 113380 686800
rect 113490 686560 113730 686800
rect 113820 686560 114060 686800
rect 114150 686560 114390 686800
rect 114480 686560 114720 686800
rect 114830 686560 115070 686800
rect 115160 686560 115400 686800
rect 115490 686560 115730 686800
rect 115820 686560 116060 686800
rect 116170 686560 116410 686800
rect 116500 686560 116740 686800
rect 116830 686560 117070 686800
rect 117160 686560 117400 686800
rect 117510 686560 117750 686800
rect 117840 686560 118080 686800
rect 118170 686560 118410 686800
rect 118500 686560 118740 686800
rect 118850 686560 119090 686800
rect 119180 686560 119420 686800
rect 119510 686560 119750 686800
rect 119840 686560 120080 686800
rect 120190 686560 120430 686800
rect 120520 686560 120760 686800
rect 120850 686560 121090 686800
rect 121180 686560 121420 686800
rect 121530 686560 121770 686800
rect 110810 686210 111050 686450
rect 111140 686210 111380 686450
rect 111470 686210 111710 686450
rect 111800 686210 112040 686450
rect 112150 686210 112390 686450
rect 112480 686210 112720 686450
rect 112810 686210 113050 686450
rect 113140 686210 113380 686450
rect 113490 686210 113730 686450
rect 113820 686210 114060 686450
rect 114150 686210 114390 686450
rect 114480 686210 114720 686450
rect 114830 686210 115070 686450
rect 115160 686210 115400 686450
rect 115490 686210 115730 686450
rect 115820 686210 116060 686450
rect 116170 686210 116410 686450
rect 116500 686210 116740 686450
rect 116830 686210 117070 686450
rect 117160 686210 117400 686450
rect 117510 686210 117750 686450
rect 117840 686210 118080 686450
rect 118170 686210 118410 686450
rect 118500 686210 118740 686450
rect 118850 686210 119090 686450
rect 119180 686210 119420 686450
rect 119510 686210 119750 686450
rect 119840 686210 120080 686450
rect 120190 686210 120430 686450
rect 120520 686210 120760 686450
rect 120850 686210 121090 686450
rect 121180 686210 121420 686450
rect 121530 686210 121770 686450
rect 110810 685880 111050 686120
rect 111140 685880 111380 686120
rect 111470 685880 111710 686120
rect 111800 685880 112040 686120
rect 112150 685880 112390 686120
rect 112480 685880 112720 686120
rect 112810 685880 113050 686120
rect 113140 685880 113380 686120
rect 113490 685880 113730 686120
rect 113820 685880 114060 686120
rect 114150 685880 114390 686120
rect 114480 685880 114720 686120
rect 114830 685880 115070 686120
rect 115160 685880 115400 686120
rect 115490 685880 115730 686120
rect 115820 685880 116060 686120
rect 116170 685880 116410 686120
rect 116500 685880 116740 686120
rect 116830 685880 117070 686120
rect 117160 685880 117400 686120
rect 117510 685880 117750 686120
rect 117840 685880 118080 686120
rect 118170 685880 118410 686120
rect 118500 685880 118740 686120
rect 118850 685880 119090 686120
rect 119180 685880 119420 686120
rect 119510 685880 119750 686120
rect 119840 685880 120080 686120
rect 120190 685880 120430 686120
rect 120520 685880 120760 686120
rect 120850 685880 121090 686120
rect 121180 685880 121420 686120
rect 121530 685880 121770 686120
rect 110810 685550 111050 685790
rect 111140 685550 111380 685790
rect 111470 685550 111710 685790
rect 111800 685550 112040 685790
rect 112150 685550 112390 685790
rect 112480 685550 112720 685790
rect 112810 685550 113050 685790
rect 113140 685550 113380 685790
rect 113490 685550 113730 685790
rect 113820 685550 114060 685790
rect 114150 685550 114390 685790
rect 114480 685550 114720 685790
rect 114830 685550 115070 685790
rect 115160 685550 115400 685790
rect 115490 685550 115730 685790
rect 115820 685550 116060 685790
rect 116170 685550 116410 685790
rect 116500 685550 116740 685790
rect 116830 685550 117070 685790
rect 117160 685550 117400 685790
rect 117510 685550 117750 685790
rect 117840 685550 118080 685790
rect 118170 685550 118410 685790
rect 118500 685550 118740 685790
rect 118850 685550 119090 685790
rect 119180 685550 119420 685790
rect 119510 685550 119750 685790
rect 119840 685550 120080 685790
rect 120190 685550 120430 685790
rect 120520 685550 120760 685790
rect 120850 685550 121090 685790
rect 121180 685550 121420 685790
rect 121530 685550 121770 685790
rect 110810 685220 111050 685460
rect 111140 685220 111380 685460
rect 111470 685220 111710 685460
rect 111800 685220 112040 685460
rect 112150 685220 112390 685460
rect 112480 685220 112720 685460
rect 112810 685220 113050 685460
rect 113140 685220 113380 685460
rect 113490 685220 113730 685460
rect 113820 685220 114060 685460
rect 114150 685220 114390 685460
rect 114480 685220 114720 685460
rect 114830 685220 115070 685460
rect 115160 685220 115400 685460
rect 115490 685220 115730 685460
rect 115820 685220 116060 685460
rect 116170 685220 116410 685460
rect 116500 685220 116740 685460
rect 116830 685220 117070 685460
rect 117160 685220 117400 685460
rect 117510 685220 117750 685460
rect 117840 685220 118080 685460
rect 118170 685220 118410 685460
rect 118500 685220 118740 685460
rect 118850 685220 119090 685460
rect 119180 685220 119420 685460
rect 119510 685220 119750 685460
rect 119840 685220 120080 685460
rect 120190 685220 120430 685460
rect 120520 685220 120760 685460
rect 120850 685220 121090 685460
rect 121180 685220 121420 685460
rect 121530 685220 121770 685460
rect 110810 684870 111050 685110
rect 111140 684870 111380 685110
rect 111470 684870 111710 685110
rect 111800 684870 112040 685110
rect 112150 684870 112390 685110
rect 112480 684870 112720 685110
rect 112810 684870 113050 685110
rect 113140 684870 113380 685110
rect 113490 684870 113730 685110
rect 113820 684870 114060 685110
rect 114150 684870 114390 685110
rect 114480 684870 114720 685110
rect 114830 684870 115070 685110
rect 115160 684870 115400 685110
rect 115490 684870 115730 685110
rect 115820 684870 116060 685110
rect 116170 684870 116410 685110
rect 116500 684870 116740 685110
rect 116830 684870 117070 685110
rect 117160 684870 117400 685110
rect 117510 684870 117750 685110
rect 117840 684870 118080 685110
rect 118170 684870 118410 685110
rect 118500 684870 118740 685110
rect 118850 684870 119090 685110
rect 119180 684870 119420 685110
rect 119510 684870 119750 685110
rect 119840 684870 120080 685110
rect 120190 684870 120430 685110
rect 120520 684870 120760 685110
rect 120850 684870 121090 685110
rect 121180 684870 121420 685110
rect 121530 684870 121770 685110
rect 110810 684540 111050 684780
rect 111140 684540 111380 684780
rect 111470 684540 111710 684780
rect 111800 684540 112040 684780
rect 112150 684540 112390 684780
rect 112480 684540 112720 684780
rect 112810 684540 113050 684780
rect 113140 684540 113380 684780
rect 113490 684540 113730 684780
rect 113820 684540 114060 684780
rect 114150 684540 114390 684780
rect 114480 684540 114720 684780
rect 114830 684540 115070 684780
rect 115160 684540 115400 684780
rect 115490 684540 115730 684780
rect 115820 684540 116060 684780
rect 116170 684540 116410 684780
rect 116500 684540 116740 684780
rect 116830 684540 117070 684780
rect 117160 684540 117400 684780
rect 117510 684540 117750 684780
rect 117840 684540 118080 684780
rect 118170 684540 118410 684780
rect 118500 684540 118740 684780
rect 118850 684540 119090 684780
rect 119180 684540 119420 684780
rect 119510 684540 119750 684780
rect 119840 684540 120080 684780
rect 120190 684540 120430 684780
rect 120520 684540 120760 684780
rect 120850 684540 121090 684780
rect 121180 684540 121420 684780
rect 121530 684540 121770 684780
rect 110810 684210 111050 684450
rect 111140 684210 111380 684450
rect 111470 684210 111710 684450
rect 111800 684210 112040 684450
rect 112150 684210 112390 684450
rect 112480 684210 112720 684450
rect 112810 684210 113050 684450
rect 113140 684210 113380 684450
rect 113490 684210 113730 684450
rect 113820 684210 114060 684450
rect 114150 684210 114390 684450
rect 114480 684210 114720 684450
rect 114830 684210 115070 684450
rect 115160 684210 115400 684450
rect 115490 684210 115730 684450
rect 115820 684210 116060 684450
rect 116170 684210 116410 684450
rect 116500 684210 116740 684450
rect 116830 684210 117070 684450
rect 117160 684210 117400 684450
rect 117510 684210 117750 684450
rect 117840 684210 118080 684450
rect 118170 684210 118410 684450
rect 118500 684210 118740 684450
rect 118850 684210 119090 684450
rect 119180 684210 119420 684450
rect 119510 684210 119750 684450
rect 119840 684210 120080 684450
rect 120190 684210 120430 684450
rect 120520 684210 120760 684450
rect 120850 684210 121090 684450
rect 121180 684210 121420 684450
rect 121530 684210 121770 684450
rect 110810 683880 111050 684120
rect 111140 683880 111380 684120
rect 111470 683880 111710 684120
rect 111800 683880 112040 684120
rect 112150 683880 112390 684120
rect 112480 683880 112720 684120
rect 112810 683880 113050 684120
rect 113140 683880 113380 684120
rect 113490 683880 113730 684120
rect 113820 683880 114060 684120
rect 114150 683880 114390 684120
rect 114480 683880 114720 684120
rect 114830 683880 115070 684120
rect 115160 683880 115400 684120
rect 115490 683880 115730 684120
rect 115820 683880 116060 684120
rect 116170 683880 116410 684120
rect 116500 683880 116740 684120
rect 116830 683880 117070 684120
rect 117160 683880 117400 684120
rect 117510 683880 117750 684120
rect 117840 683880 118080 684120
rect 118170 683880 118410 684120
rect 118500 683880 118740 684120
rect 118850 683880 119090 684120
rect 119180 683880 119420 684120
rect 119510 683880 119750 684120
rect 119840 683880 120080 684120
rect 120190 683880 120430 684120
rect 120520 683880 120760 684120
rect 120850 683880 121090 684120
rect 121180 683880 121420 684120
rect 121530 683880 121770 684120
rect 122190 694600 122430 694840
rect 122520 694600 122760 694840
rect 122850 694600 123090 694840
rect 123180 694600 123420 694840
rect 123530 694600 123770 694840
rect 123860 694600 124100 694840
rect 124190 694600 124430 694840
rect 124520 694600 124760 694840
rect 124870 694600 125110 694840
rect 125200 694600 125440 694840
rect 125530 694600 125770 694840
rect 125860 694600 126100 694840
rect 126210 694600 126450 694840
rect 126540 694600 126780 694840
rect 126870 694600 127110 694840
rect 127200 694600 127440 694840
rect 127550 694600 127790 694840
rect 127880 694600 128120 694840
rect 128210 694600 128450 694840
rect 128540 694600 128780 694840
rect 128890 694600 129130 694840
rect 129220 694600 129460 694840
rect 129550 694600 129790 694840
rect 129880 694600 130120 694840
rect 130230 694600 130470 694840
rect 130560 694600 130800 694840
rect 130890 694600 131130 694840
rect 131220 694600 131460 694840
rect 131570 694600 131810 694840
rect 131900 694600 132140 694840
rect 132230 694600 132470 694840
rect 132560 694600 132800 694840
rect 132910 694600 133150 694840
rect 122190 694250 122430 694490
rect 122520 694250 122760 694490
rect 122850 694250 123090 694490
rect 123180 694250 123420 694490
rect 123530 694250 123770 694490
rect 123860 694250 124100 694490
rect 124190 694250 124430 694490
rect 124520 694250 124760 694490
rect 124870 694250 125110 694490
rect 125200 694250 125440 694490
rect 125530 694250 125770 694490
rect 125860 694250 126100 694490
rect 126210 694250 126450 694490
rect 126540 694250 126780 694490
rect 126870 694250 127110 694490
rect 127200 694250 127440 694490
rect 127550 694250 127790 694490
rect 127880 694250 128120 694490
rect 128210 694250 128450 694490
rect 128540 694250 128780 694490
rect 128890 694250 129130 694490
rect 129220 694250 129460 694490
rect 129550 694250 129790 694490
rect 129880 694250 130120 694490
rect 130230 694250 130470 694490
rect 130560 694250 130800 694490
rect 130890 694250 131130 694490
rect 131220 694250 131460 694490
rect 131570 694250 131810 694490
rect 131900 694250 132140 694490
rect 132230 694250 132470 694490
rect 132560 694250 132800 694490
rect 132910 694250 133150 694490
rect 122190 693920 122430 694160
rect 122520 693920 122760 694160
rect 122850 693920 123090 694160
rect 123180 693920 123420 694160
rect 123530 693920 123770 694160
rect 123860 693920 124100 694160
rect 124190 693920 124430 694160
rect 124520 693920 124760 694160
rect 124870 693920 125110 694160
rect 125200 693920 125440 694160
rect 125530 693920 125770 694160
rect 125860 693920 126100 694160
rect 126210 693920 126450 694160
rect 126540 693920 126780 694160
rect 126870 693920 127110 694160
rect 127200 693920 127440 694160
rect 127550 693920 127790 694160
rect 127880 693920 128120 694160
rect 128210 693920 128450 694160
rect 128540 693920 128780 694160
rect 128890 693920 129130 694160
rect 129220 693920 129460 694160
rect 129550 693920 129790 694160
rect 129880 693920 130120 694160
rect 130230 693920 130470 694160
rect 130560 693920 130800 694160
rect 130890 693920 131130 694160
rect 131220 693920 131460 694160
rect 131570 693920 131810 694160
rect 131900 693920 132140 694160
rect 132230 693920 132470 694160
rect 132560 693920 132800 694160
rect 132910 693920 133150 694160
rect 122190 693590 122430 693830
rect 122520 693590 122760 693830
rect 122850 693590 123090 693830
rect 123180 693590 123420 693830
rect 123530 693590 123770 693830
rect 123860 693590 124100 693830
rect 124190 693590 124430 693830
rect 124520 693590 124760 693830
rect 124870 693590 125110 693830
rect 125200 693590 125440 693830
rect 125530 693590 125770 693830
rect 125860 693590 126100 693830
rect 126210 693590 126450 693830
rect 126540 693590 126780 693830
rect 126870 693590 127110 693830
rect 127200 693590 127440 693830
rect 127550 693590 127790 693830
rect 127880 693590 128120 693830
rect 128210 693590 128450 693830
rect 128540 693590 128780 693830
rect 128890 693590 129130 693830
rect 129220 693590 129460 693830
rect 129550 693590 129790 693830
rect 129880 693590 130120 693830
rect 130230 693590 130470 693830
rect 130560 693590 130800 693830
rect 130890 693590 131130 693830
rect 131220 693590 131460 693830
rect 131570 693590 131810 693830
rect 131900 693590 132140 693830
rect 132230 693590 132470 693830
rect 132560 693590 132800 693830
rect 132910 693590 133150 693830
rect 122190 693260 122430 693500
rect 122520 693260 122760 693500
rect 122850 693260 123090 693500
rect 123180 693260 123420 693500
rect 123530 693260 123770 693500
rect 123860 693260 124100 693500
rect 124190 693260 124430 693500
rect 124520 693260 124760 693500
rect 124870 693260 125110 693500
rect 125200 693260 125440 693500
rect 125530 693260 125770 693500
rect 125860 693260 126100 693500
rect 126210 693260 126450 693500
rect 126540 693260 126780 693500
rect 126870 693260 127110 693500
rect 127200 693260 127440 693500
rect 127550 693260 127790 693500
rect 127880 693260 128120 693500
rect 128210 693260 128450 693500
rect 128540 693260 128780 693500
rect 128890 693260 129130 693500
rect 129220 693260 129460 693500
rect 129550 693260 129790 693500
rect 129880 693260 130120 693500
rect 130230 693260 130470 693500
rect 130560 693260 130800 693500
rect 130890 693260 131130 693500
rect 131220 693260 131460 693500
rect 131570 693260 131810 693500
rect 131900 693260 132140 693500
rect 132230 693260 132470 693500
rect 132560 693260 132800 693500
rect 132910 693260 133150 693500
rect 122190 692910 122430 693150
rect 122520 692910 122760 693150
rect 122850 692910 123090 693150
rect 123180 692910 123420 693150
rect 123530 692910 123770 693150
rect 123860 692910 124100 693150
rect 124190 692910 124430 693150
rect 124520 692910 124760 693150
rect 124870 692910 125110 693150
rect 125200 692910 125440 693150
rect 125530 692910 125770 693150
rect 125860 692910 126100 693150
rect 126210 692910 126450 693150
rect 126540 692910 126780 693150
rect 126870 692910 127110 693150
rect 127200 692910 127440 693150
rect 127550 692910 127790 693150
rect 127880 692910 128120 693150
rect 128210 692910 128450 693150
rect 128540 692910 128780 693150
rect 128890 692910 129130 693150
rect 129220 692910 129460 693150
rect 129550 692910 129790 693150
rect 129880 692910 130120 693150
rect 130230 692910 130470 693150
rect 130560 692910 130800 693150
rect 130890 692910 131130 693150
rect 131220 692910 131460 693150
rect 131570 692910 131810 693150
rect 131900 692910 132140 693150
rect 132230 692910 132470 693150
rect 132560 692910 132800 693150
rect 132910 692910 133150 693150
rect 122190 692580 122430 692820
rect 122520 692580 122760 692820
rect 122850 692580 123090 692820
rect 123180 692580 123420 692820
rect 123530 692580 123770 692820
rect 123860 692580 124100 692820
rect 124190 692580 124430 692820
rect 124520 692580 124760 692820
rect 124870 692580 125110 692820
rect 125200 692580 125440 692820
rect 125530 692580 125770 692820
rect 125860 692580 126100 692820
rect 126210 692580 126450 692820
rect 126540 692580 126780 692820
rect 126870 692580 127110 692820
rect 127200 692580 127440 692820
rect 127550 692580 127790 692820
rect 127880 692580 128120 692820
rect 128210 692580 128450 692820
rect 128540 692580 128780 692820
rect 128890 692580 129130 692820
rect 129220 692580 129460 692820
rect 129550 692580 129790 692820
rect 129880 692580 130120 692820
rect 130230 692580 130470 692820
rect 130560 692580 130800 692820
rect 130890 692580 131130 692820
rect 131220 692580 131460 692820
rect 131570 692580 131810 692820
rect 131900 692580 132140 692820
rect 132230 692580 132470 692820
rect 132560 692580 132800 692820
rect 132910 692580 133150 692820
rect 122190 692250 122430 692490
rect 122520 692250 122760 692490
rect 122850 692250 123090 692490
rect 123180 692250 123420 692490
rect 123530 692250 123770 692490
rect 123860 692250 124100 692490
rect 124190 692250 124430 692490
rect 124520 692250 124760 692490
rect 124870 692250 125110 692490
rect 125200 692250 125440 692490
rect 125530 692250 125770 692490
rect 125860 692250 126100 692490
rect 126210 692250 126450 692490
rect 126540 692250 126780 692490
rect 126870 692250 127110 692490
rect 127200 692250 127440 692490
rect 127550 692250 127790 692490
rect 127880 692250 128120 692490
rect 128210 692250 128450 692490
rect 128540 692250 128780 692490
rect 128890 692250 129130 692490
rect 129220 692250 129460 692490
rect 129550 692250 129790 692490
rect 129880 692250 130120 692490
rect 130230 692250 130470 692490
rect 130560 692250 130800 692490
rect 130890 692250 131130 692490
rect 131220 692250 131460 692490
rect 131570 692250 131810 692490
rect 131900 692250 132140 692490
rect 132230 692250 132470 692490
rect 132560 692250 132800 692490
rect 132910 692250 133150 692490
rect 122190 691920 122430 692160
rect 122520 691920 122760 692160
rect 122850 691920 123090 692160
rect 123180 691920 123420 692160
rect 123530 691920 123770 692160
rect 123860 691920 124100 692160
rect 124190 691920 124430 692160
rect 124520 691920 124760 692160
rect 124870 691920 125110 692160
rect 125200 691920 125440 692160
rect 125530 691920 125770 692160
rect 125860 691920 126100 692160
rect 126210 691920 126450 692160
rect 126540 691920 126780 692160
rect 126870 691920 127110 692160
rect 127200 691920 127440 692160
rect 127550 691920 127790 692160
rect 127880 691920 128120 692160
rect 128210 691920 128450 692160
rect 128540 691920 128780 692160
rect 128890 691920 129130 692160
rect 129220 691920 129460 692160
rect 129550 691920 129790 692160
rect 129880 691920 130120 692160
rect 130230 691920 130470 692160
rect 130560 691920 130800 692160
rect 130890 691920 131130 692160
rect 131220 691920 131460 692160
rect 131570 691920 131810 692160
rect 131900 691920 132140 692160
rect 132230 691920 132470 692160
rect 132560 691920 132800 692160
rect 132910 691920 133150 692160
rect 122190 691570 122430 691810
rect 122520 691570 122760 691810
rect 122850 691570 123090 691810
rect 123180 691570 123420 691810
rect 123530 691570 123770 691810
rect 123860 691570 124100 691810
rect 124190 691570 124430 691810
rect 124520 691570 124760 691810
rect 124870 691570 125110 691810
rect 125200 691570 125440 691810
rect 125530 691570 125770 691810
rect 125860 691570 126100 691810
rect 126210 691570 126450 691810
rect 126540 691570 126780 691810
rect 126870 691570 127110 691810
rect 127200 691570 127440 691810
rect 127550 691570 127790 691810
rect 127880 691570 128120 691810
rect 128210 691570 128450 691810
rect 128540 691570 128780 691810
rect 128890 691570 129130 691810
rect 129220 691570 129460 691810
rect 129550 691570 129790 691810
rect 129880 691570 130120 691810
rect 130230 691570 130470 691810
rect 130560 691570 130800 691810
rect 130890 691570 131130 691810
rect 131220 691570 131460 691810
rect 131570 691570 131810 691810
rect 131900 691570 132140 691810
rect 132230 691570 132470 691810
rect 132560 691570 132800 691810
rect 132910 691570 133150 691810
rect 122190 691240 122430 691480
rect 122520 691240 122760 691480
rect 122850 691240 123090 691480
rect 123180 691240 123420 691480
rect 123530 691240 123770 691480
rect 123860 691240 124100 691480
rect 124190 691240 124430 691480
rect 124520 691240 124760 691480
rect 124870 691240 125110 691480
rect 125200 691240 125440 691480
rect 125530 691240 125770 691480
rect 125860 691240 126100 691480
rect 126210 691240 126450 691480
rect 126540 691240 126780 691480
rect 126870 691240 127110 691480
rect 127200 691240 127440 691480
rect 127550 691240 127790 691480
rect 127880 691240 128120 691480
rect 128210 691240 128450 691480
rect 128540 691240 128780 691480
rect 128890 691240 129130 691480
rect 129220 691240 129460 691480
rect 129550 691240 129790 691480
rect 129880 691240 130120 691480
rect 130230 691240 130470 691480
rect 130560 691240 130800 691480
rect 130890 691240 131130 691480
rect 131220 691240 131460 691480
rect 131570 691240 131810 691480
rect 131900 691240 132140 691480
rect 132230 691240 132470 691480
rect 132560 691240 132800 691480
rect 132910 691240 133150 691480
rect 122190 690910 122430 691150
rect 122520 690910 122760 691150
rect 122850 690910 123090 691150
rect 123180 690910 123420 691150
rect 123530 690910 123770 691150
rect 123860 690910 124100 691150
rect 124190 690910 124430 691150
rect 124520 690910 124760 691150
rect 124870 690910 125110 691150
rect 125200 690910 125440 691150
rect 125530 690910 125770 691150
rect 125860 690910 126100 691150
rect 126210 690910 126450 691150
rect 126540 690910 126780 691150
rect 126870 690910 127110 691150
rect 127200 690910 127440 691150
rect 127550 690910 127790 691150
rect 127880 690910 128120 691150
rect 128210 690910 128450 691150
rect 128540 690910 128780 691150
rect 128890 690910 129130 691150
rect 129220 690910 129460 691150
rect 129550 690910 129790 691150
rect 129880 690910 130120 691150
rect 130230 690910 130470 691150
rect 130560 690910 130800 691150
rect 130890 690910 131130 691150
rect 131220 690910 131460 691150
rect 131570 690910 131810 691150
rect 131900 690910 132140 691150
rect 132230 690910 132470 691150
rect 132560 690910 132800 691150
rect 132910 690910 133150 691150
rect 122190 690580 122430 690820
rect 122520 690580 122760 690820
rect 122850 690580 123090 690820
rect 123180 690580 123420 690820
rect 123530 690580 123770 690820
rect 123860 690580 124100 690820
rect 124190 690580 124430 690820
rect 124520 690580 124760 690820
rect 124870 690580 125110 690820
rect 125200 690580 125440 690820
rect 125530 690580 125770 690820
rect 125860 690580 126100 690820
rect 126210 690580 126450 690820
rect 126540 690580 126780 690820
rect 126870 690580 127110 690820
rect 127200 690580 127440 690820
rect 127550 690580 127790 690820
rect 127880 690580 128120 690820
rect 128210 690580 128450 690820
rect 128540 690580 128780 690820
rect 128890 690580 129130 690820
rect 129220 690580 129460 690820
rect 129550 690580 129790 690820
rect 129880 690580 130120 690820
rect 130230 690580 130470 690820
rect 130560 690580 130800 690820
rect 130890 690580 131130 690820
rect 131220 690580 131460 690820
rect 131570 690580 131810 690820
rect 131900 690580 132140 690820
rect 132230 690580 132470 690820
rect 132560 690580 132800 690820
rect 132910 690580 133150 690820
rect 122190 690230 122430 690470
rect 122520 690230 122760 690470
rect 122850 690230 123090 690470
rect 123180 690230 123420 690470
rect 123530 690230 123770 690470
rect 123860 690230 124100 690470
rect 124190 690230 124430 690470
rect 124520 690230 124760 690470
rect 124870 690230 125110 690470
rect 125200 690230 125440 690470
rect 125530 690230 125770 690470
rect 125860 690230 126100 690470
rect 126210 690230 126450 690470
rect 126540 690230 126780 690470
rect 126870 690230 127110 690470
rect 127200 690230 127440 690470
rect 127550 690230 127790 690470
rect 127880 690230 128120 690470
rect 128210 690230 128450 690470
rect 128540 690230 128780 690470
rect 128890 690230 129130 690470
rect 129220 690230 129460 690470
rect 129550 690230 129790 690470
rect 129880 690230 130120 690470
rect 130230 690230 130470 690470
rect 130560 690230 130800 690470
rect 130890 690230 131130 690470
rect 131220 690230 131460 690470
rect 131570 690230 131810 690470
rect 131900 690230 132140 690470
rect 132230 690230 132470 690470
rect 132560 690230 132800 690470
rect 132910 690230 133150 690470
rect 122190 689900 122430 690140
rect 122520 689900 122760 690140
rect 122850 689900 123090 690140
rect 123180 689900 123420 690140
rect 123530 689900 123770 690140
rect 123860 689900 124100 690140
rect 124190 689900 124430 690140
rect 124520 689900 124760 690140
rect 124870 689900 125110 690140
rect 125200 689900 125440 690140
rect 125530 689900 125770 690140
rect 125860 689900 126100 690140
rect 126210 689900 126450 690140
rect 126540 689900 126780 690140
rect 126870 689900 127110 690140
rect 127200 689900 127440 690140
rect 127550 689900 127790 690140
rect 127880 689900 128120 690140
rect 128210 689900 128450 690140
rect 128540 689900 128780 690140
rect 128890 689900 129130 690140
rect 129220 689900 129460 690140
rect 129550 689900 129790 690140
rect 129880 689900 130120 690140
rect 130230 689900 130470 690140
rect 130560 689900 130800 690140
rect 130890 689900 131130 690140
rect 131220 689900 131460 690140
rect 131570 689900 131810 690140
rect 131900 689900 132140 690140
rect 132230 689900 132470 690140
rect 132560 689900 132800 690140
rect 132910 689900 133150 690140
rect 122190 689570 122430 689810
rect 122520 689570 122760 689810
rect 122850 689570 123090 689810
rect 123180 689570 123420 689810
rect 123530 689570 123770 689810
rect 123860 689570 124100 689810
rect 124190 689570 124430 689810
rect 124520 689570 124760 689810
rect 124870 689570 125110 689810
rect 125200 689570 125440 689810
rect 125530 689570 125770 689810
rect 125860 689570 126100 689810
rect 126210 689570 126450 689810
rect 126540 689570 126780 689810
rect 126870 689570 127110 689810
rect 127200 689570 127440 689810
rect 127550 689570 127790 689810
rect 127880 689570 128120 689810
rect 128210 689570 128450 689810
rect 128540 689570 128780 689810
rect 128890 689570 129130 689810
rect 129220 689570 129460 689810
rect 129550 689570 129790 689810
rect 129880 689570 130120 689810
rect 130230 689570 130470 689810
rect 130560 689570 130800 689810
rect 130890 689570 131130 689810
rect 131220 689570 131460 689810
rect 131570 689570 131810 689810
rect 131900 689570 132140 689810
rect 132230 689570 132470 689810
rect 132560 689570 132800 689810
rect 132910 689570 133150 689810
rect 122190 689240 122430 689480
rect 122520 689240 122760 689480
rect 122850 689240 123090 689480
rect 123180 689240 123420 689480
rect 123530 689240 123770 689480
rect 123860 689240 124100 689480
rect 124190 689240 124430 689480
rect 124520 689240 124760 689480
rect 124870 689240 125110 689480
rect 125200 689240 125440 689480
rect 125530 689240 125770 689480
rect 125860 689240 126100 689480
rect 126210 689240 126450 689480
rect 126540 689240 126780 689480
rect 126870 689240 127110 689480
rect 127200 689240 127440 689480
rect 127550 689240 127790 689480
rect 127880 689240 128120 689480
rect 128210 689240 128450 689480
rect 128540 689240 128780 689480
rect 128890 689240 129130 689480
rect 129220 689240 129460 689480
rect 129550 689240 129790 689480
rect 129880 689240 130120 689480
rect 130230 689240 130470 689480
rect 130560 689240 130800 689480
rect 130890 689240 131130 689480
rect 131220 689240 131460 689480
rect 131570 689240 131810 689480
rect 131900 689240 132140 689480
rect 132230 689240 132470 689480
rect 132560 689240 132800 689480
rect 132910 689240 133150 689480
rect 122190 688890 122430 689130
rect 122520 688890 122760 689130
rect 122850 688890 123090 689130
rect 123180 688890 123420 689130
rect 123530 688890 123770 689130
rect 123860 688890 124100 689130
rect 124190 688890 124430 689130
rect 124520 688890 124760 689130
rect 124870 688890 125110 689130
rect 125200 688890 125440 689130
rect 125530 688890 125770 689130
rect 125860 688890 126100 689130
rect 126210 688890 126450 689130
rect 126540 688890 126780 689130
rect 126870 688890 127110 689130
rect 127200 688890 127440 689130
rect 127550 688890 127790 689130
rect 127880 688890 128120 689130
rect 128210 688890 128450 689130
rect 128540 688890 128780 689130
rect 128890 688890 129130 689130
rect 129220 688890 129460 689130
rect 129550 688890 129790 689130
rect 129880 688890 130120 689130
rect 130230 688890 130470 689130
rect 130560 688890 130800 689130
rect 130890 688890 131130 689130
rect 131220 688890 131460 689130
rect 131570 688890 131810 689130
rect 131900 688890 132140 689130
rect 132230 688890 132470 689130
rect 132560 688890 132800 689130
rect 132910 688890 133150 689130
rect 122190 688560 122430 688800
rect 122520 688560 122760 688800
rect 122850 688560 123090 688800
rect 123180 688560 123420 688800
rect 123530 688560 123770 688800
rect 123860 688560 124100 688800
rect 124190 688560 124430 688800
rect 124520 688560 124760 688800
rect 124870 688560 125110 688800
rect 125200 688560 125440 688800
rect 125530 688560 125770 688800
rect 125860 688560 126100 688800
rect 126210 688560 126450 688800
rect 126540 688560 126780 688800
rect 126870 688560 127110 688800
rect 127200 688560 127440 688800
rect 127550 688560 127790 688800
rect 127880 688560 128120 688800
rect 128210 688560 128450 688800
rect 128540 688560 128780 688800
rect 128890 688560 129130 688800
rect 129220 688560 129460 688800
rect 129550 688560 129790 688800
rect 129880 688560 130120 688800
rect 130230 688560 130470 688800
rect 130560 688560 130800 688800
rect 130890 688560 131130 688800
rect 131220 688560 131460 688800
rect 131570 688560 131810 688800
rect 131900 688560 132140 688800
rect 132230 688560 132470 688800
rect 132560 688560 132800 688800
rect 132910 688560 133150 688800
rect 122190 688230 122430 688470
rect 122520 688230 122760 688470
rect 122850 688230 123090 688470
rect 123180 688230 123420 688470
rect 123530 688230 123770 688470
rect 123860 688230 124100 688470
rect 124190 688230 124430 688470
rect 124520 688230 124760 688470
rect 124870 688230 125110 688470
rect 125200 688230 125440 688470
rect 125530 688230 125770 688470
rect 125860 688230 126100 688470
rect 126210 688230 126450 688470
rect 126540 688230 126780 688470
rect 126870 688230 127110 688470
rect 127200 688230 127440 688470
rect 127550 688230 127790 688470
rect 127880 688230 128120 688470
rect 128210 688230 128450 688470
rect 128540 688230 128780 688470
rect 128890 688230 129130 688470
rect 129220 688230 129460 688470
rect 129550 688230 129790 688470
rect 129880 688230 130120 688470
rect 130230 688230 130470 688470
rect 130560 688230 130800 688470
rect 130890 688230 131130 688470
rect 131220 688230 131460 688470
rect 131570 688230 131810 688470
rect 131900 688230 132140 688470
rect 132230 688230 132470 688470
rect 132560 688230 132800 688470
rect 132910 688230 133150 688470
rect 122190 687900 122430 688140
rect 122520 687900 122760 688140
rect 122850 687900 123090 688140
rect 123180 687900 123420 688140
rect 123530 687900 123770 688140
rect 123860 687900 124100 688140
rect 124190 687900 124430 688140
rect 124520 687900 124760 688140
rect 124870 687900 125110 688140
rect 125200 687900 125440 688140
rect 125530 687900 125770 688140
rect 125860 687900 126100 688140
rect 126210 687900 126450 688140
rect 126540 687900 126780 688140
rect 126870 687900 127110 688140
rect 127200 687900 127440 688140
rect 127550 687900 127790 688140
rect 127880 687900 128120 688140
rect 128210 687900 128450 688140
rect 128540 687900 128780 688140
rect 128890 687900 129130 688140
rect 129220 687900 129460 688140
rect 129550 687900 129790 688140
rect 129880 687900 130120 688140
rect 130230 687900 130470 688140
rect 130560 687900 130800 688140
rect 130890 687900 131130 688140
rect 131220 687900 131460 688140
rect 131570 687900 131810 688140
rect 131900 687900 132140 688140
rect 132230 687900 132470 688140
rect 132560 687900 132800 688140
rect 132910 687900 133150 688140
rect 122190 687550 122430 687790
rect 122520 687550 122760 687790
rect 122850 687550 123090 687790
rect 123180 687550 123420 687790
rect 123530 687550 123770 687790
rect 123860 687550 124100 687790
rect 124190 687550 124430 687790
rect 124520 687550 124760 687790
rect 124870 687550 125110 687790
rect 125200 687550 125440 687790
rect 125530 687550 125770 687790
rect 125860 687550 126100 687790
rect 126210 687550 126450 687790
rect 126540 687550 126780 687790
rect 126870 687550 127110 687790
rect 127200 687550 127440 687790
rect 127550 687550 127790 687790
rect 127880 687550 128120 687790
rect 128210 687550 128450 687790
rect 128540 687550 128780 687790
rect 128890 687550 129130 687790
rect 129220 687550 129460 687790
rect 129550 687550 129790 687790
rect 129880 687550 130120 687790
rect 130230 687550 130470 687790
rect 130560 687550 130800 687790
rect 130890 687550 131130 687790
rect 131220 687550 131460 687790
rect 131570 687550 131810 687790
rect 131900 687550 132140 687790
rect 132230 687550 132470 687790
rect 132560 687550 132800 687790
rect 132910 687550 133150 687790
rect 122190 687220 122430 687460
rect 122520 687220 122760 687460
rect 122850 687220 123090 687460
rect 123180 687220 123420 687460
rect 123530 687220 123770 687460
rect 123860 687220 124100 687460
rect 124190 687220 124430 687460
rect 124520 687220 124760 687460
rect 124870 687220 125110 687460
rect 125200 687220 125440 687460
rect 125530 687220 125770 687460
rect 125860 687220 126100 687460
rect 126210 687220 126450 687460
rect 126540 687220 126780 687460
rect 126870 687220 127110 687460
rect 127200 687220 127440 687460
rect 127550 687220 127790 687460
rect 127880 687220 128120 687460
rect 128210 687220 128450 687460
rect 128540 687220 128780 687460
rect 128890 687220 129130 687460
rect 129220 687220 129460 687460
rect 129550 687220 129790 687460
rect 129880 687220 130120 687460
rect 130230 687220 130470 687460
rect 130560 687220 130800 687460
rect 130890 687220 131130 687460
rect 131220 687220 131460 687460
rect 131570 687220 131810 687460
rect 131900 687220 132140 687460
rect 132230 687220 132470 687460
rect 132560 687220 132800 687460
rect 132910 687220 133150 687460
rect 122190 686890 122430 687130
rect 122520 686890 122760 687130
rect 122850 686890 123090 687130
rect 123180 686890 123420 687130
rect 123530 686890 123770 687130
rect 123860 686890 124100 687130
rect 124190 686890 124430 687130
rect 124520 686890 124760 687130
rect 124870 686890 125110 687130
rect 125200 686890 125440 687130
rect 125530 686890 125770 687130
rect 125860 686890 126100 687130
rect 126210 686890 126450 687130
rect 126540 686890 126780 687130
rect 126870 686890 127110 687130
rect 127200 686890 127440 687130
rect 127550 686890 127790 687130
rect 127880 686890 128120 687130
rect 128210 686890 128450 687130
rect 128540 686890 128780 687130
rect 128890 686890 129130 687130
rect 129220 686890 129460 687130
rect 129550 686890 129790 687130
rect 129880 686890 130120 687130
rect 130230 686890 130470 687130
rect 130560 686890 130800 687130
rect 130890 686890 131130 687130
rect 131220 686890 131460 687130
rect 131570 686890 131810 687130
rect 131900 686890 132140 687130
rect 132230 686890 132470 687130
rect 132560 686890 132800 687130
rect 132910 686890 133150 687130
rect 122190 686560 122430 686800
rect 122520 686560 122760 686800
rect 122850 686560 123090 686800
rect 123180 686560 123420 686800
rect 123530 686560 123770 686800
rect 123860 686560 124100 686800
rect 124190 686560 124430 686800
rect 124520 686560 124760 686800
rect 124870 686560 125110 686800
rect 125200 686560 125440 686800
rect 125530 686560 125770 686800
rect 125860 686560 126100 686800
rect 126210 686560 126450 686800
rect 126540 686560 126780 686800
rect 126870 686560 127110 686800
rect 127200 686560 127440 686800
rect 127550 686560 127790 686800
rect 127880 686560 128120 686800
rect 128210 686560 128450 686800
rect 128540 686560 128780 686800
rect 128890 686560 129130 686800
rect 129220 686560 129460 686800
rect 129550 686560 129790 686800
rect 129880 686560 130120 686800
rect 130230 686560 130470 686800
rect 130560 686560 130800 686800
rect 130890 686560 131130 686800
rect 131220 686560 131460 686800
rect 131570 686560 131810 686800
rect 131900 686560 132140 686800
rect 132230 686560 132470 686800
rect 132560 686560 132800 686800
rect 132910 686560 133150 686800
rect 122190 686210 122430 686450
rect 122520 686210 122760 686450
rect 122850 686210 123090 686450
rect 123180 686210 123420 686450
rect 123530 686210 123770 686450
rect 123860 686210 124100 686450
rect 124190 686210 124430 686450
rect 124520 686210 124760 686450
rect 124870 686210 125110 686450
rect 125200 686210 125440 686450
rect 125530 686210 125770 686450
rect 125860 686210 126100 686450
rect 126210 686210 126450 686450
rect 126540 686210 126780 686450
rect 126870 686210 127110 686450
rect 127200 686210 127440 686450
rect 127550 686210 127790 686450
rect 127880 686210 128120 686450
rect 128210 686210 128450 686450
rect 128540 686210 128780 686450
rect 128890 686210 129130 686450
rect 129220 686210 129460 686450
rect 129550 686210 129790 686450
rect 129880 686210 130120 686450
rect 130230 686210 130470 686450
rect 130560 686210 130800 686450
rect 130890 686210 131130 686450
rect 131220 686210 131460 686450
rect 131570 686210 131810 686450
rect 131900 686210 132140 686450
rect 132230 686210 132470 686450
rect 132560 686210 132800 686450
rect 132910 686210 133150 686450
rect 122190 685880 122430 686120
rect 122520 685880 122760 686120
rect 122850 685880 123090 686120
rect 123180 685880 123420 686120
rect 123530 685880 123770 686120
rect 123860 685880 124100 686120
rect 124190 685880 124430 686120
rect 124520 685880 124760 686120
rect 124870 685880 125110 686120
rect 125200 685880 125440 686120
rect 125530 685880 125770 686120
rect 125860 685880 126100 686120
rect 126210 685880 126450 686120
rect 126540 685880 126780 686120
rect 126870 685880 127110 686120
rect 127200 685880 127440 686120
rect 127550 685880 127790 686120
rect 127880 685880 128120 686120
rect 128210 685880 128450 686120
rect 128540 685880 128780 686120
rect 128890 685880 129130 686120
rect 129220 685880 129460 686120
rect 129550 685880 129790 686120
rect 129880 685880 130120 686120
rect 130230 685880 130470 686120
rect 130560 685880 130800 686120
rect 130890 685880 131130 686120
rect 131220 685880 131460 686120
rect 131570 685880 131810 686120
rect 131900 685880 132140 686120
rect 132230 685880 132470 686120
rect 132560 685880 132800 686120
rect 132910 685880 133150 686120
rect 122190 685550 122430 685790
rect 122520 685550 122760 685790
rect 122850 685550 123090 685790
rect 123180 685550 123420 685790
rect 123530 685550 123770 685790
rect 123860 685550 124100 685790
rect 124190 685550 124430 685790
rect 124520 685550 124760 685790
rect 124870 685550 125110 685790
rect 125200 685550 125440 685790
rect 125530 685550 125770 685790
rect 125860 685550 126100 685790
rect 126210 685550 126450 685790
rect 126540 685550 126780 685790
rect 126870 685550 127110 685790
rect 127200 685550 127440 685790
rect 127550 685550 127790 685790
rect 127880 685550 128120 685790
rect 128210 685550 128450 685790
rect 128540 685550 128780 685790
rect 128890 685550 129130 685790
rect 129220 685550 129460 685790
rect 129550 685550 129790 685790
rect 129880 685550 130120 685790
rect 130230 685550 130470 685790
rect 130560 685550 130800 685790
rect 130890 685550 131130 685790
rect 131220 685550 131460 685790
rect 131570 685550 131810 685790
rect 131900 685550 132140 685790
rect 132230 685550 132470 685790
rect 132560 685550 132800 685790
rect 132910 685550 133150 685790
rect 122190 685220 122430 685460
rect 122520 685220 122760 685460
rect 122850 685220 123090 685460
rect 123180 685220 123420 685460
rect 123530 685220 123770 685460
rect 123860 685220 124100 685460
rect 124190 685220 124430 685460
rect 124520 685220 124760 685460
rect 124870 685220 125110 685460
rect 125200 685220 125440 685460
rect 125530 685220 125770 685460
rect 125860 685220 126100 685460
rect 126210 685220 126450 685460
rect 126540 685220 126780 685460
rect 126870 685220 127110 685460
rect 127200 685220 127440 685460
rect 127550 685220 127790 685460
rect 127880 685220 128120 685460
rect 128210 685220 128450 685460
rect 128540 685220 128780 685460
rect 128890 685220 129130 685460
rect 129220 685220 129460 685460
rect 129550 685220 129790 685460
rect 129880 685220 130120 685460
rect 130230 685220 130470 685460
rect 130560 685220 130800 685460
rect 130890 685220 131130 685460
rect 131220 685220 131460 685460
rect 131570 685220 131810 685460
rect 131900 685220 132140 685460
rect 132230 685220 132470 685460
rect 132560 685220 132800 685460
rect 132910 685220 133150 685460
rect 122190 684870 122430 685110
rect 122520 684870 122760 685110
rect 122850 684870 123090 685110
rect 123180 684870 123420 685110
rect 123530 684870 123770 685110
rect 123860 684870 124100 685110
rect 124190 684870 124430 685110
rect 124520 684870 124760 685110
rect 124870 684870 125110 685110
rect 125200 684870 125440 685110
rect 125530 684870 125770 685110
rect 125860 684870 126100 685110
rect 126210 684870 126450 685110
rect 126540 684870 126780 685110
rect 126870 684870 127110 685110
rect 127200 684870 127440 685110
rect 127550 684870 127790 685110
rect 127880 684870 128120 685110
rect 128210 684870 128450 685110
rect 128540 684870 128780 685110
rect 128890 684870 129130 685110
rect 129220 684870 129460 685110
rect 129550 684870 129790 685110
rect 129880 684870 130120 685110
rect 130230 684870 130470 685110
rect 130560 684870 130800 685110
rect 130890 684870 131130 685110
rect 131220 684870 131460 685110
rect 131570 684870 131810 685110
rect 131900 684870 132140 685110
rect 132230 684870 132470 685110
rect 132560 684870 132800 685110
rect 132910 684870 133150 685110
rect 122190 684540 122430 684780
rect 122520 684540 122760 684780
rect 122850 684540 123090 684780
rect 123180 684540 123420 684780
rect 123530 684540 123770 684780
rect 123860 684540 124100 684780
rect 124190 684540 124430 684780
rect 124520 684540 124760 684780
rect 124870 684540 125110 684780
rect 125200 684540 125440 684780
rect 125530 684540 125770 684780
rect 125860 684540 126100 684780
rect 126210 684540 126450 684780
rect 126540 684540 126780 684780
rect 126870 684540 127110 684780
rect 127200 684540 127440 684780
rect 127550 684540 127790 684780
rect 127880 684540 128120 684780
rect 128210 684540 128450 684780
rect 128540 684540 128780 684780
rect 128890 684540 129130 684780
rect 129220 684540 129460 684780
rect 129550 684540 129790 684780
rect 129880 684540 130120 684780
rect 130230 684540 130470 684780
rect 130560 684540 130800 684780
rect 130890 684540 131130 684780
rect 131220 684540 131460 684780
rect 131570 684540 131810 684780
rect 131900 684540 132140 684780
rect 132230 684540 132470 684780
rect 132560 684540 132800 684780
rect 132910 684540 133150 684780
rect 122190 684210 122430 684450
rect 122520 684210 122760 684450
rect 122850 684210 123090 684450
rect 123180 684210 123420 684450
rect 123530 684210 123770 684450
rect 123860 684210 124100 684450
rect 124190 684210 124430 684450
rect 124520 684210 124760 684450
rect 124870 684210 125110 684450
rect 125200 684210 125440 684450
rect 125530 684210 125770 684450
rect 125860 684210 126100 684450
rect 126210 684210 126450 684450
rect 126540 684210 126780 684450
rect 126870 684210 127110 684450
rect 127200 684210 127440 684450
rect 127550 684210 127790 684450
rect 127880 684210 128120 684450
rect 128210 684210 128450 684450
rect 128540 684210 128780 684450
rect 128890 684210 129130 684450
rect 129220 684210 129460 684450
rect 129550 684210 129790 684450
rect 129880 684210 130120 684450
rect 130230 684210 130470 684450
rect 130560 684210 130800 684450
rect 130890 684210 131130 684450
rect 131220 684210 131460 684450
rect 131570 684210 131810 684450
rect 131900 684210 132140 684450
rect 132230 684210 132470 684450
rect 132560 684210 132800 684450
rect 132910 684210 133150 684450
rect 122190 683880 122430 684120
rect 122520 683880 122760 684120
rect 122850 683880 123090 684120
rect 123180 683880 123420 684120
rect 123530 683880 123770 684120
rect 123860 683880 124100 684120
rect 124190 683880 124430 684120
rect 124520 683880 124760 684120
rect 124870 683880 125110 684120
rect 125200 683880 125440 684120
rect 125530 683880 125770 684120
rect 125860 683880 126100 684120
rect 126210 683880 126450 684120
rect 126540 683880 126780 684120
rect 126870 683880 127110 684120
rect 127200 683880 127440 684120
rect 127550 683880 127790 684120
rect 127880 683880 128120 684120
rect 128210 683880 128450 684120
rect 128540 683880 128780 684120
rect 128890 683880 129130 684120
rect 129220 683880 129460 684120
rect 129550 683880 129790 684120
rect 129880 683880 130120 684120
rect 130230 683880 130470 684120
rect 130560 683880 130800 684120
rect 130890 683880 131130 684120
rect 131220 683880 131460 684120
rect 131570 683880 131810 684120
rect 131900 683880 132140 684120
rect 132230 683880 132470 684120
rect 132560 683880 132800 684120
rect 132910 683880 133150 684120
rect 133570 694600 133810 694840
rect 133900 694600 134140 694840
rect 134230 694600 134470 694840
rect 134560 694600 134800 694840
rect 134910 694600 135150 694840
rect 135240 694600 135480 694840
rect 135570 694600 135810 694840
rect 135900 694600 136140 694840
rect 136250 694600 136490 694840
rect 136580 694600 136820 694840
rect 136910 694600 137150 694840
rect 137240 694600 137480 694840
rect 137590 694600 137830 694840
rect 137920 694600 138160 694840
rect 138250 694600 138490 694840
rect 138580 694600 138820 694840
rect 138930 694600 139170 694840
rect 139260 694600 139500 694840
rect 139590 694600 139830 694840
rect 139920 694600 140160 694840
rect 140270 694600 140510 694840
rect 140600 694600 140840 694840
rect 140930 694600 141170 694840
rect 141260 694600 141500 694840
rect 141610 694600 141850 694840
rect 141940 694600 142180 694840
rect 142270 694600 142510 694840
rect 142600 694600 142840 694840
rect 142950 694600 143190 694840
rect 143280 694600 143520 694840
rect 143610 694600 143850 694840
rect 143940 694600 144180 694840
rect 144290 694600 144530 694840
rect 133570 694250 133810 694490
rect 133900 694250 134140 694490
rect 134230 694250 134470 694490
rect 134560 694250 134800 694490
rect 134910 694250 135150 694490
rect 135240 694250 135480 694490
rect 135570 694250 135810 694490
rect 135900 694250 136140 694490
rect 136250 694250 136490 694490
rect 136580 694250 136820 694490
rect 136910 694250 137150 694490
rect 137240 694250 137480 694490
rect 137590 694250 137830 694490
rect 137920 694250 138160 694490
rect 138250 694250 138490 694490
rect 138580 694250 138820 694490
rect 138930 694250 139170 694490
rect 139260 694250 139500 694490
rect 139590 694250 139830 694490
rect 139920 694250 140160 694490
rect 140270 694250 140510 694490
rect 140600 694250 140840 694490
rect 140930 694250 141170 694490
rect 141260 694250 141500 694490
rect 141610 694250 141850 694490
rect 141940 694250 142180 694490
rect 142270 694250 142510 694490
rect 142600 694250 142840 694490
rect 142950 694250 143190 694490
rect 143280 694250 143520 694490
rect 143610 694250 143850 694490
rect 143940 694250 144180 694490
rect 144290 694250 144530 694490
rect 133570 693920 133810 694160
rect 133900 693920 134140 694160
rect 134230 693920 134470 694160
rect 134560 693920 134800 694160
rect 134910 693920 135150 694160
rect 135240 693920 135480 694160
rect 135570 693920 135810 694160
rect 135900 693920 136140 694160
rect 136250 693920 136490 694160
rect 136580 693920 136820 694160
rect 136910 693920 137150 694160
rect 137240 693920 137480 694160
rect 137590 693920 137830 694160
rect 137920 693920 138160 694160
rect 138250 693920 138490 694160
rect 138580 693920 138820 694160
rect 138930 693920 139170 694160
rect 139260 693920 139500 694160
rect 139590 693920 139830 694160
rect 139920 693920 140160 694160
rect 140270 693920 140510 694160
rect 140600 693920 140840 694160
rect 140930 693920 141170 694160
rect 141260 693920 141500 694160
rect 141610 693920 141850 694160
rect 141940 693920 142180 694160
rect 142270 693920 142510 694160
rect 142600 693920 142840 694160
rect 142950 693920 143190 694160
rect 143280 693920 143520 694160
rect 143610 693920 143850 694160
rect 143940 693920 144180 694160
rect 144290 693920 144530 694160
rect 133570 693590 133810 693830
rect 133900 693590 134140 693830
rect 134230 693590 134470 693830
rect 134560 693590 134800 693830
rect 134910 693590 135150 693830
rect 135240 693590 135480 693830
rect 135570 693590 135810 693830
rect 135900 693590 136140 693830
rect 136250 693590 136490 693830
rect 136580 693590 136820 693830
rect 136910 693590 137150 693830
rect 137240 693590 137480 693830
rect 137590 693590 137830 693830
rect 137920 693590 138160 693830
rect 138250 693590 138490 693830
rect 138580 693590 138820 693830
rect 138930 693590 139170 693830
rect 139260 693590 139500 693830
rect 139590 693590 139830 693830
rect 139920 693590 140160 693830
rect 140270 693590 140510 693830
rect 140600 693590 140840 693830
rect 140930 693590 141170 693830
rect 141260 693590 141500 693830
rect 141610 693590 141850 693830
rect 141940 693590 142180 693830
rect 142270 693590 142510 693830
rect 142600 693590 142840 693830
rect 142950 693590 143190 693830
rect 143280 693590 143520 693830
rect 143610 693590 143850 693830
rect 143940 693590 144180 693830
rect 144290 693590 144530 693830
rect 133570 693260 133810 693500
rect 133900 693260 134140 693500
rect 134230 693260 134470 693500
rect 134560 693260 134800 693500
rect 134910 693260 135150 693500
rect 135240 693260 135480 693500
rect 135570 693260 135810 693500
rect 135900 693260 136140 693500
rect 136250 693260 136490 693500
rect 136580 693260 136820 693500
rect 136910 693260 137150 693500
rect 137240 693260 137480 693500
rect 137590 693260 137830 693500
rect 137920 693260 138160 693500
rect 138250 693260 138490 693500
rect 138580 693260 138820 693500
rect 138930 693260 139170 693500
rect 139260 693260 139500 693500
rect 139590 693260 139830 693500
rect 139920 693260 140160 693500
rect 140270 693260 140510 693500
rect 140600 693260 140840 693500
rect 140930 693260 141170 693500
rect 141260 693260 141500 693500
rect 141610 693260 141850 693500
rect 141940 693260 142180 693500
rect 142270 693260 142510 693500
rect 142600 693260 142840 693500
rect 142950 693260 143190 693500
rect 143280 693260 143520 693500
rect 143610 693260 143850 693500
rect 143940 693260 144180 693500
rect 144290 693260 144530 693500
rect 133570 692910 133810 693150
rect 133900 692910 134140 693150
rect 134230 692910 134470 693150
rect 134560 692910 134800 693150
rect 134910 692910 135150 693150
rect 135240 692910 135480 693150
rect 135570 692910 135810 693150
rect 135900 692910 136140 693150
rect 136250 692910 136490 693150
rect 136580 692910 136820 693150
rect 136910 692910 137150 693150
rect 137240 692910 137480 693150
rect 137590 692910 137830 693150
rect 137920 692910 138160 693150
rect 138250 692910 138490 693150
rect 138580 692910 138820 693150
rect 138930 692910 139170 693150
rect 139260 692910 139500 693150
rect 139590 692910 139830 693150
rect 139920 692910 140160 693150
rect 140270 692910 140510 693150
rect 140600 692910 140840 693150
rect 140930 692910 141170 693150
rect 141260 692910 141500 693150
rect 141610 692910 141850 693150
rect 141940 692910 142180 693150
rect 142270 692910 142510 693150
rect 142600 692910 142840 693150
rect 142950 692910 143190 693150
rect 143280 692910 143520 693150
rect 143610 692910 143850 693150
rect 143940 692910 144180 693150
rect 144290 692910 144530 693150
rect 133570 692580 133810 692820
rect 133900 692580 134140 692820
rect 134230 692580 134470 692820
rect 134560 692580 134800 692820
rect 134910 692580 135150 692820
rect 135240 692580 135480 692820
rect 135570 692580 135810 692820
rect 135900 692580 136140 692820
rect 136250 692580 136490 692820
rect 136580 692580 136820 692820
rect 136910 692580 137150 692820
rect 137240 692580 137480 692820
rect 137590 692580 137830 692820
rect 137920 692580 138160 692820
rect 138250 692580 138490 692820
rect 138580 692580 138820 692820
rect 138930 692580 139170 692820
rect 139260 692580 139500 692820
rect 139590 692580 139830 692820
rect 139920 692580 140160 692820
rect 140270 692580 140510 692820
rect 140600 692580 140840 692820
rect 140930 692580 141170 692820
rect 141260 692580 141500 692820
rect 141610 692580 141850 692820
rect 141940 692580 142180 692820
rect 142270 692580 142510 692820
rect 142600 692580 142840 692820
rect 142950 692580 143190 692820
rect 143280 692580 143520 692820
rect 143610 692580 143850 692820
rect 143940 692580 144180 692820
rect 144290 692580 144530 692820
rect 133570 692250 133810 692490
rect 133900 692250 134140 692490
rect 134230 692250 134470 692490
rect 134560 692250 134800 692490
rect 134910 692250 135150 692490
rect 135240 692250 135480 692490
rect 135570 692250 135810 692490
rect 135900 692250 136140 692490
rect 136250 692250 136490 692490
rect 136580 692250 136820 692490
rect 136910 692250 137150 692490
rect 137240 692250 137480 692490
rect 137590 692250 137830 692490
rect 137920 692250 138160 692490
rect 138250 692250 138490 692490
rect 138580 692250 138820 692490
rect 138930 692250 139170 692490
rect 139260 692250 139500 692490
rect 139590 692250 139830 692490
rect 139920 692250 140160 692490
rect 140270 692250 140510 692490
rect 140600 692250 140840 692490
rect 140930 692250 141170 692490
rect 141260 692250 141500 692490
rect 141610 692250 141850 692490
rect 141940 692250 142180 692490
rect 142270 692250 142510 692490
rect 142600 692250 142840 692490
rect 142950 692250 143190 692490
rect 143280 692250 143520 692490
rect 143610 692250 143850 692490
rect 143940 692250 144180 692490
rect 144290 692250 144530 692490
rect 133570 691920 133810 692160
rect 133900 691920 134140 692160
rect 134230 691920 134470 692160
rect 134560 691920 134800 692160
rect 134910 691920 135150 692160
rect 135240 691920 135480 692160
rect 135570 691920 135810 692160
rect 135900 691920 136140 692160
rect 136250 691920 136490 692160
rect 136580 691920 136820 692160
rect 136910 691920 137150 692160
rect 137240 691920 137480 692160
rect 137590 691920 137830 692160
rect 137920 691920 138160 692160
rect 138250 691920 138490 692160
rect 138580 691920 138820 692160
rect 138930 691920 139170 692160
rect 139260 691920 139500 692160
rect 139590 691920 139830 692160
rect 139920 691920 140160 692160
rect 140270 691920 140510 692160
rect 140600 691920 140840 692160
rect 140930 691920 141170 692160
rect 141260 691920 141500 692160
rect 141610 691920 141850 692160
rect 141940 691920 142180 692160
rect 142270 691920 142510 692160
rect 142600 691920 142840 692160
rect 142950 691920 143190 692160
rect 143280 691920 143520 692160
rect 143610 691920 143850 692160
rect 143940 691920 144180 692160
rect 144290 691920 144530 692160
rect 133570 691570 133810 691810
rect 133900 691570 134140 691810
rect 134230 691570 134470 691810
rect 134560 691570 134800 691810
rect 134910 691570 135150 691810
rect 135240 691570 135480 691810
rect 135570 691570 135810 691810
rect 135900 691570 136140 691810
rect 136250 691570 136490 691810
rect 136580 691570 136820 691810
rect 136910 691570 137150 691810
rect 137240 691570 137480 691810
rect 137590 691570 137830 691810
rect 137920 691570 138160 691810
rect 138250 691570 138490 691810
rect 138580 691570 138820 691810
rect 138930 691570 139170 691810
rect 139260 691570 139500 691810
rect 139590 691570 139830 691810
rect 139920 691570 140160 691810
rect 140270 691570 140510 691810
rect 140600 691570 140840 691810
rect 140930 691570 141170 691810
rect 141260 691570 141500 691810
rect 141610 691570 141850 691810
rect 141940 691570 142180 691810
rect 142270 691570 142510 691810
rect 142600 691570 142840 691810
rect 142950 691570 143190 691810
rect 143280 691570 143520 691810
rect 143610 691570 143850 691810
rect 143940 691570 144180 691810
rect 144290 691570 144530 691810
rect 133570 691240 133810 691480
rect 133900 691240 134140 691480
rect 134230 691240 134470 691480
rect 134560 691240 134800 691480
rect 134910 691240 135150 691480
rect 135240 691240 135480 691480
rect 135570 691240 135810 691480
rect 135900 691240 136140 691480
rect 136250 691240 136490 691480
rect 136580 691240 136820 691480
rect 136910 691240 137150 691480
rect 137240 691240 137480 691480
rect 137590 691240 137830 691480
rect 137920 691240 138160 691480
rect 138250 691240 138490 691480
rect 138580 691240 138820 691480
rect 138930 691240 139170 691480
rect 139260 691240 139500 691480
rect 139590 691240 139830 691480
rect 139920 691240 140160 691480
rect 140270 691240 140510 691480
rect 140600 691240 140840 691480
rect 140930 691240 141170 691480
rect 141260 691240 141500 691480
rect 141610 691240 141850 691480
rect 141940 691240 142180 691480
rect 142270 691240 142510 691480
rect 142600 691240 142840 691480
rect 142950 691240 143190 691480
rect 143280 691240 143520 691480
rect 143610 691240 143850 691480
rect 143940 691240 144180 691480
rect 144290 691240 144530 691480
rect 133570 690910 133810 691150
rect 133900 690910 134140 691150
rect 134230 690910 134470 691150
rect 134560 690910 134800 691150
rect 134910 690910 135150 691150
rect 135240 690910 135480 691150
rect 135570 690910 135810 691150
rect 135900 690910 136140 691150
rect 136250 690910 136490 691150
rect 136580 690910 136820 691150
rect 136910 690910 137150 691150
rect 137240 690910 137480 691150
rect 137590 690910 137830 691150
rect 137920 690910 138160 691150
rect 138250 690910 138490 691150
rect 138580 690910 138820 691150
rect 138930 690910 139170 691150
rect 139260 690910 139500 691150
rect 139590 690910 139830 691150
rect 139920 690910 140160 691150
rect 140270 690910 140510 691150
rect 140600 690910 140840 691150
rect 140930 690910 141170 691150
rect 141260 690910 141500 691150
rect 141610 690910 141850 691150
rect 141940 690910 142180 691150
rect 142270 690910 142510 691150
rect 142600 690910 142840 691150
rect 142950 690910 143190 691150
rect 143280 690910 143520 691150
rect 143610 690910 143850 691150
rect 143940 690910 144180 691150
rect 144290 690910 144530 691150
rect 133570 690580 133810 690820
rect 133900 690580 134140 690820
rect 134230 690580 134470 690820
rect 134560 690580 134800 690820
rect 134910 690580 135150 690820
rect 135240 690580 135480 690820
rect 135570 690580 135810 690820
rect 135900 690580 136140 690820
rect 136250 690580 136490 690820
rect 136580 690580 136820 690820
rect 136910 690580 137150 690820
rect 137240 690580 137480 690820
rect 137590 690580 137830 690820
rect 137920 690580 138160 690820
rect 138250 690580 138490 690820
rect 138580 690580 138820 690820
rect 138930 690580 139170 690820
rect 139260 690580 139500 690820
rect 139590 690580 139830 690820
rect 139920 690580 140160 690820
rect 140270 690580 140510 690820
rect 140600 690580 140840 690820
rect 140930 690580 141170 690820
rect 141260 690580 141500 690820
rect 141610 690580 141850 690820
rect 141940 690580 142180 690820
rect 142270 690580 142510 690820
rect 142600 690580 142840 690820
rect 142950 690580 143190 690820
rect 143280 690580 143520 690820
rect 143610 690580 143850 690820
rect 143940 690580 144180 690820
rect 144290 690580 144530 690820
rect 133570 690230 133810 690470
rect 133900 690230 134140 690470
rect 134230 690230 134470 690470
rect 134560 690230 134800 690470
rect 134910 690230 135150 690470
rect 135240 690230 135480 690470
rect 135570 690230 135810 690470
rect 135900 690230 136140 690470
rect 136250 690230 136490 690470
rect 136580 690230 136820 690470
rect 136910 690230 137150 690470
rect 137240 690230 137480 690470
rect 137590 690230 137830 690470
rect 137920 690230 138160 690470
rect 138250 690230 138490 690470
rect 138580 690230 138820 690470
rect 138930 690230 139170 690470
rect 139260 690230 139500 690470
rect 139590 690230 139830 690470
rect 139920 690230 140160 690470
rect 140270 690230 140510 690470
rect 140600 690230 140840 690470
rect 140930 690230 141170 690470
rect 141260 690230 141500 690470
rect 141610 690230 141850 690470
rect 141940 690230 142180 690470
rect 142270 690230 142510 690470
rect 142600 690230 142840 690470
rect 142950 690230 143190 690470
rect 143280 690230 143520 690470
rect 143610 690230 143850 690470
rect 143940 690230 144180 690470
rect 144290 690230 144530 690470
rect 133570 689900 133810 690140
rect 133900 689900 134140 690140
rect 134230 689900 134470 690140
rect 134560 689900 134800 690140
rect 134910 689900 135150 690140
rect 135240 689900 135480 690140
rect 135570 689900 135810 690140
rect 135900 689900 136140 690140
rect 136250 689900 136490 690140
rect 136580 689900 136820 690140
rect 136910 689900 137150 690140
rect 137240 689900 137480 690140
rect 137590 689900 137830 690140
rect 137920 689900 138160 690140
rect 138250 689900 138490 690140
rect 138580 689900 138820 690140
rect 138930 689900 139170 690140
rect 139260 689900 139500 690140
rect 139590 689900 139830 690140
rect 139920 689900 140160 690140
rect 140270 689900 140510 690140
rect 140600 689900 140840 690140
rect 140930 689900 141170 690140
rect 141260 689900 141500 690140
rect 141610 689900 141850 690140
rect 141940 689900 142180 690140
rect 142270 689900 142510 690140
rect 142600 689900 142840 690140
rect 142950 689900 143190 690140
rect 143280 689900 143520 690140
rect 143610 689900 143850 690140
rect 143940 689900 144180 690140
rect 144290 689900 144530 690140
rect 133570 689570 133810 689810
rect 133900 689570 134140 689810
rect 134230 689570 134470 689810
rect 134560 689570 134800 689810
rect 134910 689570 135150 689810
rect 135240 689570 135480 689810
rect 135570 689570 135810 689810
rect 135900 689570 136140 689810
rect 136250 689570 136490 689810
rect 136580 689570 136820 689810
rect 136910 689570 137150 689810
rect 137240 689570 137480 689810
rect 137590 689570 137830 689810
rect 137920 689570 138160 689810
rect 138250 689570 138490 689810
rect 138580 689570 138820 689810
rect 138930 689570 139170 689810
rect 139260 689570 139500 689810
rect 139590 689570 139830 689810
rect 139920 689570 140160 689810
rect 140270 689570 140510 689810
rect 140600 689570 140840 689810
rect 140930 689570 141170 689810
rect 141260 689570 141500 689810
rect 141610 689570 141850 689810
rect 141940 689570 142180 689810
rect 142270 689570 142510 689810
rect 142600 689570 142840 689810
rect 142950 689570 143190 689810
rect 143280 689570 143520 689810
rect 143610 689570 143850 689810
rect 143940 689570 144180 689810
rect 144290 689570 144530 689810
rect 133570 689240 133810 689480
rect 133900 689240 134140 689480
rect 134230 689240 134470 689480
rect 134560 689240 134800 689480
rect 134910 689240 135150 689480
rect 135240 689240 135480 689480
rect 135570 689240 135810 689480
rect 135900 689240 136140 689480
rect 136250 689240 136490 689480
rect 136580 689240 136820 689480
rect 136910 689240 137150 689480
rect 137240 689240 137480 689480
rect 137590 689240 137830 689480
rect 137920 689240 138160 689480
rect 138250 689240 138490 689480
rect 138580 689240 138820 689480
rect 138930 689240 139170 689480
rect 139260 689240 139500 689480
rect 139590 689240 139830 689480
rect 139920 689240 140160 689480
rect 140270 689240 140510 689480
rect 140600 689240 140840 689480
rect 140930 689240 141170 689480
rect 141260 689240 141500 689480
rect 141610 689240 141850 689480
rect 141940 689240 142180 689480
rect 142270 689240 142510 689480
rect 142600 689240 142840 689480
rect 142950 689240 143190 689480
rect 143280 689240 143520 689480
rect 143610 689240 143850 689480
rect 143940 689240 144180 689480
rect 144290 689240 144530 689480
rect 133570 688890 133810 689130
rect 133900 688890 134140 689130
rect 134230 688890 134470 689130
rect 134560 688890 134800 689130
rect 134910 688890 135150 689130
rect 135240 688890 135480 689130
rect 135570 688890 135810 689130
rect 135900 688890 136140 689130
rect 136250 688890 136490 689130
rect 136580 688890 136820 689130
rect 136910 688890 137150 689130
rect 137240 688890 137480 689130
rect 137590 688890 137830 689130
rect 137920 688890 138160 689130
rect 138250 688890 138490 689130
rect 138580 688890 138820 689130
rect 138930 688890 139170 689130
rect 139260 688890 139500 689130
rect 139590 688890 139830 689130
rect 139920 688890 140160 689130
rect 140270 688890 140510 689130
rect 140600 688890 140840 689130
rect 140930 688890 141170 689130
rect 141260 688890 141500 689130
rect 141610 688890 141850 689130
rect 141940 688890 142180 689130
rect 142270 688890 142510 689130
rect 142600 688890 142840 689130
rect 142950 688890 143190 689130
rect 143280 688890 143520 689130
rect 143610 688890 143850 689130
rect 143940 688890 144180 689130
rect 144290 688890 144530 689130
rect 133570 688560 133810 688800
rect 133900 688560 134140 688800
rect 134230 688560 134470 688800
rect 134560 688560 134800 688800
rect 134910 688560 135150 688800
rect 135240 688560 135480 688800
rect 135570 688560 135810 688800
rect 135900 688560 136140 688800
rect 136250 688560 136490 688800
rect 136580 688560 136820 688800
rect 136910 688560 137150 688800
rect 137240 688560 137480 688800
rect 137590 688560 137830 688800
rect 137920 688560 138160 688800
rect 138250 688560 138490 688800
rect 138580 688560 138820 688800
rect 138930 688560 139170 688800
rect 139260 688560 139500 688800
rect 139590 688560 139830 688800
rect 139920 688560 140160 688800
rect 140270 688560 140510 688800
rect 140600 688560 140840 688800
rect 140930 688560 141170 688800
rect 141260 688560 141500 688800
rect 141610 688560 141850 688800
rect 141940 688560 142180 688800
rect 142270 688560 142510 688800
rect 142600 688560 142840 688800
rect 142950 688560 143190 688800
rect 143280 688560 143520 688800
rect 143610 688560 143850 688800
rect 143940 688560 144180 688800
rect 144290 688560 144530 688800
rect 133570 688230 133810 688470
rect 133900 688230 134140 688470
rect 134230 688230 134470 688470
rect 134560 688230 134800 688470
rect 134910 688230 135150 688470
rect 135240 688230 135480 688470
rect 135570 688230 135810 688470
rect 135900 688230 136140 688470
rect 136250 688230 136490 688470
rect 136580 688230 136820 688470
rect 136910 688230 137150 688470
rect 137240 688230 137480 688470
rect 137590 688230 137830 688470
rect 137920 688230 138160 688470
rect 138250 688230 138490 688470
rect 138580 688230 138820 688470
rect 138930 688230 139170 688470
rect 139260 688230 139500 688470
rect 139590 688230 139830 688470
rect 139920 688230 140160 688470
rect 140270 688230 140510 688470
rect 140600 688230 140840 688470
rect 140930 688230 141170 688470
rect 141260 688230 141500 688470
rect 141610 688230 141850 688470
rect 141940 688230 142180 688470
rect 142270 688230 142510 688470
rect 142600 688230 142840 688470
rect 142950 688230 143190 688470
rect 143280 688230 143520 688470
rect 143610 688230 143850 688470
rect 143940 688230 144180 688470
rect 144290 688230 144530 688470
rect 133570 687900 133810 688140
rect 133900 687900 134140 688140
rect 134230 687900 134470 688140
rect 134560 687900 134800 688140
rect 134910 687900 135150 688140
rect 135240 687900 135480 688140
rect 135570 687900 135810 688140
rect 135900 687900 136140 688140
rect 136250 687900 136490 688140
rect 136580 687900 136820 688140
rect 136910 687900 137150 688140
rect 137240 687900 137480 688140
rect 137590 687900 137830 688140
rect 137920 687900 138160 688140
rect 138250 687900 138490 688140
rect 138580 687900 138820 688140
rect 138930 687900 139170 688140
rect 139260 687900 139500 688140
rect 139590 687900 139830 688140
rect 139920 687900 140160 688140
rect 140270 687900 140510 688140
rect 140600 687900 140840 688140
rect 140930 687900 141170 688140
rect 141260 687900 141500 688140
rect 141610 687900 141850 688140
rect 141940 687900 142180 688140
rect 142270 687900 142510 688140
rect 142600 687900 142840 688140
rect 142950 687900 143190 688140
rect 143280 687900 143520 688140
rect 143610 687900 143850 688140
rect 143940 687900 144180 688140
rect 144290 687900 144530 688140
rect 133570 687550 133810 687790
rect 133900 687550 134140 687790
rect 134230 687550 134470 687790
rect 134560 687550 134800 687790
rect 134910 687550 135150 687790
rect 135240 687550 135480 687790
rect 135570 687550 135810 687790
rect 135900 687550 136140 687790
rect 136250 687550 136490 687790
rect 136580 687550 136820 687790
rect 136910 687550 137150 687790
rect 137240 687550 137480 687790
rect 137590 687550 137830 687790
rect 137920 687550 138160 687790
rect 138250 687550 138490 687790
rect 138580 687550 138820 687790
rect 138930 687550 139170 687790
rect 139260 687550 139500 687790
rect 139590 687550 139830 687790
rect 139920 687550 140160 687790
rect 140270 687550 140510 687790
rect 140600 687550 140840 687790
rect 140930 687550 141170 687790
rect 141260 687550 141500 687790
rect 141610 687550 141850 687790
rect 141940 687550 142180 687790
rect 142270 687550 142510 687790
rect 142600 687550 142840 687790
rect 142950 687550 143190 687790
rect 143280 687550 143520 687790
rect 143610 687550 143850 687790
rect 143940 687550 144180 687790
rect 144290 687550 144530 687790
rect 133570 687220 133810 687460
rect 133900 687220 134140 687460
rect 134230 687220 134470 687460
rect 134560 687220 134800 687460
rect 134910 687220 135150 687460
rect 135240 687220 135480 687460
rect 135570 687220 135810 687460
rect 135900 687220 136140 687460
rect 136250 687220 136490 687460
rect 136580 687220 136820 687460
rect 136910 687220 137150 687460
rect 137240 687220 137480 687460
rect 137590 687220 137830 687460
rect 137920 687220 138160 687460
rect 138250 687220 138490 687460
rect 138580 687220 138820 687460
rect 138930 687220 139170 687460
rect 139260 687220 139500 687460
rect 139590 687220 139830 687460
rect 139920 687220 140160 687460
rect 140270 687220 140510 687460
rect 140600 687220 140840 687460
rect 140930 687220 141170 687460
rect 141260 687220 141500 687460
rect 141610 687220 141850 687460
rect 141940 687220 142180 687460
rect 142270 687220 142510 687460
rect 142600 687220 142840 687460
rect 142950 687220 143190 687460
rect 143280 687220 143520 687460
rect 143610 687220 143850 687460
rect 143940 687220 144180 687460
rect 144290 687220 144530 687460
rect 133570 686890 133810 687130
rect 133900 686890 134140 687130
rect 134230 686890 134470 687130
rect 134560 686890 134800 687130
rect 134910 686890 135150 687130
rect 135240 686890 135480 687130
rect 135570 686890 135810 687130
rect 135900 686890 136140 687130
rect 136250 686890 136490 687130
rect 136580 686890 136820 687130
rect 136910 686890 137150 687130
rect 137240 686890 137480 687130
rect 137590 686890 137830 687130
rect 137920 686890 138160 687130
rect 138250 686890 138490 687130
rect 138580 686890 138820 687130
rect 138930 686890 139170 687130
rect 139260 686890 139500 687130
rect 139590 686890 139830 687130
rect 139920 686890 140160 687130
rect 140270 686890 140510 687130
rect 140600 686890 140840 687130
rect 140930 686890 141170 687130
rect 141260 686890 141500 687130
rect 141610 686890 141850 687130
rect 141940 686890 142180 687130
rect 142270 686890 142510 687130
rect 142600 686890 142840 687130
rect 142950 686890 143190 687130
rect 143280 686890 143520 687130
rect 143610 686890 143850 687130
rect 143940 686890 144180 687130
rect 144290 686890 144530 687130
rect 133570 686560 133810 686800
rect 133900 686560 134140 686800
rect 134230 686560 134470 686800
rect 134560 686560 134800 686800
rect 134910 686560 135150 686800
rect 135240 686560 135480 686800
rect 135570 686560 135810 686800
rect 135900 686560 136140 686800
rect 136250 686560 136490 686800
rect 136580 686560 136820 686800
rect 136910 686560 137150 686800
rect 137240 686560 137480 686800
rect 137590 686560 137830 686800
rect 137920 686560 138160 686800
rect 138250 686560 138490 686800
rect 138580 686560 138820 686800
rect 138930 686560 139170 686800
rect 139260 686560 139500 686800
rect 139590 686560 139830 686800
rect 139920 686560 140160 686800
rect 140270 686560 140510 686800
rect 140600 686560 140840 686800
rect 140930 686560 141170 686800
rect 141260 686560 141500 686800
rect 141610 686560 141850 686800
rect 141940 686560 142180 686800
rect 142270 686560 142510 686800
rect 142600 686560 142840 686800
rect 142950 686560 143190 686800
rect 143280 686560 143520 686800
rect 143610 686560 143850 686800
rect 143940 686560 144180 686800
rect 144290 686560 144530 686800
rect 133570 686210 133810 686450
rect 133900 686210 134140 686450
rect 134230 686210 134470 686450
rect 134560 686210 134800 686450
rect 134910 686210 135150 686450
rect 135240 686210 135480 686450
rect 135570 686210 135810 686450
rect 135900 686210 136140 686450
rect 136250 686210 136490 686450
rect 136580 686210 136820 686450
rect 136910 686210 137150 686450
rect 137240 686210 137480 686450
rect 137590 686210 137830 686450
rect 137920 686210 138160 686450
rect 138250 686210 138490 686450
rect 138580 686210 138820 686450
rect 138930 686210 139170 686450
rect 139260 686210 139500 686450
rect 139590 686210 139830 686450
rect 139920 686210 140160 686450
rect 140270 686210 140510 686450
rect 140600 686210 140840 686450
rect 140930 686210 141170 686450
rect 141260 686210 141500 686450
rect 141610 686210 141850 686450
rect 141940 686210 142180 686450
rect 142270 686210 142510 686450
rect 142600 686210 142840 686450
rect 142950 686210 143190 686450
rect 143280 686210 143520 686450
rect 143610 686210 143850 686450
rect 143940 686210 144180 686450
rect 144290 686210 144530 686450
rect 133570 685880 133810 686120
rect 133900 685880 134140 686120
rect 134230 685880 134470 686120
rect 134560 685880 134800 686120
rect 134910 685880 135150 686120
rect 135240 685880 135480 686120
rect 135570 685880 135810 686120
rect 135900 685880 136140 686120
rect 136250 685880 136490 686120
rect 136580 685880 136820 686120
rect 136910 685880 137150 686120
rect 137240 685880 137480 686120
rect 137590 685880 137830 686120
rect 137920 685880 138160 686120
rect 138250 685880 138490 686120
rect 138580 685880 138820 686120
rect 138930 685880 139170 686120
rect 139260 685880 139500 686120
rect 139590 685880 139830 686120
rect 139920 685880 140160 686120
rect 140270 685880 140510 686120
rect 140600 685880 140840 686120
rect 140930 685880 141170 686120
rect 141260 685880 141500 686120
rect 141610 685880 141850 686120
rect 141940 685880 142180 686120
rect 142270 685880 142510 686120
rect 142600 685880 142840 686120
rect 142950 685880 143190 686120
rect 143280 685880 143520 686120
rect 143610 685880 143850 686120
rect 143940 685880 144180 686120
rect 144290 685880 144530 686120
rect 133570 685550 133810 685790
rect 133900 685550 134140 685790
rect 134230 685550 134470 685790
rect 134560 685550 134800 685790
rect 134910 685550 135150 685790
rect 135240 685550 135480 685790
rect 135570 685550 135810 685790
rect 135900 685550 136140 685790
rect 136250 685550 136490 685790
rect 136580 685550 136820 685790
rect 136910 685550 137150 685790
rect 137240 685550 137480 685790
rect 137590 685550 137830 685790
rect 137920 685550 138160 685790
rect 138250 685550 138490 685790
rect 138580 685550 138820 685790
rect 138930 685550 139170 685790
rect 139260 685550 139500 685790
rect 139590 685550 139830 685790
rect 139920 685550 140160 685790
rect 140270 685550 140510 685790
rect 140600 685550 140840 685790
rect 140930 685550 141170 685790
rect 141260 685550 141500 685790
rect 141610 685550 141850 685790
rect 141940 685550 142180 685790
rect 142270 685550 142510 685790
rect 142600 685550 142840 685790
rect 142950 685550 143190 685790
rect 143280 685550 143520 685790
rect 143610 685550 143850 685790
rect 143940 685550 144180 685790
rect 144290 685550 144530 685790
rect 133570 685220 133810 685460
rect 133900 685220 134140 685460
rect 134230 685220 134470 685460
rect 134560 685220 134800 685460
rect 134910 685220 135150 685460
rect 135240 685220 135480 685460
rect 135570 685220 135810 685460
rect 135900 685220 136140 685460
rect 136250 685220 136490 685460
rect 136580 685220 136820 685460
rect 136910 685220 137150 685460
rect 137240 685220 137480 685460
rect 137590 685220 137830 685460
rect 137920 685220 138160 685460
rect 138250 685220 138490 685460
rect 138580 685220 138820 685460
rect 138930 685220 139170 685460
rect 139260 685220 139500 685460
rect 139590 685220 139830 685460
rect 139920 685220 140160 685460
rect 140270 685220 140510 685460
rect 140600 685220 140840 685460
rect 140930 685220 141170 685460
rect 141260 685220 141500 685460
rect 141610 685220 141850 685460
rect 141940 685220 142180 685460
rect 142270 685220 142510 685460
rect 142600 685220 142840 685460
rect 142950 685220 143190 685460
rect 143280 685220 143520 685460
rect 143610 685220 143850 685460
rect 143940 685220 144180 685460
rect 144290 685220 144530 685460
rect 133570 684870 133810 685110
rect 133900 684870 134140 685110
rect 134230 684870 134470 685110
rect 134560 684870 134800 685110
rect 134910 684870 135150 685110
rect 135240 684870 135480 685110
rect 135570 684870 135810 685110
rect 135900 684870 136140 685110
rect 136250 684870 136490 685110
rect 136580 684870 136820 685110
rect 136910 684870 137150 685110
rect 137240 684870 137480 685110
rect 137590 684870 137830 685110
rect 137920 684870 138160 685110
rect 138250 684870 138490 685110
rect 138580 684870 138820 685110
rect 138930 684870 139170 685110
rect 139260 684870 139500 685110
rect 139590 684870 139830 685110
rect 139920 684870 140160 685110
rect 140270 684870 140510 685110
rect 140600 684870 140840 685110
rect 140930 684870 141170 685110
rect 141260 684870 141500 685110
rect 141610 684870 141850 685110
rect 141940 684870 142180 685110
rect 142270 684870 142510 685110
rect 142600 684870 142840 685110
rect 142950 684870 143190 685110
rect 143280 684870 143520 685110
rect 143610 684870 143850 685110
rect 143940 684870 144180 685110
rect 144290 684870 144530 685110
rect 133570 684540 133810 684780
rect 133900 684540 134140 684780
rect 134230 684540 134470 684780
rect 134560 684540 134800 684780
rect 134910 684540 135150 684780
rect 135240 684540 135480 684780
rect 135570 684540 135810 684780
rect 135900 684540 136140 684780
rect 136250 684540 136490 684780
rect 136580 684540 136820 684780
rect 136910 684540 137150 684780
rect 137240 684540 137480 684780
rect 137590 684540 137830 684780
rect 137920 684540 138160 684780
rect 138250 684540 138490 684780
rect 138580 684540 138820 684780
rect 138930 684540 139170 684780
rect 139260 684540 139500 684780
rect 139590 684540 139830 684780
rect 139920 684540 140160 684780
rect 140270 684540 140510 684780
rect 140600 684540 140840 684780
rect 140930 684540 141170 684780
rect 141260 684540 141500 684780
rect 141610 684540 141850 684780
rect 141940 684540 142180 684780
rect 142270 684540 142510 684780
rect 142600 684540 142840 684780
rect 142950 684540 143190 684780
rect 143280 684540 143520 684780
rect 143610 684540 143850 684780
rect 143940 684540 144180 684780
rect 144290 684540 144530 684780
rect 133570 684210 133810 684450
rect 133900 684210 134140 684450
rect 134230 684210 134470 684450
rect 134560 684210 134800 684450
rect 134910 684210 135150 684450
rect 135240 684210 135480 684450
rect 135570 684210 135810 684450
rect 135900 684210 136140 684450
rect 136250 684210 136490 684450
rect 136580 684210 136820 684450
rect 136910 684210 137150 684450
rect 137240 684210 137480 684450
rect 137590 684210 137830 684450
rect 137920 684210 138160 684450
rect 138250 684210 138490 684450
rect 138580 684210 138820 684450
rect 138930 684210 139170 684450
rect 139260 684210 139500 684450
rect 139590 684210 139830 684450
rect 139920 684210 140160 684450
rect 140270 684210 140510 684450
rect 140600 684210 140840 684450
rect 140930 684210 141170 684450
rect 141260 684210 141500 684450
rect 141610 684210 141850 684450
rect 141940 684210 142180 684450
rect 142270 684210 142510 684450
rect 142600 684210 142840 684450
rect 142950 684210 143190 684450
rect 143280 684210 143520 684450
rect 143610 684210 143850 684450
rect 143940 684210 144180 684450
rect 144290 684210 144530 684450
rect 133570 683880 133810 684120
rect 133900 683880 134140 684120
rect 134230 683880 134470 684120
rect 134560 683880 134800 684120
rect 134910 683880 135150 684120
rect 135240 683880 135480 684120
rect 135570 683880 135810 684120
rect 135900 683880 136140 684120
rect 136250 683880 136490 684120
rect 136580 683880 136820 684120
rect 136910 683880 137150 684120
rect 137240 683880 137480 684120
rect 137590 683880 137830 684120
rect 137920 683880 138160 684120
rect 138250 683880 138490 684120
rect 138580 683880 138820 684120
rect 138930 683880 139170 684120
rect 139260 683880 139500 684120
rect 139590 683880 139830 684120
rect 139920 683880 140160 684120
rect 140270 683880 140510 684120
rect 140600 683880 140840 684120
rect 140930 683880 141170 684120
rect 141260 683880 141500 684120
rect 141610 683880 141850 684120
rect 141940 683880 142180 684120
rect 142270 683880 142510 684120
rect 142600 683880 142840 684120
rect 142950 683880 143190 684120
rect 143280 683880 143520 684120
rect 143610 683880 143850 684120
rect 143940 683880 144180 684120
rect 144290 683880 144530 684120
rect 144950 694600 145190 694840
rect 145280 694600 145520 694840
rect 145610 694600 145850 694840
rect 145940 694600 146180 694840
rect 146290 694600 146530 694840
rect 146620 694600 146860 694840
rect 146950 694600 147190 694840
rect 147280 694600 147520 694840
rect 147630 694600 147870 694840
rect 147960 694600 148200 694840
rect 148290 694600 148530 694840
rect 148620 694600 148860 694840
rect 148970 694600 149210 694840
rect 149300 694600 149540 694840
rect 149630 694600 149870 694840
rect 149960 694600 150200 694840
rect 150310 694600 150550 694840
rect 150640 694600 150880 694840
rect 150970 694600 151210 694840
rect 151300 694600 151540 694840
rect 151650 694600 151890 694840
rect 151980 694600 152220 694840
rect 152310 694600 152550 694840
rect 152640 694600 152880 694840
rect 152990 694600 153230 694840
rect 153320 694600 153560 694840
rect 153650 694600 153890 694840
rect 153980 694600 154220 694840
rect 154330 694600 154570 694840
rect 154660 694600 154900 694840
rect 154990 694600 155230 694840
rect 155320 694600 155560 694840
rect 155670 694600 155910 694840
rect 144950 694250 145190 694490
rect 145280 694250 145520 694490
rect 145610 694250 145850 694490
rect 145940 694250 146180 694490
rect 146290 694250 146530 694490
rect 146620 694250 146860 694490
rect 146950 694250 147190 694490
rect 147280 694250 147520 694490
rect 147630 694250 147870 694490
rect 147960 694250 148200 694490
rect 148290 694250 148530 694490
rect 148620 694250 148860 694490
rect 148970 694250 149210 694490
rect 149300 694250 149540 694490
rect 149630 694250 149870 694490
rect 149960 694250 150200 694490
rect 150310 694250 150550 694490
rect 150640 694250 150880 694490
rect 150970 694250 151210 694490
rect 151300 694250 151540 694490
rect 151650 694250 151890 694490
rect 151980 694250 152220 694490
rect 152310 694250 152550 694490
rect 152640 694250 152880 694490
rect 152990 694250 153230 694490
rect 153320 694250 153560 694490
rect 153650 694250 153890 694490
rect 153980 694250 154220 694490
rect 154330 694250 154570 694490
rect 154660 694250 154900 694490
rect 154990 694250 155230 694490
rect 155320 694250 155560 694490
rect 155670 694250 155910 694490
rect 144950 693920 145190 694160
rect 145280 693920 145520 694160
rect 145610 693920 145850 694160
rect 145940 693920 146180 694160
rect 146290 693920 146530 694160
rect 146620 693920 146860 694160
rect 146950 693920 147190 694160
rect 147280 693920 147520 694160
rect 147630 693920 147870 694160
rect 147960 693920 148200 694160
rect 148290 693920 148530 694160
rect 148620 693920 148860 694160
rect 148970 693920 149210 694160
rect 149300 693920 149540 694160
rect 149630 693920 149870 694160
rect 149960 693920 150200 694160
rect 150310 693920 150550 694160
rect 150640 693920 150880 694160
rect 150970 693920 151210 694160
rect 151300 693920 151540 694160
rect 151650 693920 151890 694160
rect 151980 693920 152220 694160
rect 152310 693920 152550 694160
rect 152640 693920 152880 694160
rect 152990 693920 153230 694160
rect 153320 693920 153560 694160
rect 153650 693920 153890 694160
rect 153980 693920 154220 694160
rect 154330 693920 154570 694160
rect 154660 693920 154900 694160
rect 154990 693920 155230 694160
rect 155320 693920 155560 694160
rect 155670 693920 155910 694160
rect 144950 693590 145190 693830
rect 145280 693590 145520 693830
rect 145610 693590 145850 693830
rect 145940 693590 146180 693830
rect 146290 693590 146530 693830
rect 146620 693590 146860 693830
rect 146950 693590 147190 693830
rect 147280 693590 147520 693830
rect 147630 693590 147870 693830
rect 147960 693590 148200 693830
rect 148290 693590 148530 693830
rect 148620 693590 148860 693830
rect 148970 693590 149210 693830
rect 149300 693590 149540 693830
rect 149630 693590 149870 693830
rect 149960 693590 150200 693830
rect 150310 693590 150550 693830
rect 150640 693590 150880 693830
rect 150970 693590 151210 693830
rect 151300 693590 151540 693830
rect 151650 693590 151890 693830
rect 151980 693590 152220 693830
rect 152310 693590 152550 693830
rect 152640 693590 152880 693830
rect 152990 693590 153230 693830
rect 153320 693590 153560 693830
rect 153650 693590 153890 693830
rect 153980 693590 154220 693830
rect 154330 693590 154570 693830
rect 154660 693590 154900 693830
rect 154990 693590 155230 693830
rect 155320 693590 155560 693830
rect 155670 693590 155910 693830
rect 144950 693260 145190 693500
rect 145280 693260 145520 693500
rect 145610 693260 145850 693500
rect 145940 693260 146180 693500
rect 146290 693260 146530 693500
rect 146620 693260 146860 693500
rect 146950 693260 147190 693500
rect 147280 693260 147520 693500
rect 147630 693260 147870 693500
rect 147960 693260 148200 693500
rect 148290 693260 148530 693500
rect 148620 693260 148860 693500
rect 148970 693260 149210 693500
rect 149300 693260 149540 693500
rect 149630 693260 149870 693500
rect 149960 693260 150200 693500
rect 150310 693260 150550 693500
rect 150640 693260 150880 693500
rect 150970 693260 151210 693500
rect 151300 693260 151540 693500
rect 151650 693260 151890 693500
rect 151980 693260 152220 693500
rect 152310 693260 152550 693500
rect 152640 693260 152880 693500
rect 152990 693260 153230 693500
rect 153320 693260 153560 693500
rect 153650 693260 153890 693500
rect 153980 693260 154220 693500
rect 154330 693260 154570 693500
rect 154660 693260 154900 693500
rect 154990 693260 155230 693500
rect 155320 693260 155560 693500
rect 155670 693260 155910 693500
rect 144950 692910 145190 693150
rect 145280 692910 145520 693150
rect 145610 692910 145850 693150
rect 145940 692910 146180 693150
rect 146290 692910 146530 693150
rect 146620 692910 146860 693150
rect 146950 692910 147190 693150
rect 147280 692910 147520 693150
rect 147630 692910 147870 693150
rect 147960 692910 148200 693150
rect 148290 692910 148530 693150
rect 148620 692910 148860 693150
rect 148970 692910 149210 693150
rect 149300 692910 149540 693150
rect 149630 692910 149870 693150
rect 149960 692910 150200 693150
rect 150310 692910 150550 693150
rect 150640 692910 150880 693150
rect 150970 692910 151210 693150
rect 151300 692910 151540 693150
rect 151650 692910 151890 693150
rect 151980 692910 152220 693150
rect 152310 692910 152550 693150
rect 152640 692910 152880 693150
rect 152990 692910 153230 693150
rect 153320 692910 153560 693150
rect 153650 692910 153890 693150
rect 153980 692910 154220 693150
rect 154330 692910 154570 693150
rect 154660 692910 154900 693150
rect 154990 692910 155230 693150
rect 155320 692910 155560 693150
rect 155670 692910 155910 693150
rect 144950 692580 145190 692820
rect 145280 692580 145520 692820
rect 145610 692580 145850 692820
rect 145940 692580 146180 692820
rect 146290 692580 146530 692820
rect 146620 692580 146860 692820
rect 146950 692580 147190 692820
rect 147280 692580 147520 692820
rect 147630 692580 147870 692820
rect 147960 692580 148200 692820
rect 148290 692580 148530 692820
rect 148620 692580 148860 692820
rect 148970 692580 149210 692820
rect 149300 692580 149540 692820
rect 149630 692580 149870 692820
rect 149960 692580 150200 692820
rect 150310 692580 150550 692820
rect 150640 692580 150880 692820
rect 150970 692580 151210 692820
rect 151300 692580 151540 692820
rect 151650 692580 151890 692820
rect 151980 692580 152220 692820
rect 152310 692580 152550 692820
rect 152640 692580 152880 692820
rect 152990 692580 153230 692820
rect 153320 692580 153560 692820
rect 153650 692580 153890 692820
rect 153980 692580 154220 692820
rect 154330 692580 154570 692820
rect 154660 692580 154900 692820
rect 154990 692580 155230 692820
rect 155320 692580 155560 692820
rect 155670 692580 155910 692820
rect 144950 692250 145190 692490
rect 145280 692250 145520 692490
rect 145610 692250 145850 692490
rect 145940 692250 146180 692490
rect 146290 692250 146530 692490
rect 146620 692250 146860 692490
rect 146950 692250 147190 692490
rect 147280 692250 147520 692490
rect 147630 692250 147870 692490
rect 147960 692250 148200 692490
rect 148290 692250 148530 692490
rect 148620 692250 148860 692490
rect 148970 692250 149210 692490
rect 149300 692250 149540 692490
rect 149630 692250 149870 692490
rect 149960 692250 150200 692490
rect 150310 692250 150550 692490
rect 150640 692250 150880 692490
rect 150970 692250 151210 692490
rect 151300 692250 151540 692490
rect 151650 692250 151890 692490
rect 151980 692250 152220 692490
rect 152310 692250 152550 692490
rect 152640 692250 152880 692490
rect 152990 692250 153230 692490
rect 153320 692250 153560 692490
rect 153650 692250 153890 692490
rect 153980 692250 154220 692490
rect 154330 692250 154570 692490
rect 154660 692250 154900 692490
rect 154990 692250 155230 692490
rect 155320 692250 155560 692490
rect 155670 692250 155910 692490
rect 144950 691920 145190 692160
rect 145280 691920 145520 692160
rect 145610 691920 145850 692160
rect 145940 691920 146180 692160
rect 146290 691920 146530 692160
rect 146620 691920 146860 692160
rect 146950 691920 147190 692160
rect 147280 691920 147520 692160
rect 147630 691920 147870 692160
rect 147960 691920 148200 692160
rect 148290 691920 148530 692160
rect 148620 691920 148860 692160
rect 148970 691920 149210 692160
rect 149300 691920 149540 692160
rect 149630 691920 149870 692160
rect 149960 691920 150200 692160
rect 150310 691920 150550 692160
rect 150640 691920 150880 692160
rect 150970 691920 151210 692160
rect 151300 691920 151540 692160
rect 151650 691920 151890 692160
rect 151980 691920 152220 692160
rect 152310 691920 152550 692160
rect 152640 691920 152880 692160
rect 152990 691920 153230 692160
rect 153320 691920 153560 692160
rect 153650 691920 153890 692160
rect 153980 691920 154220 692160
rect 154330 691920 154570 692160
rect 154660 691920 154900 692160
rect 154990 691920 155230 692160
rect 155320 691920 155560 692160
rect 155670 691920 155910 692160
rect 144950 691570 145190 691810
rect 145280 691570 145520 691810
rect 145610 691570 145850 691810
rect 145940 691570 146180 691810
rect 146290 691570 146530 691810
rect 146620 691570 146860 691810
rect 146950 691570 147190 691810
rect 147280 691570 147520 691810
rect 147630 691570 147870 691810
rect 147960 691570 148200 691810
rect 148290 691570 148530 691810
rect 148620 691570 148860 691810
rect 148970 691570 149210 691810
rect 149300 691570 149540 691810
rect 149630 691570 149870 691810
rect 149960 691570 150200 691810
rect 150310 691570 150550 691810
rect 150640 691570 150880 691810
rect 150970 691570 151210 691810
rect 151300 691570 151540 691810
rect 151650 691570 151890 691810
rect 151980 691570 152220 691810
rect 152310 691570 152550 691810
rect 152640 691570 152880 691810
rect 152990 691570 153230 691810
rect 153320 691570 153560 691810
rect 153650 691570 153890 691810
rect 153980 691570 154220 691810
rect 154330 691570 154570 691810
rect 154660 691570 154900 691810
rect 154990 691570 155230 691810
rect 155320 691570 155560 691810
rect 155670 691570 155910 691810
rect 144950 691240 145190 691480
rect 145280 691240 145520 691480
rect 145610 691240 145850 691480
rect 145940 691240 146180 691480
rect 146290 691240 146530 691480
rect 146620 691240 146860 691480
rect 146950 691240 147190 691480
rect 147280 691240 147520 691480
rect 147630 691240 147870 691480
rect 147960 691240 148200 691480
rect 148290 691240 148530 691480
rect 148620 691240 148860 691480
rect 148970 691240 149210 691480
rect 149300 691240 149540 691480
rect 149630 691240 149870 691480
rect 149960 691240 150200 691480
rect 150310 691240 150550 691480
rect 150640 691240 150880 691480
rect 150970 691240 151210 691480
rect 151300 691240 151540 691480
rect 151650 691240 151890 691480
rect 151980 691240 152220 691480
rect 152310 691240 152550 691480
rect 152640 691240 152880 691480
rect 152990 691240 153230 691480
rect 153320 691240 153560 691480
rect 153650 691240 153890 691480
rect 153980 691240 154220 691480
rect 154330 691240 154570 691480
rect 154660 691240 154900 691480
rect 154990 691240 155230 691480
rect 155320 691240 155560 691480
rect 155670 691240 155910 691480
rect 144950 690910 145190 691150
rect 145280 690910 145520 691150
rect 145610 690910 145850 691150
rect 145940 690910 146180 691150
rect 146290 690910 146530 691150
rect 146620 690910 146860 691150
rect 146950 690910 147190 691150
rect 147280 690910 147520 691150
rect 147630 690910 147870 691150
rect 147960 690910 148200 691150
rect 148290 690910 148530 691150
rect 148620 690910 148860 691150
rect 148970 690910 149210 691150
rect 149300 690910 149540 691150
rect 149630 690910 149870 691150
rect 149960 690910 150200 691150
rect 150310 690910 150550 691150
rect 150640 690910 150880 691150
rect 150970 690910 151210 691150
rect 151300 690910 151540 691150
rect 151650 690910 151890 691150
rect 151980 690910 152220 691150
rect 152310 690910 152550 691150
rect 152640 690910 152880 691150
rect 152990 690910 153230 691150
rect 153320 690910 153560 691150
rect 153650 690910 153890 691150
rect 153980 690910 154220 691150
rect 154330 690910 154570 691150
rect 154660 690910 154900 691150
rect 154990 690910 155230 691150
rect 155320 690910 155560 691150
rect 155670 690910 155910 691150
rect 144950 690580 145190 690820
rect 145280 690580 145520 690820
rect 145610 690580 145850 690820
rect 145940 690580 146180 690820
rect 146290 690580 146530 690820
rect 146620 690580 146860 690820
rect 146950 690580 147190 690820
rect 147280 690580 147520 690820
rect 147630 690580 147870 690820
rect 147960 690580 148200 690820
rect 148290 690580 148530 690820
rect 148620 690580 148860 690820
rect 148970 690580 149210 690820
rect 149300 690580 149540 690820
rect 149630 690580 149870 690820
rect 149960 690580 150200 690820
rect 150310 690580 150550 690820
rect 150640 690580 150880 690820
rect 150970 690580 151210 690820
rect 151300 690580 151540 690820
rect 151650 690580 151890 690820
rect 151980 690580 152220 690820
rect 152310 690580 152550 690820
rect 152640 690580 152880 690820
rect 152990 690580 153230 690820
rect 153320 690580 153560 690820
rect 153650 690580 153890 690820
rect 153980 690580 154220 690820
rect 154330 690580 154570 690820
rect 154660 690580 154900 690820
rect 154990 690580 155230 690820
rect 155320 690580 155560 690820
rect 155670 690580 155910 690820
rect 144950 690230 145190 690470
rect 145280 690230 145520 690470
rect 145610 690230 145850 690470
rect 145940 690230 146180 690470
rect 146290 690230 146530 690470
rect 146620 690230 146860 690470
rect 146950 690230 147190 690470
rect 147280 690230 147520 690470
rect 147630 690230 147870 690470
rect 147960 690230 148200 690470
rect 148290 690230 148530 690470
rect 148620 690230 148860 690470
rect 148970 690230 149210 690470
rect 149300 690230 149540 690470
rect 149630 690230 149870 690470
rect 149960 690230 150200 690470
rect 150310 690230 150550 690470
rect 150640 690230 150880 690470
rect 150970 690230 151210 690470
rect 151300 690230 151540 690470
rect 151650 690230 151890 690470
rect 151980 690230 152220 690470
rect 152310 690230 152550 690470
rect 152640 690230 152880 690470
rect 152990 690230 153230 690470
rect 153320 690230 153560 690470
rect 153650 690230 153890 690470
rect 153980 690230 154220 690470
rect 154330 690230 154570 690470
rect 154660 690230 154900 690470
rect 154990 690230 155230 690470
rect 155320 690230 155560 690470
rect 155670 690230 155910 690470
rect 144950 689900 145190 690140
rect 145280 689900 145520 690140
rect 145610 689900 145850 690140
rect 145940 689900 146180 690140
rect 146290 689900 146530 690140
rect 146620 689900 146860 690140
rect 146950 689900 147190 690140
rect 147280 689900 147520 690140
rect 147630 689900 147870 690140
rect 147960 689900 148200 690140
rect 148290 689900 148530 690140
rect 148620 689900 148860 690140
rect 148970 689900 149210 690140
rect 149300 689900 149540 690140
rect 149630 689900 149870 690140
rect 149960 689900 150200 690140
rect 150310 689900 150550 690140
rect 150640 689900 150880 690140
rect 150970 689900 151210 690140
rect 151300 689900 151540 690140
rect 151650 689900 151890 690140
rect 151980 689900 152220 690140
rect 152310 689900 152550 690140
rect 152640 689900 152880 690140
rect 152990 689900 153230 690140
rect 153320 689900 153560 690140
rect 153650 689900 153890 690140
rect 153980 689900 154220 690140
rect 154330 689900 154570 690140
rect 154660 689900 154900 690140
rect 154990 689900 155230 690140
rect 155320 689900 155560 690140
rect 155670 689900 155910 690140
rect 144950 689570 145190 689810
rect 145280 689570 145520 689810
rect 145610 689570 145850 689810
rect 145940 689570 146180 689810
rect 146290 689570 146530 689810
rect 146620 689570 146860 689810
rect 146950 689570 147190 689810
rect 147280 689570 147520 689810
rect 147630 689570 147870 689810
rect 147960 689570 148200 689810
rect 148290 689570 148530 689810
rect 148620 689570 148860 689810
rect 148970 689570 149210 689810
rect 149300 689570 149540 689810
rect 149630 689570 149870 689810
rect 149960 689570 150200 689810
rect 150310 689570 150550 689810
rect 150640 689570 150880 689810
rect 150970 689570 151210 689810
rect 151300 689570 151540 689810
rect 151650 689570 151890 689810
rect 151980 689570 152220 689810
rect 152310 689570 152550 689810
rect 152640 689570 152880 689810
rect 152990 689570 153230 689810
rect 153320 689570 153560 689810
rect 153650 689570 153890 689810
rect 153980 689570 154220 689810
rect 154330 689570 154570 689810
rect 154660 689570 154900 689810
rect 154990 689570 155230 689810
rect 155320 689570 155560 689810
rect 155670 689570 155910 689810
rect 144950 689240 145190 689480
rect 145280 689240 145520 689480
rect 145610 689240 145850 689480
rect 145940 689240 146180 689480
rect 146290 689240 146530 689480
rect 146620 689240 146860 689480
rect 146950 689240 147190 689480
rect 147280 689240 147520 689480
rect 147630 689240 147870 689480
rect 147960 689240 148200 689480
rect 148290 689240 148530 689480
rect 148620 689240 148860 689480
rect 148970 689240 149210 689480
rect 149300 689240 149540 689480
rect 149630 689240 149870 689480
rect 149960 689240 150200 689480
rect 150310 689240 150550 689480
rect 150640 689240 150880 689480
rect 150970 689240 151210 689480
rect 151300 689240 151540 689480
rect 151650 689240 151890 689480
rect 151980 689240 152220 689480
rect 152310 689240 152550 689480
rect 152640 689240 152880 689480
rect 152990 689240 153230 689480
rect 153320 689240 153560 689480
rect 153650 689240 153890 689480
rect 153980 689240 154220 689480
rect 154330 689240 154570 689480
rect 154660 689240 154900 689480
rect 154990 689240 155230 689480
rect 155320 689240 155560 689480
rect 155670 689240 155910 689480
rect 144950 688890 145190 689130
rect 145280 688890 145520 689130
rect 145610 688890 145850 689130
rect 145940 688890 146180 689130
rect 146290 688890 146530 689130
rect 146620 688890 146860 689130
rect 146950 688890 147190 689130
rect 147280 688890 147520 689130
rect 147630 688890 147870 689130
rect 147960 688890 148200 689130
rect 148290 688890 148530 689130
rect 148620 688890 148860 689130
rect 148970 688890 149210 689130
rect 149300 688890 149540 689130
rect 149630 688890 149870 689130
rect 149960 688890 150200 689130
rect 150310 688890 150550 689130
rect 150640 688890 150880 689130
rect 150970 688890 151210 689130
rect 151300 688890 151540 689130
rect 151650 688890 151890 689130
rect 151980 688890 152220 689130
rect 152310 688890 152550 689130
rect 152640 688890 152880 689130
rect 152990 688890 153230 689130
rect 153320 688890 153560 689130
rect 153650 688890 153890 689130
rect 153980 688890 154220 689130
rect 154330 688890 154570 689130
rect 154660 688890 154900 689130
rect 154990 688890 155230 689130
rect 155320 688890 155560 689130
rect 155670 688890 155910 689130
rect 144950 688560 145190 688800
rect 145280 688560 145520 688800
rect 145610 688560 145850 688800
rect 145940 688560 146180 688800
rect 146290 688560 146530 688800
rect 146620 688560 146860 688800
rect 146950 688560 147190 688800
rect 147280 688560 147520 688800
rect 147630 688560 147870 688800
rect 147960 688560 148200 688800
rect 148290 688560 148530 688800
rect 148620 688560 148860 688800
rect 148970 688560 149210 688800
rect 149300 688560 149540 688800
rect 149630 688560 149870 688800
rect 149960 688560 150200 688800
rect 150310 688560 150550 688800
rect 150640 688560 150880 688800
rect 150970 688560 151210 688800
rect 151300 688560 151540 688800
rect 151650 688560 151890 688800
rect 151980 688560 152220 688800
rect 152310 688560 152550 688800
rect 152640 688560 152880 688800
rect 152990 688560 153230 688800
rect 153320 688560 153560 688800
rect 153650 688560 153890 688800
rect 153980 688560 154220 688800
rect 154330 688560 154570 688800
rect 154660 688560 154900 688800
rect 154990 688560 155230 688800
rect 155320 688560 155560 688800
rect 155670 688560 155910 688800
rect 144950 688230 145190 688470
rect 145280 688230 145520 688470
rect 145610 688230 145850 688470
rect 145940 688230 146180 688470
rect 146290 688230 146530 688470
rect 146620 688230 146860 688470
rect 146950 688230 147190 688470
rect 147280 688230 147520 688470
rect 147630 688230 147870 688470
rect 147960 688230 148200 688470
rect 148290 688230 148530 688470
rect 148620 688230 148860 688470
rect 148970 688230 149210 688470
rect 149300 688230 149540 688470
rect 149630 688230 149870 688470
rect 149960 688230 150200 688470
rect 150310 688230 150550 688470
rect 150640 688230 150880 688470
rect 150970 688230 151210 688470
rect 151300 688230 151540 688470
rect 151650 688230 151890 688470
rect 151980 688230 152220 688470
rect 152310 688230 152550 688470
rect 152640 688230 152880 688470
rect 152990 688230 153230 688470
rect 153320 688230 153560 688470
rect 153650 688230 153890 688470
rect 153980 688230 154220 688470
rect 154330 688230 154570 688470
rect 154660 688230 154900 688470
rect 154990 688230 155230 688470
rect 155320 688230 155560 688470
rect 155670 688230 155910 688470
rect 144950 687900 145190 688140
rect 145280 687900 145520 688140
rect 145610 687900 145850 688140
rect 145940 687900 146180 688140
rect 146290 687900 146530 688140
rect 146620 687900 146860 688140
rect 146950 687900 147190 688140
rect 147280 687900 147520 688140
rect 147630 687900 147870 688140
rect 147960 687900 148200 688140
rect 148290 687900 148530 688140
rect 148620 687900 148860 688140
rect 148970 687900 149210 688140
rect 149300 687900 149540 688140
rect 149630 687900 149870 688140
rect 149960 687900 150200 688140
rect 150310 687900 150550 688140
rect 150640 687900 150880 688140
rect 150970 687900 151210 688140
rect 151300 687900 151540 688140
rect 151650 687900 151890 688140
rect 151980 687900 152220 688140
rect 152310 687900 152550 688140
rect 152640 687900 152880 688140
rect 152990 687900 153230 688140
rect 153320 687900 153560 688140
rect 153650 687900 153890 688140
rect 153980 687900 154220 688140
rect 154330 687900 154570 688140
rect 154660 687900 154900 688140
rect 154990 687900 155230 688140
rect 155320 687900 155560 688140
rect 155670 687900 155910 688140
rect 144950 687550 145190 687790
rect 145280 687550 145520 687790
rect 145610 687550 145850 687790
rect 145940 687550 146180 687790
rect 146290 687550 146530 687790
rect 146620 687550 146860 687790
rect 146950 687550 147190 687790
rect 147280 687550 147520 687790
rect 147630 687550 147870 687790
rect 147960 687550 148200 687790
rect 148290 687550 148530 687790
rect 148620 687550 148860 687790
rect 148970 687550 149210 687790
rect 149300 687550 149540 687790
rect 149630 687550 149870 687790
rect 149960 687550 150200 687790
rect 150310 687550 150550 687790
rect 150640 687550 150880 687790
rect 150970 687550 151210 687790
rect 151300 687550 151540 687790
rect 151650 687550 151890 687790
rect 151980 687550 152220 687790
rect 152310 687550 152550 687790
rect 152640 687550 152880 687790
rect 152990 687550 153230 687790
rect 153320 687550 153560 687790
rect 153650 687550 153890 687790
rect 153980 687550 154220 687790
rect 154330 687550 154570 687790
rect 154660 687550 154900 687790
rect 154990 687550 155230 687790
rect 155320 687550 155560 687790
rect 155670 687550 155910 687790
rect 144950 687220 145190 687460
rect 145280 687220 145520 687460
rect 145610 687220 145850 687460
rect 145940 687220 146180 687460
rect 146290 687220 146530 687460
rect 146620 687220 146860 687460
rect 146950 687220 147190 687460
rect 147280 687220 147520 687460
rect 147630 687220 147870 687460
rect 147960 687220 148200 687460
rect 148290 687220 148530 687460
rect 148620 687220 148860 687460
rect 148970 687220 149210 687460
rect 149300 687220 149540 687460
rect 149630 687220 149870 687460
rect 149960 687220 150200 687460
rect 150310 687220 150550 687460
rect 150640 687220 150880 687460
rect 150970 687220 151210 687460
rect 151300 687220 151540 687460
rect 151650 687220 151890 687460
rect 151980 687220 152220 687460
rect 152310 687220 152550 687460
rect 152640 687220 152880 687460
rect 152990 687220 153230 687460
rect 153320 687220 153560 687460
rect 153650 687220 153890 687460
rect 153980 687220 154220 687460
rect 154330 687220 154570 687460
rect 154660 687220 154900 687460
rect 154990 687220 155230 687460
rect 155320 687220 155560 687460
rect 155670 687220 155910 687460
rect 144950 686890 145190 687130
rect 145280 686890 145520 687130
rect 145610 686890 145850 687130
rect 145940 686890 146180 687130
rect 146290 686890 146530 687130
rect 146620 686890 146860 687130
rect 146950 686890 147190 687130
rect 147280 686890 147520 687130
rect 147630 686890 147870 687130
rect 147960 686890 148200 687130
rect 148290 686890 148530 687130
rect 148620 686890 148860 687130
rect 148970 686890 149210 687130
rect 149300 686890 149540 687130
rect 149630 686890 149870 687130
rect 149960 686890 150200 687130
rect 150310 686890 150550 687130
rect 150640 686890 150880 687130
rect 150970 686890 151210 687130
rect 151300 686890 151540 687130
rect 151650 686890 151890 687130
rect 151980 686890 152220 687130
rect 152310 686890 152550 687130
rect 152640 686890 152880 687130
rect 152990 686890 153230 687130
rect 153320 686890 153560 687130
rect 153650 686890 153890 687130
rect 153980 686890 154220 687130
rect 154330 686890 154570 687130
rect 154660 686890 154900 687130
rect 154990 686890 155230 687130
rect 155320 686890 155560 687130
rect 155670 686890 155910 687130
rect 144950 686560 145190 686800
rect 145280 686560 145520 686800
rect 145610 686560 145850 686800
rect 145940 686560 146180 686800
rect 146290 686560 146530 686800
rect 146620 686560 146860 686800
rect 146950 686560 147190 686800
rect 147280 686560 147520 686800
rect 147630 686560 147870 686800
rect 147960 686560 148200 686800
rect 148290 686560 148530 686800
rect 148620 686560 148860 686800
rect 148970 686560 149210 686800
rect 149300 686560 149540 686800
rect 149630 686560 149870 686800
rect 149960 686560 150200 686800
rect 150310 686560 150550 686800
rect 150640 686560 150880 686800
rect 150970 686560 151210 686800
rect 151300 686560 151540 686800
rect 151650 686560 151890 686800
rect 151980 686560 152220 686800
rect 152310 686560 152550 686800
rect 152640 686560 152880 686800
rect 152990 686560 153230 686800
rect 153320 686560 153560 686800
rect 153650 686560 153890 686800
rect 153980 686560 154220 686800
rect 154330 686560 154570 686800
rect 154660 686560 154900 686800
rect 154990 686560 155230 686800
rect 155320 686560 155560 686800
rect 155670 686560 155910 686800
rect 144950 686210 145190 686450
rect 145280 686210 145520 686450
rect 145610 686210 145850 686450
rect 145940 686210 146180 686450
rect 146290 686210 146530 686450
rect 146620 686210 146860 686450
rect 146950 686210 147190 686450
rect 147280 686210 147520 686450
rect 147630 686210 147870 686450
rect 147960 686210 148200 686450
rect 148290 686210 148530 686450
rect 148620 686210 148860 686450
rect 148970 686210 149210 686450
rect 149300 686210 149540 686450
rect 149630 686210 149870 686450
rect 149960 686210 150200 686450
rect 150310 686210 150550 686450
rect 150640 686210 150880 686450
rect 150970 686210 151210 686450
rect 151300 686210 151540 686450
rect 151650 686210 151890 686450
rect 151980 686210 152220 686450
rect 152310 686210 152550 686450
rect 152640 686210 152880 686450
rect 152990 686210 153230 686450
rect 153320 686210 153560 686450
rect 153650 686210 153890 686450
rect 153980 686210 154220 686450
rect 154330 686210 154570 686450
rect 154660 686210 154900 686450
rect 154990 686210 155230 686450
rect 155320 686210 155560 686450
rect 155670 686210 155910 686450
rect 144950 685880 145190 686120
rect 145280 685880 145520 686120
rect 145610 685880 145850 686120
rect 145940 685880 146180 686120
rect 146290 685880 146530 686120
rect 146620 685880 146860 686120
rect 146950 685880 147190 686120
rect 147280 685880 147520 686120
rect 147630 685880 147870 686120
rect 147960 685880 148200 686120
rect 148290 685880 148530 686120
rect 148620 685880 148860 686120
rect 148970 685880 149210 686120
rect 149300 685880 149540 686120
rect 149630 685880 149870 686120
rect 149960 685880 150200 686120
rect 150310 685880 150550 686120
rect 150640 685880 150880 686120
rect 150970 685880 151210 686120
rect 151300 685880 151540 686120
rect 151650 685880 151890 686120
rect 151980 685880 152220 686120
rect 152310 685880 152550 686120
rect 152640 685880 152880 686120
rect 152990 685880 153230 686120
rect 153320 685880 153560 686120
rect 153650 685880 153890 686120
rect 153980 685880 154220 686120
rect 154330 685880 154570 686120
rect 154660 685880 154900 686120
rect 154990 685880 155230 686120
rect 155320 685880 155560 686120
rect 155670 685880 155910 686120
rect 144950 685550 145190 685790
rect 145280 685550 145520 685790
rect 145610 685550 145850 685790
rect 145940 685550 146180 685790
rect 146290 685550 146530 685790
rect 146620 685550 146860 685790
rect 146950 685550 147190 685790
rect 147280 685550 147520 685790
rect 147630 685550 147870 685790
rect 147960 685550 148200 685790
rect 148290 685550 148530 685790
rect 148620 685550 148860 685790
rect 148970 685550 149210 685790
rect 149300 685550 149540 685790
rect 149630 685550 149870 685790
rect 149960 685550 150200 685790
rect 150310 685550 150550 685790
rect 150640 685550 150880 685790
rect 150970 685550 151210 685790
rect 151300 685550 151540 685790
rect 151650 685550 151890 685790
rect 151980 685550 152220 685790
rect 152310 685550 152550 685790
rect 152640 685550 152880 685790
rect 152990 685550 153230 685790
rect 153320 685550 153560 685790
rect 153650 685550 153890 685790
rect 153980 685550 154220 685790
rect 154330 685550 154570 685790
rect 154660 685550 154900 685790
rect 154990 685550 155230 685790
rect 155320 685550 155560 685790
rect 155670 685550 155910 685790
rect 144950 685220 145190 685460
rect 145280 685220 145520 685460
rect 145610 685220 145850 685460
rect 145940 685220 146180 685460
rect 146290 685220 146530 685460
rect 146620 685220 146860 685460
rect 146950 685220 147190 685460
rect 147280 685220 147520 685460
rect 147630 685220 147870 685460
rect 147960 685220 148200 685460
rect 148290 685220 148530 685460
rect 148620 685220 148860 685460
rect 148970 685220 149210 685460
rect 149300 685220 149540 685460
rect 149630 685220 149870 685460
rect 149960 685220 150200 685460
rect 150310 685220 150550 685460
rect 150640 685220 150880 685460
rect 150970 685220 151210 685460
rect 151300 685220 151540 685460
rect 151650 685220 151890 685460
rect 151980 685220 152220 685460
rect 152310 685220 152550 685460
rect 152640 685220 152880 685460
rect 152990 685220 153230 685460
rect 153320 685220 153560 685460
rect 153650 685220 153890 685460
rect 153980 685220 154220 685460
rect 154330 685220 154570 685460
rect 154660 685220 154900 685460
rect 154990 685220 155230 685460
rect 155320 685220 155560 685460
rect 155670 685220 155910 685460
rect 144950 684870 145190 685110
rect 145280 684870 145520 685110
rect 145610 684870 145850 685110
rect 145940 684870 146180 685110
rect 146290 684870 146530 685110
rect 146620 684870 146860 685110
rect 146950 684870 147190 685110
rect 147280 684870 147520 685110
rect 147630 684870 147870 685110
rect 147960 684870 148200 685110
rect 148290 684870 148530 685110
rect 148620 684870 148860 685110
rect 148970 684870 149210 685110
rect 149300 684870 149540 685110
rect 149630 684870 149870 685110
rect 149960 684870 150200 685110
rect 150310 684870 150550 685110
rect 150640 684870 150880 685110
rect 150970 684870 151210 685110
rect 151300 684870 151540 685110
rect 151650 684870 151890 685110
rect 151980 684870 152220 685110
rect 152310 684870 152550 685110
rect 152640 684870 152880 685110
rect 152990 684870 153230 685110
rect 153320 684870 153560 685110
rect 153650 684870 153890 685110
rect 153980 684870 154220 685110
rect 154330 684870 154570 685110
rect 154660 684870 154900 685110
rect 154990 684870 155230 685110
rect 155320 684870 155560 685110
rect 155670 684870 155910 685110
rect 144950 684540 145190 684780
rect 145280 684540 145520 684780
rect 145610 684540 145850 684780
rect 145940 684540 146180 684780
rect 146290 684540 146530 684780
rect 146620 684540 146860 684780
rect 146950 684540 147190 684780
rect 147280 684540 147520 684780
rect 147630 684540 147870 684780
rect 147960 684540 148200 684780
rect 148290 684540 148530 684780
rect 148620 684540 148860 684780
rect 148970 684540 149210 684780
rect 149300 684540 149540 684780
rect 149630 684540 149870 684780
rect 149960 684540 150200 684780
rect 150310 684540 150550 684780
rect 150640 684540 150880 684780
rect 150970 684540 151210 684780
rect 151300 684540 151540 684780
rect 151650 684540 151890 684780
rect 151980 684540 152220 684780
rect 152310 684540 152550 684780
rect 152640 684540 152880 684780
rect 152990 684540 153230 684780
rect 153320 684540 153560 684780
rect 153650 684540 153890 684780
rect 153980 684540 154220 684780
rect 154330 684540 154570 684780
rect 154660 684540 154900 684780
rect 154990 684540 155230 684780
rect 155320 684540 155560 684780
rect 155670 684540 155910 684780
rect 144950 684210 145190 684450
rect 145280 684210 145520 684450
rect 145610 684210 145850 684450
rect 145940 684210 146180 684450
rect 146290 684210 146530 684450
rect 146620 684210 146860 684450
rect 146950 684210 147190 684450
rect 147280 684210 147520 684450
rect 147630 684210 147870 684450
rect 147960 684210 148200 684450
rect 148290 684210 148530 684450
rect 148620 684210 148860 684450
rect 148970 684210 149210 684450
rect 149300 684210 149540 684450
rect 149630 684210 149870 684450
rect 149960 684210 150200 684450
rect 150310 684210 150550 684450
rect 150640 684210 150880 684450
rect 150970 684210 151210 684450
rect 151300 684210 151540 684450
rect 151650 684210 151890 684450
rect 151980 684210 152220 684450
rect 152310 684210 152550 684450
rect 152640 684210 152880 684450
rect 152990 684210 153230 684450
rect 153320 684210 153560 684450
rect 153650 684210 153890 684450
rect 153980 684210 154220 684450
rect 154330 684210 154570 684450
rect 154660 684210 154900 684450
rect 154990 684210 155230 684450
rect 155320 684210 155560 684450
rect 155670 684210 155910 684450
rect 144950 683880 145190 684120
rect 145280 683880 145520 684120
rect 145610 683880 145850 684120
rect 145940 683880 146180 684120
rect 146290 683880 146530 684120
rect 146620 683880 146860 684120
rect 146950 683880 147190 684120
rect 147280 683880 147520 684120
rect 147630 683880 147870 684120
rect 147960 683880 148200 684120
rect 148290 683880 148530 684120
rect 148620 683880 148860 684120
rect 148970 683880 149210 684120
rect 149300 683880 149540 684120
rect 149630 683880 149870 684120
rect 149960 683880 150200 684120
rect 150310 683880 150550 684120
rect 150640 683880 150880 684120
rect 150970 683880 151210 684120
rect 151300 683880 151540 684120
rect 151650 683880 151890 684120
rect 151980 683880 152220 684120
rect 152310 683880 152550 684120
rect 152640 683880 152880 684120
rect 152990 683880 153230 684120
rect 153320 683880 153560 684120
rect 153650 683880 153890 684120
rect 153980 683880 154220 684120
rect 154330 683880 154570 684120
rect 154660 683880 154900 684120
rect 154990 683880 155230 684120
rect 155320 683880 155560 684120
rect 155670 683880 155910 684120
rect 110810 683040 111050 683280
rect 111160 683040 111400 683280
rect 111490 683040 111730 683280
rect 111820 683040 112060 683280
rect 112150 683040 112390 683280
rect 112500 683040 112740 683280
rect 112830 683040 113070 683280
rect 113160 683040 113400 683280
rect 113490 683040 113730 683280
rect 113840 683040 114080 683280
rect 114170 683040 114410 683280
rect 114500 683040 114740 683280
rect 114830 683040 115070 683280
rect 115180 683040 115420 683280
rect 115510 683040 115750 683280
rect 115840 683040 116080 683280
rect 116170 683040 116410 683280
rect 116520 683040 116760 683280
rect 116850 683040 117090 683280
rect 117180 683040 117420 683280
rect 117510 683040 117750 683280
rect 117860 683040 118100 683280
rect 118190 683040 118430 683280
rect 118520 683040 118760 683280
rect 118850 683040 119090 683280
rect 119200 683040 119440 683280
rect 119530 683040 119770 683280
rect 119860 683040 120100 683280
rect 120190 683040 120430 683280
rect 120540 683040 120780 683280
rect 120870 683040 121110 683280
rect 121200 683040 121440 683280
rect 121530 683040 121770 683280
rect 110810 682710 111050 682950
rect 111160 682710 111400 682950
rect 111490 682710 111730 682950
rect 111820 682710 112060 682950
rect 112150 682710 112390 682950
rect 112500 682710 112740 682950
rect 112830 682710 113070 682950
rect 113160 682710 113400 682950
rect 113490 682710 113730 682950
rect 113840 682710 114080 682950
rect 114170 682710 114410 682950
rect 114500 682710 114740 682950
rect 114830 682710 115070 682950
rect 115180 682710 115420 682950
rect 115510 682710 115750 682950
rect 115840 682710 116080 682950
rect 116170 682710 116410 682950
rect 116520 682710 116760 682950
rect 116850 682710 117090 682950
rect 117180 682710 117420 682950
rect 117510 682710 117750 682950
rect 117860 682710 118100 682950
rect 118190 682710 118430 682950
rect 118520 682710 118760 682950
rect 118850 682710 119090 682950
rect 119200 682710 119440 682950
rect 119530 682710 119770 682950
rect 119860 682710 120100 682950
rect 120190 682710 120430 682950
rect 120540 682710 120780 682950
rect 120870 682710 121110 682950
rect 121200 682710 121440 682950
rect 121530 682710 121770 682950
rect 110810 682380 111050 682620
rect 111160 682380 111400 682620
rect 111490 682380 111730 682620
rect 111820 682380 112060 682620
rect 112150 682380 112390 682620
rect 112500 682380 112740 682620
rect 112830 682380 113070 682620
rect 113160 682380 113400 682620
rect 113490 682380 113730 682620
rect 113840 682380 114080 682620
rect 114170 682380 114410 682620
rect 114500 682380 114740 682620
rect 114830 682380 115070 682620
rect 115180 682380 115420 682620
rect 115510 682380 115750 682620
rect 115840 682380 116080 682620
rect 116170 682380 116410 682620
rect 116520 682380 116760 682620
rect 116850 682380 117090 682620
rect 117180 682380 117420 682620
rect 117510 682380 117750 682620
rect 117860 682380 118100 682620
rect 118190 682380 118430 682620
rect 118520 682380 118760 682620
rect 118850 682380 119090 682620
rect 119200 682380 119440 682620
rect 119530 682380 119770 682620
rect 119860 682380 120100 682620
rect 120190 682380 120430 682620
rect 120540 682380 120780 682620
rect 120870 682380 121110 682620
rect 121200 682380 121440 682620
rect 121530 682380 121770 682620
rect 110810 682050 111050 682290
rect 111160 682050 111400 682290
rect 111490 682050 111730 682290
rect 111820 682050 112060 682290
rect 112150 682050 112390 682290
rect 112500 682050 112740 682290
rect 112830 682050 113070 682290
rect 113160 682050 113400 682290
rect 113490 682050 113730 682290
rect 113840 682050 114080 682290
rect 114170 682050 114410 682290
rect 114500 682050 114740 682290
rect 114830 682050 115070 682290
rect 115180 682050 115420 682290
rect 115510 682050 115750 682290
rect 115840 682050 116080 682290
rect 116170 682050 116410 682290
rect 116520 682050 116760 682290
rect 116850 682050 117090 682290
rect 117180 682050 117420 682290
rect 117510 682050 117750 682290
rect 117860 682050 118100 682290
rect 118190 682050 118430 682290
rect 118520 682050 118760 682290
rect 118850 682050 119090 682290
rect 119200 682050 119440 682290
rect 119530 682050 119770 682290
rect 119860 682050 120100 682290
rect 120190 682050 120430 682290
rect 120540 682050 120780 682290
rect 120870 682050 121110 682290
rect 121200 682050 121440 682290
rect 121530 682050 121770 682290
rect 110810 681700 111050 681940
rect 111160 681700 111400 681940
rect 111490 681700 111730 681940
rect 111820 681700 112060 681940
rect 112150 681700 112390 681940
rect 112500 681700 112740 681940
rect 112830 681700 113070 681940
rect 113160 681700 113400 681940
rect 113490 681700 113730 681940
rect 113840 681700 114080 681940
rect 114170 681700 114410 681940
rect 114500 681700 114740 681940
rect 114830 681700 115070 681940
rect 115180 681700 115420 681940
rect 115510 681700 115750 681940
rect 115840 681700 116080 681940
rect 116170 681700 116410 681940
rect 116520 681700 116760 681940
rect 116850 681700 117090 681940
rect 117180 681700 117420 681940
rect 117510 681700 117750 681940
rect 117860 681700 118100 681940
rect 118190 681700 118430 681940
rect 118520 681700 118760 681940
rect 118850 681700 119090 681940
rect 119200 681700 119440 681940
rect 119530 681700 119770 681940
rect 119860 681700 120100 681940
rect 120190 681700 120430 681940
rect 120540 681700 120780 681940
rect 120870 681700 121110 681940
rect 121200 681700 121440 681940
rect 121530 681700 121770 681940
rect 110810 681370 111050 681610
rect 111160 681370 111400 681610
rect 111490 681370 111730 681610
rect 111820 681370 112060 681610
rect 112150 681370 112390 681610
rect 112500 681370 112740 681610
rect 112830 681370 113070 681610
rect 113160 681370 113400 681610
rect 113490 681370 113730 681610
rect 113840 681370 114080 681610
rect 114170 681370 114410 681610
rect 114500 681370 114740 681610
rect 114830 681370 115070 681610
rect 115180 681370 115420 681610
rect 115510 681370 115750 681610
rect 115840 681370 116080 681610
rect 116170 681370 116410 681610
rect 116520 681370 116760 681610
rect 116850 681370 117090 681610
rect 117180 681370 117420 681610
rect 117510 681370 117750 681610
rect 117860 681370 118100 681610
rect 118190 681370 118430 681610
rect 118520 681370 118760 681610
rect 118850 681370 119090 681610
rect 119200 681370 119440 681610
rect 119530 681370 119770 681610
rect 119860 681370 120100 681610
rect 120190 681370 120430 681610
rect 120540 681370 120780 681610
rect 120870 681370 121110 681610
rect 121200 681370 121440 681610
rect 121530 681370 121770 681610
rect 110810 681040 111050 681280
rect 111160 681040 111400 681280
rect 111490 681040 111730 681280
rect 111820 681040 112060 681280
rect 112150 681040 112390 681280
rect 112500 681040 112740 681280
rect 112830 681040 113070 681280
rect 113160 681040 113400 681280
rect 113490 681040 113730 681280
rect 113840 681040 114080 681280
rect 114170 681040 114410 681280
rect 114500 681040 114740 681280
rect 114830 681040 115070 681280
rect 115180 681040 115420 681280
rect 115510 681040 115750 681280
rect 115840 681040 116080 681280
rect 116170 681040 116410 681280
rect 116520 681040 116760 681280
rect 116850 681040 117090 681280
rect 117180 681040 117420 681280
rect 117510 681040 117750 681280
rect 117860 681040 118100 681280
rect 118190 681040 118430 681280
rect 118520 681040 118760 681280
rect 118850 681040 119090 681280
rect 119200 681040 119440 681280
rect 119530 681040 119770 681280
rect 119860 681040 120100 681280
rect 120190 681040 120430 681280
rect 120540 681040 120780 681280
rect 120870 681040 121110 681280
rect 121200 681040 121440 681280
rect 121530 681040 121770 681280
rect 110810 680710 111050 680950
rect 111160 680710 111400 680950
rect 111490 680710 111730 680950
rect 111820 680710 112060 680950
rect 112150 680710 112390 680950
rect 112500 680710 112740 680950
rect 112830 680710 113070 680950
rect 113160 680710 113400 680950
rect 113490 680710 113730 680950
rect 113840 680710 114080 680950
rect 114170 680710 114410 680950
rect 114500 680710 114740 680950
rect 114830 680710 115070 680950
rect 115180 680710 115420 680950
rect 115510 680710 115750 680950
rect 115840 680710 116080 680950
rect 116170 680710 116410 680950
rect 116520 680710 116760 680950
rect 116850 680710 117090 680950
rect 117180 680710 117420 680950
rect 117510 680710 117750 680950
rect 117860 680710 118100 680950
rect 118190 680710 118430 680950
rect 118520 680710 118760 680950
rect 118850 680710 119090 680950
rect 119200 680710 119440 680950
rect 119530 680710 119770 680950
rect 119860 680710 120100 680950
rect 120190 680710 120430 680950
rect 120540 680710 120780 680950
rect 120870 680710 121110 680950
rect 121200 680710 121440 680950
rect 121530 680710 121770 680950
rect 110810 680360 111050 680600
rect 111160 680360 111400 680600
rect 111490 680360 111730 680600
rect 111820 680360 112060 680600
rect 112150 680360 112390 680600
rect 112500 680360 112740 680600
rect 112830 680360 113070 680600
rect 113160 680360 113400 680600
rect 113490 680360 113730 680600
rect 113840 680360 114080 680600
rect 114170 680360 114410 680600
rect 114500 680360 114740 680600
rect 114830 680360 115070 680600
rect 115180 680360 115420 680600
rect 115510 680360 115750 680600
rect 115840 680360 116080 680600
rect 116170 680360 116410 680600
rect 116520 680360 116760 680600
rect 116850 680360 117090 680600
rect 117180 680360 117420 680600
rect 117510 680360 117750 680600
rect 117860 680360 118100 680600
rect 118190 680360 118430 680600
rect 118520 680360 118760 680600
rect 118850 680360 119090 680600
rect 119200 680360 119440 680600
rect 119530 680360 119770 680600
rect 119860 680360 120100 680600
rect 120190 680360 120430 680600
rect 120540 680360 120780 680600
rect 120870 680360 121110 680600
rect 121200 680360 121440 680600
rect 121530 680360 121770 680600
rect 110810 680030 111050 680270
rect 111160 680030 111400 680270
rect 111490 680030 111730 680270
rect 111820 680030 112060 680270
rect 112150 680030 112390 680270
rect 112500 680030 112740 680270
rect 112830 680030 113070 680270
rect 113160 680030 113400 680270
rect 113490 680030 113730 680270
rect 113840 680030 114080 680270
rect 114170 680030 114410 680270
rect 114500 680030 114740 680270
rect 114830 680030 115070 680270
rect 115180 680030 115420 680270
rect 115510 680030 115750 680270
rect 115840 680030 116080 680270
rect 116170 680030 116410 680270
rect 116520 680030 116760 680270
rect 116850 680030 117090 680270
rect 117180 680030 117420 680270
rect 117510 680030 117750 680270
rect 117860 680030 118100 680270
rect 118190 680030 118430 680270
rect 118520 680030 118760 680270
rect 118850 680030 119090 680270
rect 119200 680030 119440 680270
rect 119530 680030 119770 680270
rect 119860 680030 120100 680270
rect 120190 680030 120430 680270
rect 120540 680030 120780 680270
rect 120870 680030 121110 680270
rect 121200 680030 121440 680270
rect 121530 680030 121770 680270
rect 110810 679700 111050 679940
rect 111160 679700 111400 679940
rect 111490 679700 111730 679940
rect 111820 679700 112060 679940
rect 112150 679700 112390 679940
rect 112500 679700 112740 679940
rect 112830 679700 113070 679940
rect 113160 679700 113400 679940
rect 113490 679700 113730 679940
rect 113840 679700 114080 679940
rect 114170 679700 114410 679940
rect 114500 679700 114740 679940
rect 114830 679700 115070 679940
rect 115180 679700 115420 679940
rect 115510 679700 115750 679940
rect 115840 679700 116080 679940
rect 116170 679700 116410 679940
rect 116520 679700 116760 679940
rect 116850 679700 117090 679940
rect 117180 679700 117420 679940
rect 117510 679700 117750 679940
rect 117860 679700 118100 679940
rect 118190 679700 118430 679940
rect 118520 679700 118760 679940
rect 118850 679700 119090 679940
rect 119200 679700 119440 679940
rect 119530 679700 119770 679940
rect 119860 679700 120100 679940
rect 120190 679700 120430 679940
rect 120540 679700 120780 679940
rect 120870 679700 121110 679940
rect 121200 679700 121440 679940
rect 121530 679700 121770 679940
rect 110810 679370 111050 679610
rect 111160 679370 111400 679610
rect 111490 679370 111730 679610
rect 111820 679370 112060 679610
rect 112150 679370 112390 679610
rect 112500 679370 112740 679610
rect 112830 679370 113070 679610
rect 113160 679370 113400 679610
rect 113490 679370 113730 679610
rect 113840 679370 114080 679610
rect 114170 679370 114410 679610
rect 114500 679370 114740 679610
rect 114830 679370 115070 679610
rect 115180 679370 115420 679610
rect 115510 679370 115750 679610
rect 115840 679370 116080 679610
rect 116170 679370 116410 679610
rect 116520 679370 116760 679610
rect 116850 679370 117090 679610
rect 117180 679370 117420 679610
rect 117510 679370 117750 679610
rect 117860 679370 118100 679610
rect 118190 679370 118430 679610
rect 118520 679370 118760 679610
rect 118850 679370 119090 679610
rect 119200 679370 119440 679610
rect 119530 679370 119770 679610
rect 119860 679370 120100 679610
rect 120190 679370 120430 679610
rect 120540 679370 120780 679610
rect 120870 679370 121110 679610
rect 121200 679370 121440 679610
rect 121530 679370 121770 679610
rect 110810 679020 111050 679260
rect 111160 679020 111400 679260
rect 111490 679020 111730 679260
rect 111820 679020 112060 679260
rect 112150 679020 112390 679260
rect 112500 679020 112740 679260
rect 112830 679020 113070 679260
rect 113160 679020 113400 679260
rect 113490 679020 113730 679260
rect 113840 679020 114080 679260
rect 114170 679020 114410 679260
rect 114500 679020 114740 679260
rect 114830 679020 115070 679260
rect 115180 679020 115420 679260
rect 115510 679020 115750 679260
rect 115840 679020 116080 679260
rect 116170 679020 116410 679260
rect 116520 679020 116760 679260
rect 116850 679020 117090 679260
rect 117180 679020 117420 679260
rect 117510 679020 117750 679260
rect 117860 679020 118100 679260
rect 118190 679020 118430 679260
rect 118520 679020 118760 679260
rect 118850 679020 119090 679260
rect 119200 679020 119440 679260
rect 119530 679020 119770 679260
rect 119860 679020 120100 679260
rect 120190 679020 120430 679260
rect 120540 679020 120780 679260
rect 120870 679020 121110 679260
rect 121200 679020 121440 679260
rect 121530 679020 121770 679260
rect 110810 678690 111050 678930
rect 111160 678690 111400 678930
rect 111490 678690 111730 678930
rect 111820 678690 112060 678930
rect 112150 678690 112390 678930
rect 112500 678690 112740 678930
rect 112830 678690 113070 678930
rect 113160 678690 113400 678930
rect 113490 678690 113730 678930
rect 113840 678690 114080 678930
rect 114170 678690 114410 678930
rect 114500 678690 114740 678930
rect 114830 678690 115070 678930
rect 115180 678690 115420 678930
rect 115510 678690 115750 678930
rect 115840 678690 116080 678930
rect 116170 678690 116410 678930
rect 116520 678690 116760 678930
rect 116850 678690 117090 678930
rect 117180 678690 117420 678930
rect 117510 678690 117750 678930
rect 117860 678690 118100 678930
rect 118190 678690 118430 678930
rect 118520 678690 118760 678930
rect 118850 678690 119090 678930
rect 119200 678690 119440 678930
rect 119530 678690 119770 678930
rect 119860 678690 120100 678930
rect 120190 678690 120430 678930
rect 120540 678690 120780 678930
rect 120870 678690 121110 678930
rect 121200 678690 121440 678930
rect 121530 678690 121770 678930
rect 110810 678360 111050 678600
rect 111160 678360 111400 678600
rect 111490 678360 111730 678600
rect 111820 678360 112060 678600
rect 112150 678360 112390 678600
rect 112500 678360 112740 678600
rect 112830 678360 113070 678600
rect 113160 678360 113400 678600
rect 113490 678360 113730 678600
rect 113840 678360 114080 678600
rect 114170 678360 114410 678600
rect 114500 678360 114740 678600
rect 114830 678360 115070 678600
rect 115180 678360 115420 678600
rect 115510 678360 115750 678600
rect 115840 678360 116080 678600
rect 116170 678360 116410 678600
rect 116520 678360 116760 678600
rect 116850 678360 117090 678600
rect 117180 678360 117420 678600
rect 117510 678360 117750 678600
rect 117860 678360 118100 678600
rect 118190 678360 118430 678600
rect 118520 678360 118760 678600
rect 118850 678360 119090 678600
rect 119200 678360 119440 678600
rect 119530 678360 119770 678600
rect 119860 678360 120100 678600
rect 120190 678360 120430 678600
rect 120540 678360 120780 678600
rect 120870 678360 121110 678600
rect 121200 678360 121440 678600
rect 121530 678360 121770 678600
rect 110810 678030 111050 678270
rect 111160 678030 111400 678270
rect 111490 678030 111730 678270
rect 111820 678030 112060 678270
rect 112150 678030 112390 678270
rect 112500 678030 112740 678270
rect 112830 678030 113070 678270
rect 113160 678030 113400 678270
rect 113490 678030 113730 678270
rect 113840 678030 114080 678270
rect 114170 678030 114410 678270
rect 114500 678030 114740 678270
rect 114830 678030 115070 678270
rect 115180 678030 115420 678270
rect 115510 678030 115750 678270
rect 115840 678030 116080 678270
rect 116170 678030 116410 678270
rect 116520 678030 116760 678270
rect 116850 678030 117090 678270
rect 117180 678030 117420 678270
rect 117510 678030 117750 678270
rect 117860 678030 118100 678270
rect 118190 678030 118430 678270
rect 118520 678030 118760 678270
rect 118850 678030 119090 678270
rect 119200 678030 119440 678270
rect 119530 678030 119770 678270
rect 119860 678030 120100 678270
rect 120190 678030 120430 678270
rect 120540 678030 120780 678270
rect 120870 678030 121110 678270
rect 121200 678030 121440 678270
rect 121530 678030 121770 678270
rect 110810 677680 111050 677920
rect 111160 677680 111400 677920
rect 111490 677680 111730 677920
rect 111820 677680 112060 677920
rect 112150 677680 112390 677920
rect 112500 677680 112740 677920
rect 112830 677680 113070 677920
rect 113160 677680 113400 677920
rect 113490 677680 113730 677920
rect 113840 677680 114080 677920
rect 114170 677680 114410 677920
rect 114500 677680 114740 677920
rect 114830 677680 115070 677920
rect 115180 677680 115420 677920
rect 115510 677680 115750 677920
rect 115840 677680 116080 677920
rect 116170 677680 116410 677920
rect 116520 677680 116760 677920
rect 116850 677680 117090 677920
rect 117180 677680 117420 677920
rect 117510 677680 117750 677920
rect 117860 677680 118100 677920
rect 118190 677680 118430 677920
rect 118520 677680 118760 677920
rect 118850 677680 119090 677920
rect 119200 677680 119440 677920
rect 119530 677680 119770 677920
rect 119860 677680 120100 677920
rect 120190 677680 120430 677920
rect 120540 677680 120780 677920
rect 120870 677680 121110 677920
rect 121200 677680 121440 677920
rect 121530 677680 121770 677920
rect 110810 677350 111050 677590
rect 111160 677350 111400 677590
rect 111490 677350 111730 677590
rect 111820 677350 112060 677590
rect 112150 677350 112390 677590
rect 112500 677350 112740 677590
rect 112830 677350 113070 677590
rect 113160 677350 113400 677590
rect 113490 677350 113730 677590
rect 113840 677350 114080 677590
rect 114170 677350 114410 677590
rect 114500 677350 114740 677590
rect 114830 677350 115070 677590
rect 115180 677350 115420 677590
rect 115510 677350 115750 677590
rect 115840 677350 116080 677590
rect 116170 677350 116410 677590
rect 116520 677350 116760 677590
rect 116850 677350 117090 677590
rect 117180 677350 117420 677590
rect 117510 677350 117750 677590
rect 117860 677350 118100 677590
rect 118190 677350 118430 677590
rect 118520 677350 118760 677590
rect 118850 677350 119090 677590
rect 119200 677350 119440 677590
rect 119530 677350 119770 677590
rect 119860 677350 120100 677590
rect 120190 677350 120430 677590
rect 120540 677350 120780 677590
rect 120870 677350 121110 677590
rect 121200 677350 121440 677590
rect 121530 677350 121770 677590
rect 110810 677020 111050 677260
rect 111160 677020 111400 677260
rect 111490 677020 111730 677260
rect 111820 677020 112060 677260
rect 112150 677020 112390 677260
rect 112500 677020 112740 677260
rect 112830 677020 113070 677260
rect 113160 677020 113400 677260
rect 113490 677020 113730 677260
rect 113840 677020 114080 677260
rect 114170 677020 114410 677260
rect 114500 677020 114740 677260
rect 114830 677020 115070 677260
rect 115180 677020 115420 677260
rect 115510 677020 115750 677260
rect 115840 677020 116080 677260
rect 116170 677020 116410 677260
rect 116520 677020 116760 677260
rect 116850 677020 117090 677260
rect 117180 677020 117420 677260
rect 117510 677020 117750 677260
rect 117860 677020 118100 677260
rect 118190 677020 118430 677260
rect 118520 677020 118760 677260
rect 118850 677020 119090 677260
rect 119200 677020 119440 677260
rect 119530 677020 119770 677260
rect 119860 677020 120100 677260
rect 120190 677020 120430 677260
rect 120540 677020 120780 677260
rect 120870 677020 121110 677260
rect 121200 677020 121440 677260
rect 121530 677020 121770 677260
rect 110810 676690 111050 676930
rect 111160 676690 111400 676930
rect 111490 676690 111730 676930
rect 111820 676690 112060 676930
rect 112150 676690 112390 676930
rect 112500 676690 112740 676930
rect 112830 676690 113070 676930
rect 113160 676690 113400 676930
rect 113490 676690 113730 676930
rect 113840 676690 114080 676930
rect 114170 676690 114410 676930
rect 114500 676690 114740 676930
rect 114830 676690 115070 676930
rect 115180 676690 115420 676930
rect 115510 676690 115750 676930
rect 115840 676690 116080 676930
rect 116170 676690 116410 676930
rect 116520 676690 116760 676930
rect 116850 676690 117090 676930
rect 117180 676690 117420 676930
rect 117510 676690 117750 676930
rect 117860 676690 118100 676930
rect 118190 676690 118430 676930
rect 118520 676690 118760 676930
rect 118850 676690 119090 676930
rect 119200 676690 119440 676930
rect 119530 676690 119770 676930
rect 119860 676690 120100 676930
rect 120190 676690 120430 676930
rect 120540 676690 120780 676930
rect 120870 676690 121110 676930
rect 121200 676690 121440 676930
rect 121530 676690 121770 676930
rect 110810 676340 111050 676580
rect 111160 676340 111400 676580
rect 111490 676340 111730 676580
rect 111820 676340 112060 676580
rect 112150 676340 112390 676580
rect 112500 676340 112740 676580
rect 112830 676340 113070 676580
rect 113160 676340 113400 676580
rect 113490 676340 113730 676580
rect 113840 676340 114080 676580
rect 114170 676340 114410 676580
rect 114500 676340 114740 676580
rect 114830 676340 115070 676580
rect 115180 676340 115420 676580
rect 115510 676340 115750 676580
rect 115840 676340 116080 676580
rect 116170 676340 116410 676580
rect 116520 676340 116760 676580
rect 116850 676340 117090 676580
rect 117180 676340 117420 676580
rect 117510 676340 117750 676580
rect 117860 676340 118100 676580
rect 118190 676340 118430 676580
rect 118520 676340 118760 676580
rect 118850 676340 119090 676580
rect 119200 676340 119440 676580
rect 119530 676340 119770 676580
rect 119860 676340 120100 676580
rect 120190 676340 120430 676580
rect 120540 676340 120780 676580
rect 120870 676340 121110 676580
rect 121200 676340 121440 676580
rect 121530 676340 121770 676580
rect 110810 676010 111050 676250
rect 111160 676010 111400 676250
rect 111490 676010 111730 676250
rect 111820 676010 112060 676250
rect 112150 676010 112390 676250
rect 112500 676010 112740 676250
rect 112830 676010 113070 676250
rect 113160 676010 113400 676250
rect 113490 676010 113730 676250
rect 113840 676010 114080 676250
rect 114170 676010 114410 676250
rect 114500 676010 114740 676250
rect 114830 676010 115070 676250
rect 115180 676010 115420 676250
rect 115510 676010 115750 676250
rect 115840 676010 116080 676250
rect 116170 676010 116410 676250
rect 116520 676010 116760 676250
rect 116850 676010 117090 676250
rect 117180 676010 117420 676250
rect 117510 676010 117750 676250
rect 117860 676010 118100 676250
rect 118190 676010 118430 676250
rect 118520 676010 118760 676250
rect 118850 676010 119090 676250
rect 119200 676010 119440 676250
rect 119530 676010 119770 676250
rect 119860 676010 120100 676250
rect 120190 676010 120430 676250
rect 120540 676010 120780 676250
rect 120870 676010 121110 676250
rect 121200 676010 121440 676250
rect 121530 676010 121770 676250
rect 110810 675680 111050 675920
rect 111160 675680 111400 675920
rect 111490 675680 111730 675920
rect 111820 675680 112060 675920
rect 112150 675680 112390 675920
rect 112500 675680 112740 675920
rect 112830 675680 113070 675920
rect 113160 675680 113400 675920
rect 113490 675680 113730 675920
rect 113840 675680 114080 675920
rect 114170 675680 114410 675920
rect 114500 675680 114740 675920
rect 114830 675680 115070 675920
rect 115180 675680 115420 675920
rect 115510 675680 115750 675920
rect 115840 675680 116080 675920
rect 116170 675680 116410 675920
rect 116520 675680 116760 675920
rect 116850 675680 117090 675920
rect 117180 675680 117420 675920
rect 117510 675680 117750 675920
rect 117860 675680 118100 675920
rect 118190 675680 118430 675920
rect 118520 675680 118760 675920
rect 118850 675680 119090 675920
rect 119200 675680 119440 675920
rect 119530 675680 119770 675920
rect 119860 675680 120100 675920
rect 120190 675680 120430 675920
rect 120540 675680 120780 675920
rect 120870 675680 121110 675920
rect 121200 675680 121440 675920
rect 121530 675680 121770 675920
rect 110810 675350 111050 675590
rect 111160 675350 111400 675590
rect 111490 675350 111730 675590
rect 111820 675350 112060 675590
rect 112150 675350 112390 675590
rect 112500 675350 112740 675590
rect 112830 675350 113070 675590
rect 113160 675350 113400 675590
rect 113490 675350 113730 675590
rect 113840 675350 114080 675590
rect 114170 675350 114410 675590
rect 114500 675350 114740 675590
rect 114830 675350 115070 675590
rect 115180 675350 115420 675590
rect 115510 675350 115750 675590
rect 115840 675350 116080 675590
rect 116170 675350 116410 675590
rect 116520 675350 116760 675590
rect 116850 675350 117090 675590
rect 117180 675350 117420 675590
rect 117510 675350 117750 675590
rect 117860 675350 118100 675590
rect 118190 675350 118430 675590
rect 118520 675350 118760 675590
rect 118850 675350 119090 675590
rect 119200 675350 119440 675590
rect 119530 675350 119770 675590
rect 119860 675350 120100 675590
rect 120190 675350 120430 675590
rect 120540 675350 120780 675590
rect 120870 675350 121110 675590
rect 121200 675350 121440 675590
rect 121530 675350 121770 675590
rect 110810 675000 111050 675240
rect 111160 675000 111400 675240
rect 111490 675000 111730 675240
rect 111820 675000 112060 675240
rect 112150 675000 112390 675240
rect 112500 675000 112740 675240
rect 112830 675000 113070 675240
rect 113160 675000 113400 675240
rect 113490 675000 113730 675240
rect 113840 675000 114080 675240
rect 114170 675000 114410 675240
rect 114500 675000 114740 675240
rect 114830 675000 115070 675240
rect 115180 675000 115420 675240
rect 115510 675000 115750 675240
rect 115840 675000 116080 675240
rect 116170 675000 116410 675240
rect 116520 675000 116760 675240
rect 116850 675000 117090 675240
rect 117180 675000 117420 675240
rect 117510 675000 117750 675240
rect 117860 675000 118100 675240
rect 118190 675000 118430 675240
rect 118520 675000 118760 675240
rect 118850 675000 119090 675240
rect 119200 675000 119440 675240
rect 119530 675000 119770 675240
rect 119860 675000 120100 675240
rect 120190 675000 120430 675240
rect 120540 675000 120780 675240
rect 120870 675000 121110 675240
rect 121200 675000 121440 675240
rect 121530 675000 121770 675240
rect 110810 674670 111050 674910
rect 111160 674670 111400 674910
rect 111490 674670 111730 674910
rect 111820 674670 112060 674910
rect 112150 674670 112390 674910
rect 112500 674670 112740 674910
rect 112830 674670 113070 674910
rect 113160 674670 113400 674910
rect 113490 674670 113730 674910
rect 113840 674670 114080 674910
rect 114170 674670 114410 674910
rect 114500 674670 114740 674910
rect 114830 674670 115070 674910
rect 115180 674670 115420 674910
rect 115510 674670 115750 674910
rect 115840 674670 116080 674910
rect 116170 674670 116410 674910
rect 116520 674670 116760 674910
rect 116850 674670 117090 674910
rect 117180 674670 117420 674910
rect 117510 674670 117750 674910
rect 117860 674670 118100 674910
rect 118190 674670 118430 674910
rect 118520 674670 118760 674910
rect 118850 674670 119090 674910
rect 119200 674670 119440 674910
rect 119530 674670 119770 674910
rect 119860 674670 120100 674910
rect 120190 674670 120430 674910
rect 120540 674670 120780 674910
rect 120870 674670 121110 674910
rect 121200 674670 121440 674910
rect 121530 674670 121770 674910
rect 110810 674340 111050 674580
rect 111160 674340 111400 674580
rect 111490 674340 111730 674580
rect 111820 674340 112060 674580
rect 112150 674340 112390 674580
rect 112500 674340 112740 674580
rect 112830 674340 113070 674580
rect 113160 674340 113400 674580
rect 113490 674340 113730 674580
rect 113840 674340 114080 674580
rect 114170 674340 114410 674580
rect 114500 674340 114740 674580
rect 114830 674340 115070 674580
rect 115180 674340 115420 674580
rect 115510 674340 115750 674580
rect 115840 674340 116080 674580
rect 116170 674340 116410 674580
rect 116520 674340 116760 674580
rect 116850 674340 117090 674580
rect 117180 674340 117420 674580
rect 117510 674340 117750 674580
rect 117860 674340 118100 674580
rect 118190 674340 118430 674580
rect 118520 674340 118760 674580
rect 118850 674340 119090 674580
rect 119200 674340 119440 674580
rect 119530 674340 119770 674580
rect 119860 674340 120100 674580
rect 120190 674340 120430 674580
rect 120540 674340 120780 674580
rect 120870 674340 121110 674580
rect 121200 674340 121440 674580
rect 121530 674340 121770 674580
rect 110810 674010 111050 674250
rect 111160 674010 111400 674250
rect 111490 674010 111730 674250
rect 111820 674010 112060 674250
rect 112150 674010 112390 674250
rect 112500 674010 112740 674250
rect 112830 674010 113070 674250
rect 113160 674010 113400 674250
rect 113490 674010 113730 674250
rect 113840 674010 114080 674250
rect 114170 674010 114410 674250
rect 114500 674010 114740 674250
rect 114830 674010 115070 674250
rect 115180 674010 115420 674250
rect 115510 674010 115750 674250
rect 115840 674010 116080 674250
rect 116170 674010 116410 674250
rect 116520 674010 116760 674250
rect 116850 674010 117090 674250
rect 117180 674010 117420 674250
rect 117510 674010 117750 674250
rect 117860 674010 118100 674250
rect 118190 674010 118430 674250
rect 118520 674010 118760 674250
rect 118850 674010 119090 674250
rect 119200 674010 119440 674250
rect 119530 674010 119770 674250
rect 119860 674010 120100 674250
rect 120190 674010 120430 674250
rect 120540 674010 120780 674250
rect 120870 674010 121110 674250
rect 121200 674010 121440 674250
rect 121530 674010 121770 674250
rect 110810 673660 111050 673900
rect 111160 673660 111400 673900
rect 111490 673660 111730 673900
rect 111820 673660 112060 673900
rect 112150 673660 112390 673900
rect 112500 673660 112740 673900
rect 112830 673660 113070 673900
rect 113160 673660 113400 673900
rect 113490 673660 113730 673900
rect 113840 673660 114080 673900
rect 114170 673660 114410 673900
rect 114500 673660 114740 673900
rect 114830 673660 115070 673900
rect 115180 673660 115420 673900
rect 115510 673660 115750 673900
rect 115840 673660 116080 673900
rect 116170 673660 116410 673900
rect 116520 673660 116760 673900
rect 116850 673660 117090 673900
rect 117180 673660 117420 673900
rect 117510 673660 117750 673900
rect 117860 673660 118100 673900
rect 118190 673660 118430 673900
rect 118520 673660 118760 673900
rect 118850 673660 119090 673900
rect 119200 673660 119440 673900
rect 119530 673660 119770 673900
rect 119860 673660 120100 673900
rect 120190 673660 120430 673900
rect 120540 673660 120780 673900
rect 120870 673660 121110 673900
rect 121200 673660 121440 673900
rect 121530 673660 121770 673900
rect 110810 673330 111050 673570
rect 111160 673330 111400 673570
rect 111490 673330 111730 673570
rect 111820 673330 112060 673570
rect 112150 673330 112390 673570
rect 112500 673330 112740 673570
rect 112830 673330 113070 673570
rect 113160 673330 113400 673570
rect 113490 673330 113730 673570
rect 113840 673330 114080 673570
rect 114170 673330 114410 673570
rect 114500 673330 114740 673570
rect 114830 673330 115070 673570
rect 115180 673330 115420 673570
rect 115510 673330 115750 673570
rect 115840 673330 116080 673570
rect 116170 673330 116410 673570
rect 116520 673330 116760 673570
rect 116850 673330 117090 673570
rect 117180 673330 117420 673570
rect 117510 673330 117750 673570
rect 117860 673330 118100 673570
rect 118190 673330 118430 673570
rect 118520 673330 118760 673570
rect 118850 673330 119090 673570
rect 119200 673330 119440 673570
rect 119530 673330 119770 673570
rect 119860 673330 120100 673570
rect 120190 673330 120430 673570
rect 120540 673330 120780 673570
rect 120870 673330 121110 673570
rect 121200 673330 121440 673570
rect 121530 673330 121770 673570
rect 110810 673000 111050 673240
rect 111160 673000 111400 673240
rect 111490 673000 111730 673240
rect 111820 673000 112060 673240
rect 112150 673000 112390 673240
rect 112500 673000 112740 673240
rect 112830 673000 113070 673240
rect 113160 673000 113400 673240
rect 113490 673000 113730 673240
rect 113840 673000 114080 673240
rect 114170 673000 114410 673240
rect 114500 673000 114740 673240
rect 114830 673000 115070 673240
rect 115180 673000 115420 673240
rect 115510 673000 115750 673240
rect 115840 673000 116080 673240
rect 116170 673000 116410 673240
rect 116520 673000 116760 673240
rect 116850 673000 117090 673240
rect 117180 673000 117420 673240
rect 117510 673000 117750 673240
rect 117860 673000 118100 673240
rect 118190 673000 118430 673240
rect 118520 673000 118760 673240
rect 118850 673000 119090 673240
rect 119200 673000 119440 673240
rect 119530 673000 119770 673240
rect 119860 673000 120100 673240
rect 120190 673000 120430 673240
rect 120540 673000 120780 673240
rect 120870 673000 121110 673240
rect 121200 673000 121440 673240
rect 121530 673000 121770 673240
rect 110810 672670 111050 672910
rect 111160 672670 111400 672910
rect 111490 672670 111730 672910
rect 111820 672670 112060 672910
rect 112150 672670 112390 672910
rect 112500 672670 112740 672910
rect 112830 672670 113070 672910
rect 113160 672670 113400 672910
rect 113490 672670 113730 672910
rect 113840 672670 114080 672910
rect 114170 672670 114410 672910
rect 114500 672670 114740 672910
rect 114830 672670 115070 672910
rect 115180 672670 115420 672910
rect 115510 672670 115750 672910
rect 115840 672670 116080 672910
rect 116170 672670 116410 672910
rect 116520 672670 116760 672910
rect 116850 672670 117090 672910
rect 117180 672670 117420 672910
rect 117510 672670 117750 672910
rect 117860 672670 118100 672910
rect 118190 672670 118430 672910
rect 118520 672670 118760 672910
rect 118850 672670 119090 672910
rect 119200 672670 119440 672910
rect 119530 672670 119770 672910
rect 119860 672670 120100 672910
rect 120190 672670 120430 672910
rect 120540 672670 120780 672910
rect 120870 672670 121110 672910
rect 121200 672670 121440 672910
rect 121530 672670 121770 672910
rect 110810 672320 111050 672560
rect 111160 672320 111400 672560
rect 111490 672320 111730 672560
rect 111820 672320 112060 672560
rect 112150 672320 112390 672560
rect 112500 672320 112740 672560
rect 112830 672320 113070 672560
rect 113160 672320 113400 672560
rect 113490 672320 113730 672560
rect 113840 672320 114080 672560
rect 114170 672320 114410 672560
rect 114500 672320 114740 672560
rect 114830 672320 115070 672560
rect 115180 672320 115420 672560
rect 115510 672320 115750 672560
rect 115840 672320 116080 672560
rect 116170 672320 116410 672560
rect 116520 672320 116760 672560
rect 116850 672320 117090 672560
rect 117180 672320 117420 672560
rect 117510 672320 117750 672560
rect 117860 672320 118100 672560
rect 118190 672320 118430 672560
rect 118520 672320 118760 672560
rect 118850 672320 119090 672560
rect 119200 672320 119440 672560
rect 119530 672320 119770 672560
rect 119860 672320 120100 672560
rect 120190 672320 120430 672560
rect 120540 672320 120780 672560
rect 120870 672320 121110 672560
rect 121200 672320 121440 672560
rect 121530 672320 121770 672560
rect 122190 683040 122430 683280
rect 122540 683040 122780 683280
rect 122870 683040 123110 683280
rect 123200 683040 123440 683280
rect 123530 683040 123770 683280
rect 123880 683040 124120 683280
rect 124210 683040 124450 683280
rect 124540 683040 124780 683280
rect 124870 683040 125110 683280
rect 125220 683040 125460 683280
rect 125550 683040 125790 683280
rect 125880 683040 126120 683280
rect 126210 683040 126450 683280
rect 126560 683040 126800 683280
rect 126890 683040 127130 683280
rect 127220 683040 127460 683280
rect 127550 683040 127790 683280
rect 127900 683040 128140 683280
rect 128230 683040 128470 683280
rect 128560 683040 128800 683280
rect 128890 683040 129130 683280
rect 129240 683040 129480 683280
rect 129570 683040 129810 683280
rect 129900 683040 130140 683280
rect 130230 683040 130470 683280
rect 130580 683040 130820 683280
rect 130910 683040 131150 683280
rect 131240 683040 131480 683280
rect 131570 683040 131810 683280
rect 131920 683040 132160 683280
rect 132250 683040 132490 683280
rect 132580 683040 132820 683280
rect 132910 683040 133150 683280
rect 122190 682710 122430 682950
rect 122540 682710 122780 682950
rect 122870 682710 123110 682950
rect 123200 682710 123440 682950
rect 123530 682710 123770 682950
rect 123880 682710 124120 682950
rect 124210 682710 124450 682950
rect 124540 682710 124780 682950
rect 124870 682710 125110 682950
rect 125220 682710 125460 682950
rect 125550 682710 125790 682950
rect 125880 682710 126120 682950
rect 126210 682710 126450 682950
rect 126560 682710 126800 682950
rect 126890 682710 127130 682950
rect 127220 682710 127460 682950
rect 127550 682710 127790 682950
rect 127900 682710 128140 682950
rect 128230 682710 128470 682950
rect 128560 682710 128800 682950
rect 128890 682710 129130 682950
rect 129240 682710 129480 682950
rect 129570 682710 129810 682950
rect 129900 682710 130140 682950
rect 130230 682710 130470 682950
rect 130580 682710 130820 682950
rect 130910 682710 131150 682950
rect 131240 682710 131480 682950
rect 131570 682710 131810 682950
rect 131920 682710 132160 682950
rect 132250 682710 132490 682950
rect 132580 682710 132820 682950
rect 132910 682710 133150 682950
rect 122190 682380 122430 682620
rect 122540 682380 122780 682620
rect 122870 682380 123110 682620
rect 123200 682380 123440 682620
rect 123530 682380 123770 682620
rect 123880 682380 124120 682620
rect 124210 682380 124450 682620
rect 124540 682380 124780 682620
rect 124870 682380 125110 682620
rect 125220 682380 125460 682620
rect 125550 682380 125790 682620
rect 125880 682380 126120 682620
rect 126210 682380 126450 682620
rect 126560 682380 126800 682620
rect 126890 682380 127130 682620
rect 127220 682380 127460 682620
rect 127550 682380 127790 682620
rect 127900 682380 128140 682620
rect 128230 682380 128470 682620
rect 128560 682380 128800 682620
rect 128890 682380 129130 682620
rect 129240 682380 129480 682620
rect 129570 682380 129810 682620
rect 129900 682380 130140 682620
rect 130230 682380 130470 682620
rect 130580 682380 130820 682620
rect 130910 682380 131150 682620
rect 131240 682380 131480 682620
rect 131570 682380 131810 682620
rect 131920 682380 132160 682620
rect 132250 682380 132490 682620
rect 132580 682380 132820 682620
rect 132910 682380 133150 682620
rect 122190 682050 122430 682290
rect 122540 682050 122780 682290
rect 122870 682050 123110 682290
rect 123200 682050 123440 682290
rect 123530 682050 123770 682290
rect 123880 682050 124120 682290
rect 124210 682050 124450 682290
rect 124540 682050 124780 682290
rect 124870 682050 125110 682290
rect 125220 682050 125460 682290
rect 125550 682050 125790 682290
rect 125880 682050 126120 682290
rect 126210 682050 126450 682290
rect 126560 682050 126800 682290
rect 126890 682050 127130 682290
rect 127220 682050 127460 682290
rect 127550 682050 127790 682290
rect 127900 682050 128140 682290
rect 128230 682050 128470 682290
rect 128560 682050 128800 682290
rect 128890 682050 129130 682290
rect 129240 682050 129480 682290
rect 129570 682050 129810 682290
rect 129900 682050 130140 682290
rect 130230 682050 130470 682290
rect 130580 682050 130820 682290
rect 130910 682050 131150 682290
rect 131240 682050 131480 682290
rect 131570 682050 131810 682290
rect 131920 682050 132160 682290
rect 132250 682050 132490 682290
rect 132580 682050 132820 682290
rect 132910 682050 133150 682290
rect 122190 681700 122430 681940
rect 122540 681700 122780 681940
rect 122870 681700 123110 681940
rect 123200 681700 123440 681940
rect 123530 681700 123770 681940
rect 123880 681700 124120 681940
rect 124210 681700 124450 681940
rect 124540 681700 124780 681940
rect 124870 681700 125110 681940
rect 125220 681700 125460 681940
rect 125550 681700 125790 681940
rect 125880 681700 126120 681940
rect 126210 681700 126450 681940
rect 126560 681700 126800 681940
rect 126890 681700 127130 681940
rect 127220 681700 127460 681940
rect 127550 681700 127790 681940
rect 127900 681700 128140 681940
rect 128230 681700 128470 681940
rect 128560 681700 128800 681940
rect 128890 681700 129130 681940
rect 129240 681700 129480 681940
rect 129570 681700 129810 681940
rect 129900 681700 130140 681940
rect 130230 681700 130470 681940
rect 130580 681700 130820 681940
rect 130910 681700 131150 681940
rect 131240 681700 131480 681940
rect 131570 681700 131810 681940
rect 131920 681700 132160 681940
rect 132250 681700 132490 681940
rect 132580 681700 132820 681940
rect 132910 681700 133150 681940
rect 122190 681370 122430 681610
rect 122540 681370 122780 681610
rect 122870 681370 123110 681610
rect 123200 681370 123440 681610
rect 123530 681370 123770 681610
rect 123880 681370 124120 681610
rect 124210 681370 124450 681610
rect 124540 681370 124780 681610
rect 124870 681370 125110 681610
rect 125220 681370 125460 681610
rect 125550 681370 125790 681610
rect 125880 681370 126120 681610
rect 126210 681370 126450 681610
rect 126560 681370 126800 681610
rect 126890 681370 127130 681610
rect 127220 681370 127460 681610
rect 127550 681370 127790 681610
rect 127900 681370 128140 681610
rect 128230 681370 128470 681610
rect 128560 681370 128800 681610
rect 128890 681370 129130 681610
rect 129240 681370 129480 681610
rect 129570 681370 129810 681610
rect 129900 681370 130140 681610
rect 130230 681370 130470 681610
rect 130580 681370 130820 681610
rect 130910 681370 131150 681610
rect 131240 681370 131480 681610
rect 131570 681370 131810 681610
rect 131920 681370 132160 681610
rect 132250 681370 132490 681610
rect 132580 681370 132820 681610
rect 132910 681370 133150 681610
rect 122190 681040 122430 681280
rect 122540 681040 122780 681280
rect 122870 681040 123110 681280
rect 123200 681040 123440 681280
rect 123530 681040 123770 681280
rect 123880 681040 124120 681280
rect 124210 681040 124450 681280
rect 124540 681040 124780 681280
rect 124870 681040 125110 681280
rect 125220 681040 125460 681280
rect 125550 681040 125790 681280
rect 125880 681040 126120 681280
rect 126210 681040 126450 681280
rect 126560 681040 126800 681280
rect 126890 681040 127130 681280
rect 127220 681040 127460 681280
rect 127550 681040 127790 681280
rect 127900 681040 128140 681280
rect 128230 681040 128470 681280
rect 128560 681040 128800 681280
rect 128890 681040 129130 681280
rect 129240 681040 129480 681280
rect 129570 681040 129810 681280
rect 129900 681040 130140 681280
rect 130230 681040 130470 681280
rect 130580 681040 130820 681280
rect 130910 681040 131150 681280
rect 131240 681040 131480 681280
rect 131570 681040 131810 681280
rect 131920 681040 132160 681280
rect 132250 681040 132490 681280
rect 132580 681040 132820 681280
rect 132910 681040 133150 681280
rect 122190 680710 122430 680950
rect 122540 680710 122780 680950
rect 122870 680710 123110 680950
rect 123200 680710 123440 680950
rect 123530 680710 123770 680950
rect 123880 680710 124120 680950
rect 124210 680710 124450 680950
rect 124540 680710 124780 680950
rect 124870 680710 125110 680950
rect 125220 680710 125460 680950
rect 125550 680710 125790 680950
rect 125880 680710 126120 680950
rect 126210 680710 126450 680950
rect 126560 680710 126800 680950
rect 126890 680710 127130 680950
rect 127220 680710 127460 680950
rect 127550 680710 127790 680950
rect 127900 680710 128140 680950
rect 128230 680710 128470 680950
rect 128560 680710 128800 680950
rect 128890 680710 129130 680950
rect 129240 680710 129480 680950
rect 129570 680710 129810 680950
rect 129900 680710 130140 680950
rect 130230 680710 130470 680950
rect 130580 680710 130820 680950
rect 130910 680710 131150 680950
rect 131240 680710 131480 680950
rect 131570 680710 131810 680950
rect 131920 680710 132160 680950
rect 132250 680710 132490 680950
rect 132580 680710 132820 680950
rect 132910 680710 133150 680950
rect 122190 680360 122430 680600
rect 122540 680360 122780 680600
rect 122870 680360 123110 680600
rect 123200 680360 123440 680600
rect 123530 680360 123770 680600
rect 123880 680360 124120 680600
rect 124210 680360 124450 680600
rect 124540 680360 124780 680600
rect 124870 680360 125110 680600
rect 125220 680360 125460 680600
rect 125550 680360 125790 680600
rect 125880 680360 126120 680600
rect 126210 680360 126450 680600
rect 126560 680360 126800 680600
rect 126890 680360 127130 680600
rect 127220 680360 127460 680600
rect 127550 680360 127790 680600
rect 127900 680360 128140 680600
rect 128230 680360 128470 680600
rect 128560 680360 128800 680600
rect 128890 680360 129130 680600
rect 129240 680360 129480 680600
rect 129570 680360 129810 680600
rect 129900 680360 130140 680600
rect 130230 680360 130470 680600
rect 130580 680360 130820 680600
rect 130910 680360 131150 680600
rect 131240 680360 131480 680600
rect 131570 680360 131810 680600
rect 131920 680360 132160 680600
rect 132250 680360 132490 680600
rect 132580 680360 132820 680600
rect 132910 680360 133150 680600
rect 122190 680030 122430 680270
rect 122540 680030 122780 680270
rect 122870 680030 123110 680270
rect 123200 680030 123440 680270
rect 123530 680030 123770 680270
rect 123880 680030 124120 680270
rect 124210 680030 124450 680270
rect 124540 680030 124780 680270
rect 124870 680030 125110 680270
rect 125220 680030 125460 680270
rect 125550 680030 125790 680270
rect 125880 680030 126120 680270
rect 126210 680030 126450 680270
rect 126560 680030 126800 680270
rect 126890 680030 127130 680270
rect 127220 680030 127460 680270
rect 127550 680030 127790 680270
rect 127900 680030 128140 680270
rect 128230 680030 128470 680270
rect 128560 680030 128800 680270
rect 128890 680030 129130 680270
rect 129240 680030 129480 680270
rect 129570 680030 129810 680270
rect 129900 680030 130140 680270
rect 130230 680030 130470 680270
rect 130580 680030 130820 680270
rect 130910 680030 131150 680270
rect 131240 680030 131480 680270
rect 131570 680030 131810 680270
rect 131920 680030 132160 680270
rect 132250 680030 132490 680270
rect 132580 680030 132820 680270
rect 132910 680030 133150 680270
rect 122190 679700 122430 679940
rect 122540 679700 122780 679940
rect 122870 679700 123110 679940
rect 123200 679700 123440 679940
rect 123530 679700 123770 679940
rect 123880 679700 124120 679940
rect 124210 679700 124450 679940
rect 124540 679700 124780 679940
rect 124870 679700 125110 679940
rect 125220 679700 125460 679940
rect 125550 679700 125790 679940
rect 125880 679700 126120 679940
rect 126210 679700 126450 679940
rect 126560 679700 126800 679940
rect 126890 679700 127130 679940
rect 127220 679700 127460 679940
rect 127550 679700 127790 679940
rect 127900 679700 128140 679940
rect 128230 679700 128470 679940
rect 128560 679700 128800 679940
rect 128890 679700 129130 679940
rect 129240 679700 129480 679940
rect 129570 679700 129810 679940
rect 129900 679700 130140 679940
rect 130230 679700 130470 679940
rect 130580 679700 130820 679940
rect 130910 679700 131150 679940
rect 131240 679700 131480 679940
rect 131570 679700 131810 679940
rect 131920 679700 132160 679940
rect 132250 679700 132490 679940
rect 132580 679700 132820 679940
rect 132910 679700 133150 679940
rect 122190 679370 122430 679610
rect 122540 679370 122780 679610
rect 122870 679370 123110 679610
rect 123200 679370 123440 679610
rect 123530 679370 123770 679610
rect 123880 679370 124120 679610
rect 124210 679370 124450 679610
rect 124540 679370 124780 679610
rect 124870 679370 125110 679610
rect 125220 679370 125460 679610
rect 125550 679370 125790 679610
rect 125880 679370 126120 679610
rect 126210 679370 126450 679610
rect 126560 679370 126800 679610
rect 126890 679370 127130 679610
rect 127220 679370 127460 679610
rect 127550 679370 127790 679610
rect 127900 679370 128140 679610
rect 128230 679370 128470 679610
rect 128560 679370 128800 679610
rect 128890 679370 129130 679610
rect 129240 679370 129480 679610
rect 129570 679370 129810 679610
rect 129900 679370 130140 679610
rect 130230 679370 130470 679610
rect 130580 679370 130820 679610
rect 130910 679370 131150 679610
rect 131240 679370 131480 679610
rect 131570 679370 131810 679610
rect 131920 679370 132160 679610
rect 132250 679370 132490 679610
rect 132580 679370 132820 679610
rect 132910 679370 133150 679610
rect 122190 679020 122430 679260
rect 122540 679020 122780 679260
rect 122870 679020 123110 679260
rect 123200 679020 123440 679260
rect 123530 679020 123770 679260
rect 123880 679020 124120 679260
rect 124210 679020 124450 679260
rect 124540 679020 124780 679260
rect 124870 679020 125110 679260
rect 125220 679020 125460 679260
rect 125550 679020 125790 679260
rect 125880 679020 126120 679260
rect 126210 679020 126450 679260
rect 126560 679020 126800 679260
rect 126890 679020 127130 679260
rect 127220 679020 127460 679260
rect 127550 679020 127790 679260
rect 127900 679020 128140 679260
rect 128230 679020 128470 679260
rect 128560 679020 128800 679260
rect 128890 679020 129130 679260
rect 129240 679020 129480 679260
rect 129570 679020 129810 679260
rect 129900 679020 130140 679260
rect 130230 679020 130470 679260
rect 130580 679020 130820 679260
rect 130910 679020 131150 679260
rect 131240 679020 131480 679260
rect 131570 679020 131810 679260
rect 131920 679020 132160 679260
rect 132250 679020 132490 679260
rect 132580 679020 132820 679260
rect 132910 679020 133150 679260
rect 122190 678690 122430 678930
rect 122540 678690 122780 678930
rect 122870 678690 123110 678930
rect 123200 678690 123440 678930
rect 123530 678690 123770 678930
rect 123880 678690 124120 678930
rect 124210 678690 124450 678930
rect 124540 678690 124780 678930
rect 124870 678690 125110 678930
rect 125220 678690 125460 678930
rect 125550 678690 125790 678930
rect 125880 678690 126120 678930
rect 126210 678690 126450 678930
rect 126560 678690 126800 678930
rect 126890 678690 127130 678930
rect 127220 678690 127460 678930
rect 127550 678690 127790 678930
rect 127900 678690 128140 678930
rect 128230 678690 128470 678930
rect 128560 678690 128800 678930
rect 128890 678690 129130 678930
rect 129240 678690 129480 678930
rect 129570 678690 129810 678930
rect 129900 678690 130140 678930
rect 130230 678690 130470 678930
rect 130580 678690 130820 678930
rect 130910 678690 131150 678930
rect 131240 678690 131480 678930
rect 131570 678690 131810 678930
rect 131920 678690 132160 678930
rect 132250 678690 132490 678930
rect 132580 678690 132820 678930
rect 132910 678690 133150 678930
rect 122190 678360 122430 678600
rect 122540 678360 122780 678600
rect 122870 678360 123110 678600
rect 123200 678360 123440 678600
rect 123530 678360 123770 678600
rect 123880 678360 124120 678600
rect 124210 678360 124450 678600
rect 124540 678360 124780 678600
rect 124870 678360 125110 678600
rect 125220 678360 125460 678600
rect 125550 678360 125790 678600
rect 125880 678360 126120 678600
rect 126210 678360 126450 678600
rect 126560 678360 126800 678600
rect 126890 678360 127130 678600
rect 127220 678360 127460 678600
rect 127550 678360 127790 678600
rect 127900 678360 128140 678600
rect 128230 678360 128470 678600
rect 128560 678360 128800 678600
rect 128890 678360 129130 678600
rect 129240 678360 129480 678600
rect 129570 678360 129810 678600
rect 129900 678360 130140 678600
rect 130230 678360 130470 678600
rect 130580 678360 130820 678600
rect 130910 678360 131150 678600
rect 131240 678360 131480 678600
rect 131570 678360 131810 678600
rect 131920 678360 132160 678600
rect 132250 678360 132490 678600
rect 132580 678360 132820 678600
rect 132910 678360 133150 678600
rect 122190 678030 122430 678270
rect 122540 678030 122780 678270
rect 122870 678030 123110 678270
rect 123200 678030 123440 678270
rect 123530 678030 123770 678270
rect 123880 678030 124120 678270
rect 124210 678030 124450 678270
rect 124540 678030 124780 678270
rect 124870 678030 125110 678270
rect 125220 678030 125460 678270
rect 125550 678030 125790 678270
rect 125880 678030 126120 678270
rect 126210 678030 126450 678270
rect 126560 678030 126800 678270
rect 126890 678030 127130 678270
rect 127220 678030 127460 678270
rect 127550 678030 127790 678270
rect 127900 678030 128140 678270
rect 128230 678030 128470 678270
rect 128560 678030 128800 678270
rect 128890 678030 129130 678270
rect 129240 678030 129480 678270
rect 129570 678030 129810 678270
rect 129900 678030 130140 678270
rect 130230 678030 130470 678270
rect 130580 678030 130820 678270
rect 130910 678030 131150 678270
rect 131240 678030 131480 678270
rect 131570 678030 131810 678270
rect 131920 678030 132160 678270
rect 132250 678030 132490 678270
rect 132580 678030 132820 678270
rect 132910 678030 133150 678270
rect 122190 677680 122430 677920
rect 122540 677680 122780 677920
rect 122870 677680 123110 677920
rect 123200 677680 123440 677920
rect 123530 677680 123770 677920
rect 123880 677680 124120 677920
rect 124210 677680 124450 677920
rect 124540 677680 124780 677920
rect 124870 677680 125110 677920
rect 125220 677680 125460 677920
rect 125550 677680 125790 677920
rect 125880 677680 126120 677920
rect 126210 677680 126450 677920
rect 126560 677680 126800 677920
rect 126890 677680 127130 677920
rect 127220 677680 127460 677920
rect 127550 677680 127790 677920
rect 127900 677680 128140 677920
rect 128230 677680 128470 677920
rect 128560 677680 128800 677920
rect 128890 677680 129130 677920
rect 129240 677680 129480 677920
rect 129570 677680 129810 677920
rect 129900 677680 130140 677920
rect 130230 677680 130470 677920
rect 130580 677680 130820 677920
rect 130910 677680 131150 677920
rect 131240 677680 131480 677920
rect 131570 677680 131810 677920
rect 131920 677680 132160 677920
rect 132250 677680 132490 677920
rect 132580 677680 132820 677920
rect 132910 677680 133150 677920
rect 122190 677350 122430 677590
rect 122540 677350 122780 677590
rect 122870 677350 123110 677590
rect 123200 677350 123440 677590
rect 123530 677350 123770 677590
rect 123880 677350 124120 677590
rect 124210 677350 124450 677590
rect 124540 677350 124780 677590
rect 124870 677350 125110 677590
rect 125220 677350 125460 677590
rect 125550 677350 125790 677590
rect 125880 677350 126120 677590
rect 126210 677350 126450 677590
rect 126560 677350 126800 677590
rect 126890 677350 127130 677590
rect 127220 677350 127460 677590
rect 127550 677350 127790 677590
rect 127900 677350 128140 677590
rect 128230 677350 128470 677590
rect 128560 677350 128800 677590
rect 128890 677350 129130 677590
rect 129240 677350 129480 677590
rect 129570 677350 129810 677590
rect 129900 677350 130140 677590
rect 130230 677350 130470 677590
rect 130580 677350 130820 677590
rect 130910 677350 131150 677590
rect 131240 677350 131480 677590
rect 131570 677350 131810 677590
rect 131920 677350 132160 677590
rect 132250 677350 132490 677590
rect 132580 677350 132820 677590
rect 132910 677350 133150 677590
rect 122190 677020 122430 677260
rect 122540 677020 122780 677260
rect 122870 677020 123110 677260
rect 123200 677020 123440 677260
rect 123530 677020 123770 677260
rect 123880 677020 124120 677260
rect 124210 677020 124450 677260
rect 124540 677020 124780 677260
rect 124870 677020 125110 677260
rect 125220 677020 125460 677260
rect 125550 677020 125790 677260
rect 125880 677020 126120 677260
rect 126210 677020 126450 677260
rect 126560 677020 126800 677260
rect 126890 677020 127130 677260
rect 127220 677020 127460 677260
rect 127550 677020 127790 677260
rect 127900 677020 128140 677260
rect 128230 677020 128470 677260
rect 128560 677020 128800 677260
rect 128890 677020 129130 677260
rect 129240 677020 129480 677260
rect 129570 677020 129810 677260
rect 129900 677020 130140 677260
rect 130230 677020 130470 677260
rect 130580 677020 130820 677260
rect 130910 677020 131150 677260
rect 131240 677020 131480 677260
rect 131570 677020 131810 677260
rect 131920 677020 132160 677260
rect 132250 677020 132490 677260
rect 132580 677020 132820 677260
rect 132910 677020 133150 677260
rect 122190 676690 122430 676930
rect 122540 676690 122780 676930
rect 122870 676690 123110 676930
rect 123200 676690 123440 676930
rect 123530 676690 123770 676930
rect 123880 676690 124120 676930
rect 124210 676690 124450 676930
rect 124540 676690 124780 676930
rect 124870 676690 125110 676930
rect 125220 676690 125460 676930
rect 125550 676690 125790 676930
rect 125880 676690 126120 676930
rect 126210 676690 126450 676930
rect 126560 676690 126800 676930
rect 126890 676690 127130 676930
rect 127220 676690 127460 676930
rect 127550 676690 127790 676930
rect 127900 676690 128140 676930
rect 128230 676690 128470 676930
rect 128560 676690 128800 676930
rect 128890 676690 129130 676930
rect 129240 676690 129480 676930
rect 129570 676690 129810 676930
rect 129900 676690 130140 676930
rect 130230 676690 130470 676930
rect 130580 676690 130820 676930
rect 130910 676690 131150 676930
rect 131240 676690 131480 676930
rect 131570 676690 131810 676930
rect 131920 676690 132160 676930
rect 132250 676690 132490 676930
rect 132580 676690 132820 676930
rect 132910 676690 133150 676930
rect 122190 676340 122430 676580
rect 122540 676340 122780 676580
rect 122870 676340 123110 676580
rect 123200 676340 123440 676580
rect 123530 676340 123770 676580
rect 123880 676340 124120 676580
rect 124210 676340 124450 676580
rect 124540 676340 124780 676580
rect 124870 676340 125110 676580
rect 125220 676340 125460 676580
rect 125550 676340 125790 676580
rect 125880 676340 126120 676580
rect 126210 676340 126450 676580
rect 126560 676340 126800 676580
rect 126890 676340 127130 676580
rect 127220 676340 127460 676580
rect 127550 676340 127790 676580
rect 127900 676340 128140 676580
rect 128230 676340 128470 676580
rect 128560 676340 128800 676580
rect 128890 676340 129130 676580
rect 129240 676340 129480 676580
rect 129570 676340 129810 676580
rect 129900 676340 130140 676580
rect 130230 676340 130470 676580
rect 130580 676340 130820 676580
rect 130910 676340 131150 676580
rect 131240 676340 131480 676580
rect 131570 676340 131810 676580
rect 131920 676340 132160 676580
rect 132250 676340 132490 676580
rect 132580 676340 132820 676580
rect 132910 676340 133150 676580
rect 122190 676010 122430 676250
rect 122540 676010 122780 676250
rect 122870 676010 123110 676250
rect 123200 676010 123440 676250
rect 123530 676010 123770 676250
rect 123880 676010 124120 676250
rect 124210 676010 124450 676250
rect 124540 676010 124780 676250
rect 124870 676010 125110 676250
rect 125220 676010 125460 676250
rect 125550 676010 125790 676250
rect 125880 676010 126120 676250
rect 126210 676010 126450 676250
rect 126560 676010 126800 676250
rect 126890 676010 127130 676250
rect 127220 676010 127460 676250
rect 127550 676010 127790 676250
rect 127900 676010 128140 676250
rect 128230 676010 128470 676250
rect 128560 676010 128800 676250
rect 128890 676010 129130 676250
rect 129240 676010 129480 676250
rect 129570 676010 129810 676250
rect 129900 676010 130140 676250
rect 130230 676010 130470 676250
rect 130580 676010 130820 676250
rect 130910 676010 131150 676250
rect 131240 676010 131480 676250
rect 131570 676010 131810 676250
rect 131920 676010 132160 676250
rect 132250 676010 132490 676250
rect 132580 676010 132820 676250
rect 132910 676010 133150 676250
rect 122190 675680 122430 675920
rect 122540 675680 122780 675920
rect 122870 675680 123110 675920
rect 123200 675680 123440 675920
rect 123530 675680 123770 675920
rect 123880 675680 124120 675920
rect 124210 675680 124450 675920
rect 124540 675680 124780 675920
rect 124870 675680 125110 675920
rect 125220 675680 125460 675920
rect 125550 675680 125790 675920
rect 125880 675680 126120 675920
rect 126210 675680 126450 675920
rect 126560 675680 126800 675920
rect 126890 675680 127130 675920
rect 127220 675680 127460 675920
rect 127550 675680 127790 675920
rect 127900 675680 128140 675920
rect 128230 675680 128470 675920
rect 128560 675680 128800 675920
rect 128890 675680 129130 675920
rect 129240 675680 129480 675920
rect 129570 675680 129810 675920
rect 129900 675680 130140 675920
rect 130230 675680 130470 675920
rect 130580 675680 130820 675920
rect 130910 675680 131150 675920
rect 131240 675680 131480 675920
rect 131570 675680 131810 675920
rect 131920 675680 132160 675920
rect 132250 675680 132490 675920
rect 132580 675680 132820 675920
rect 132910 675680 133150 675920
rect 122190 675350 122430 675590
rect 122540 675350 122780 675590
rect 122870 675350 123110 675590
rect 123200 675350 123440 675590
rect 123530 675350 123770 675590
rect 123880 675350 124120 675590
rect 124210 675350 124450 675590
rect 124540 675350 124780 675590
rect 124870 675350 125110 675590
rect 125220 675350 125460 675590
rect 125550 675350 125790 675590
rect 125880 675350 126120 675590
rect 126210 675350 126450 675590
rect 126560 675350 126800 675590
rect 126890 675350 127130 675590
rect 127220 675350 127460 675590
rect 127550 675350 127790 675590
rect 127900 675350 128140 675590
rect 128230 675350 128470 675590
rect 128560 675350 128800 675590
rect 128890 675350 129130 675590
rect 129240 675350 129480 675590
rect 129570 675350 129810 675590
rect 129900 675350 130140 675590
rect 130230 675350 130470 675590
rect 130580 675350 130820 675590
rect 130910 675350 131150 675590
rect 131240 675350 131480 675590
rect 131570 675350 131810 675590
rect 131920 675350 132160 675590
rect 132250 675350 132490 675590
rect 132580 675350 132820 675590
rect 132910 675350 133150 675590
rect 122190 675000 122430 675240
rect 122540 675000 122780 675240
rect 122870 675000 123110 675240
rect 123200 675000 123440 675240
rect 123530 675000 123770 675240
rect 123880 675000 124120 675240
rect 124210 675000 124450 675240
rect 124540 675000 124780 675240
rect 124870 675000 125110 675240
rect 125220 675000 125460 675240
rect 125550 675000 125790 675240
rect 125880 675000 126120 675240
rect 126210 675000 126450 675240
rect 126560 675000 126800 675240
rect 126890 675000 127130 675240
rect 127220 675000 127460 675240
rect 127550 675000 127790 675240
rect 127900 675000 128140 675240
rect 128230 675000 128470 675240
rect 128560 675000 128800 675240
rect 128890 675000 129130 675240
rect 129240 675000 129480 675240
rect 129570 675000 129810 675240
rect 129900 675000 130140 675240
rect 130230 675000 130470 675240
rect 130580 675000 130820 675240
rect 130910 675000 131150 675240
rect 131240 675000 131480 675240
rect 131570 675000 131810 675240
rect 131920 675000 132160 675240
rect 132250 675000 132490 675240
rect 132580 675000 132820 675240
rect 132910 675000 133150 675240
rect 122190 674670 122430 674910
rect 122540 674670 122780 674910
rect 122870 674670 123110 674910
rect 123200 674670 123440 674910
rect 123530 674670 123770 674910
rect 123880 674670 124120 674910
rect 124210 674670 124450 674910
rect 124540 674670 124780 674910
rect 124870 674670 125110 674910
rect 125220 674670 125460 674910
rect 125550 674670 125790 674910
rect 125880 674670 126120 674910
rect 126210 674670 126450 674910
rect 126560 674670 126800 674910
rect 126890 674670 127130 674910
rect 127220 674670 127460 674910
rect 127550 674670 127790 674910
rect 127900 674670 128140 674910
rect 128230 674670 128470 674910
rect 128560 674670 128800 674910
rect 128890 674670 129130 674910
rect 129240 674670 129480 674910
rect 129570 674670 129810 674910
rect 129900 674670 130140 674910
rect 130230 674670 130470 674910
rect 130580 674670 130820 674910
rect 130910 674670 131150 674910
rect 131240 674670 131480 674910
rect 131570 674670 131810 674910
rect 131920 674670 132160 674910
rect 132250 674670 132490 674910
rect 132580 674670 132820 674910
rect 132910 674670 133150 674910
rect 122190 674340 122430 674580
rect 122540 674340 122780 674580
rect 122870 674340 123110 674580
rect 123200 674340 123440 674580
rect 123530 674340 123770 674580
rect 123880 674340 124120 674580
rect 124210 674340 124450 674580
rect 124540 674340 124780 674580
rect 124870 674340 125110 674580
rect 125220 674340 125460 674580
rect 125550 674340 125790 674580
rect 125880 674340 126120 674580
rect 126210 674340 126450 674580
rect 126560 674340 126800 674580
rect 126890 674340 127130 674580
rect 127220 674340 127460 674580
rect 127550 674340 127790 674580
rect 127900 674340 128140 674580
rect 128230 674340 128470 674580
rect 128560 674340 128800 674580
rect 128890 674340 129130 674580
rect 129240 674340 129480 674580
rect 129570 674340 129810 674580
rect 129900 674340 130140 674580
rect 130230 674340 130470 674580
rect 130580 674340 130820 674580
rect 130910 674340 131150 674580
rect 131240 674340 131480 674580
rect 131570 674340 131810 674580
rect 131920 674340 132160 674580
rect 132250 674340 132490 674580
rect 132580 674340 132820 674580
rect 132910 674340 133150 674580
rect 122190 674010 122430 674250
rect 122540 674010 122780 674250
rect 122870 674010 123110 674250
rect 123200 674010 123440 674250
rect 123530 674010 123770 674250
rect 123880 674010 124120 674250
rect 124210 674010 124450 674250
rect 124540 674010 124780 674250
rect 124870 674010 125110 674250
rect 125220 674010 125460 674250
rect 125550 674010 125790 674250
rect 125880 674010 126120 674250
rect 126210 674010 126450 674250
rect 126560 674010 126800 674250
rect 126890 674010 127130 674250
rect 127220 674010 127460 674250
rect 127550 674010 127790 674250
rect 127900 674010 128140 674250
rect 128230 674010 128470 674250
rect 128560 674010 128800 674250
rect 128890 674010 129130 674250
rect 129240 674010 129480 674250
rect 129570 674010 129810 674250
rect 129900 674010 130140 674250
rect 130230 674010 130470 674250
rect 130580 674010 130820 674250
rect 130910 674010 131150 674250
rect 131240 674010 131480 674250
rect 131570 674010 131810 674250
rect 131920 674010 132160 674250
rect 132250 674010 132490 674250
rect 132580 674010 132820 674250
rect 132910 674010 133150 674250
rect 122190 673660 122430 673900
rect 122540 673660 122780 673900
rect 122870 673660 123110 673900
rect 123200 673660 123440 673900
rect 123530 673660 123770 673900
rect 123880 673660 124120 673900
rect 124210 673660 124450 673900
rect 124540 673660 124780 673900
rect 124870 673660 125110 673900
rect 125220 673660 125460 673900
rect 125550 673660 125790 673900
rect 125880 673660 126120 673900
rect 126210 673660 126450 673900
rect 126560 673660 126800 673900
rect 126890 673660 127130 673900
rect 127220 673660 127460 673900
rect 127550 673660 127790 673900
rect 127900 673660 128140 673900
rect 128230 673660 128470 673900
rect 128560 673660 128800 673900
rect 128890 673660 129130 673900
rect 129240 673660 129480 673900
rect 129570 673660 129810 673900
rect 129900 673660 130140 673900
rect 130230 673660 130470 673900
rect 130580 673660 130820 673900
rect 130910 673660 131150 673900
rect 131240 673660 131480 673900
rect 131570 673660 131810 673900
rect 131920 673660 132160 673900
rect 132250 673660 132490 673900
rect 132580 673660 132820 673900
rect 132910 673660 133150 673900
rect 122190 673330 122430 673570
rect 122540 673330 122780 673570
rect 122870 673330 123110 673570
rect 123200 673330 123440 673570
rect 123530 673330 123770 673570
rect 123880 673330 124120 673570
rect 124210 673330 124450 673570
rect 124540 673330 124780 673570
rect 124870 673330 125110 673570
rect 125220 673330 125460 673570
rect 125550 673330 125790 673570
rect 125880 673330 126120 673570
rect 126210 673330 126450 673570
rect 126560 673330 126800 673570
rect 126890 673330 127130 673570
rect 127220 673330 127460 673570
rect 127550 673330 127790 673570
rect 127900 673330 128140 673570
rect 128230 673330 128470 673570
rect 128560 673330 128800 673570
rect 128890 673330 129130 673570
rect 129240 673330 129480 673570
rect 129570 673330 129810 673570
rect 129900 673330 130140 673570
rect 130230 673330 130470 673570
rect 130580 673330 130820 673570
rect 130910 673330 131150 673570
rect 131240 673330 131480 673570
rect 131570 673330 131810 673570
rect 131920 673330 132160 673570
rect 132250 673330 132490 673570
rect 132580 673330 132820 673570
rect 132910 673330 133150 673570
rect 122190 673000 122430 673240
rect 122540 673000 122780 673240
rect 122870 673000 123110 673240
rect 123200 673000 123440 673240
rect 123530 673000 123770 673240
rect 123880 673000 124120 673240
rect 124210 673000 124450 673240
rect 124540 673000 124780 673240
rect 124870 673000 125110 673240
rect 125220 673000 125460 673240
rect 125550 673000 125790 673240
rect 125880 673000 126120 673240
rect 126210 673000 126450 673240
rect 126560 673000 126800 673240
rect 126890 673000 127130 673240
rect 127220 673000 127460 673240
rect 127550 673000 127790 673240
rect 127900 673000 128140 673240
rect 128230 673000 128470 673240
rect 128560 673000 128800 673240
rect 128890 673000 129130 673240
rect 129240 673000 129480 673240
rect 129570 673000 129810 673240
rect 129900 673000 130140 673240
rect 130230 673000 130470 673240
rect 130580 673000 130820 673240
rect 130910 673000 131150 673240
rect 131240 673000 131480 673240
rect 131570 673000 131810 673240
rect 131920 673000 132160 673240
rect 132250 673000 132490 673240
rect 132580 673000 132820 673240
rect 132910 673000 133150 673240
rect 122190 672670 122430 672910
rect 122540 672670 122780 672910
rect 122870 672670 123110 672910
rect 123200 672670 123440 672910
rect 123530 672670 123770 672910
rect 123880 672670 124120 672910
rect 124210 672670 124450 672910
rect 124540 672670 124780 672910
rect 124870 672670 125110 672910
rect 125220 672670 125460 672910
rect 125550 672670 125790 672910
rect 125880 672670 126120 672910
rect 126210 672670 126450 672910
rect 126560 672670 126800 672910
rect 126890 672670 127130 672910
rect 127220 672670 127460 672910
rect 127550 672670 127790 672910
rect 127900 672670 128140 672910
rect 128230 672670 128470 672910
rect 128560 672670 128800 672910
rect 128890 672670 129130 672910
rect 129240 672670 129480 672910
rect 129570 672670 129810 672910
rect 129900 672670 130140 672910
rect 130230 672670 130470 672910
rect 130580 672670 130820 672910
rect 130910 672670 131150 672910
rect 131240 672670 131480 672910
rect 131570 672670 131810 672910
rect 131920 672670 132160 672910
rect 132250 672670 132490 672910
rect 132580 672670 132820 672910
rect 132910 672670 133150 672910
rect 122190 672320 122430 672560
rect 122540 672320 122780 672560
rect 122870 672320 123110 672560
rect 123200 672320 123440 672560
rect 123530 672320 123770 672560
rect 123880 672320 124120 672560
rect 124210 672320 124450 672560
rect 124540 672320 124780 672560
rect 124870 672320 125110 672560
rect 125220 672320 125460 672560
rect 125550 672320 125790 672560
rect 125880 672320 126120 672560
rect 126210 672320 126450 672560
rect 126560 672320 126800 672560
rect 126890 672320 127130 672560
rect 127220 672320 127460 672560
rect 127550 672320 127790 672560
rect 127900 672320 128140 672560
rect 128230 672320 128470 672560
rect 128560 672320 128800 672560
rect 128890 672320 129130 672560
rect 129240 672320 129480 672560
rect 129570 672320 129810 672560
rect 129900 672320 130140 672560
rect 130230 672320 130470 672560
rect 130580 672320 130820 672560
rect 130910 672320 131150 672560
rect 131240 672320 131480 672560
rect 131570 672320 131810 672560
rect 131920 672320 132160 672560
rect 132250 672320 132490 672560
rect 132580 672320 132820 672560
rect 132910 672320 133150 672560
rect 133570 683040 133810 683280
rect 133920 683040 134160 683280
rect 134250 683040 134490 683280
rect 134580 683040 134820 683280
rect 134910 683040 135150 683280
rect 135260 683040 135500 683280
rect 135590 683040 135830 683280
rect 135920 683040 136160 683280
rect 136250 683040 136490 683280
rect 136600 683040 136840 683280
rect 136930 683040 137170 683280
rect 137260 683040 137500 683280
rect 137590 683040 137830 683280
rect 137940 683040 138180 683280
rect 138270 683040 138510 683280
rect 138600 683040 138840 683280
rect 138930 683040 139170 683280
rect 139280 683040 139520 683280
rect 139610 683040 139850 683280
rect 139940 683040 140180 683280
rect 140270 683040 140510 683280
rect 140620 683040 140860 683280
rect 140950 683040 141190 683280
rect 141280 683040 141520 683280
rect 141610 683040 141850 683280
rect 141960 683040 142200 683280
rect 142290 683040 142530 683280
rect 142620 683040 142860 683280
rect 142950 683040 143190 683280
rect 143300 683040 143540 683280
rect 143630 683040 143870 683280
rect 143960 683040 144200 683280
rect 144290 683040 144530 683280
rect 133570 682710 133810 682950
rect 133920 682710 134160 682950
rect 134250 682710 134490 682950
rect 134580 682710 134820 682950
rect 134910 682710 135150 682950
rect 135260 682710 135500 682950
rect 135590 682710 135830 682950
rect 135920 682710 136160 682950
rect 136250 682710 136490 682950
rect 136600 682710 136840 682950
rect 136930 682710 137170 682950
rect 137260 682710 137500 682950
rect 137590 682710 137830 682950
rect 137940 682710 138180 682950
rect 138270 682710 138510 682950
rect 138600 682710 138840 682950
rect 138930 682710 139170 682950
rect 139280 682710 139520 682950
rect 139610 682710 139850 682950
rect 139940 682710 140180 682950
rect 140270 682710 140510 682950
rect 140620 682710 140860 682950
rect 140950 682710 141190 682950
rect 141280 682710 141520 682950
rect 141610 682710 141850 682950
rect 141960 682710 142200 682950
rect 142290 682710 142530 682950
rect 142620 682710 142860 682950
rect 142950 682710 143190 682950
rect 143300 682710 143540 682950
rect 143630 682710 143870 682950
rect 143960 682710 144200 682950
rect 144290 682710 144530 682950
rect 133570 682380 133810 682620
rect 133920 682380 134160 682620
rect 134250 682380 134490 682620
rect 134580 682380 134820 682620
rect 134910 682380 135150 682620
rect 135260 682380 135500 682620
rect 135590 682380 135830 682620
rect 135920 682380 136160 682620
rect 136250 682380 136490 682620
rect 136600 682380 136840 682620
rect 136930 682380 137170 682620
rect 137260 682380 137500 682620
rect 137590 682380 137830 682620
rect 137940 682380 138180 682620
rect 138270 682380 138510 682620
rect 138600 682380 138840 682620
rect 138930 682380 139170 682620
rect 139280 682380 139520 682620
rect 139610 682380 139850 682620
rect 139940 682380 140180 682620
rect 140270 682380 140510 682620
rect 140620 682380 140860 682620
rect 140950 682380 141190 682620
rect 141280 682380 141520 682620
rect 141610 682380 141850 682620
rect 141960 682380 142200 682620
rect 142290 682380 142530 682620
rect 142620 682380 142860 682620
rect 142950 682380 143190 682620
rect 143300 682380 143540 682620
rect 143630 682380 143870 682620
rect 143960 682380 144200 682620
rect 144290 682380 144530 682620
rect 133570 682050 133810 682290
rect 133920 682050 134160 682290
rect 134250 682050 134490 682290
rect 134580 682050 134820 682290
rect 134910 682050 135150 682290
rect 135260 682050 135500 682290
rect 135590 682050 135830 682290
rect 135920 682050 136160 682290
rect 136250 682050 136490 682290
rect 136600 682050 136840 682290
rect 136930 682050 137170 682290
rect 137260 682050 137500 682290
rect 137590 682050 137830 682290
rect 137940 682050 138180 682290
rect 138270 682050 138510 682290
rect 138600 682050 138840 682290
rect 138930 682050 139170 682290
rect 139280 682050 139520 682290
rect 139610 682050 139850 682290
rect 139940 682050 140180 682290
rect 140270 682050 140510 682290
rect 140620 682050 140860 682290
rect 140950 682050 141190 682290
rect 141280 682050 141520 682290
rect 141610 682050 141850 682290
rect 141960 682050 142200 682290
rect 142290 682050 142530 682290
rect 142620 682050 142860 682290
rect 142950 682050 143190 682290
rect 143300 682050 143540 682290
rect 143630 682050 143870 682290
rect 143960 682050 144200 682290
rect 144290 682050 144530 682290
rect 133570 681700 133810 681940
rect 133920 681700 134160 681940
rect 134250 681700 134490 681940
rect 134580 681700 134820 681940
rect 134910 681700 135150 681940
rect 135260 681700 135500 681940
rect 135590 681700 135830 681940
rect 135920 681700 136160 681940
rect 136250 681700 136490 681940
rect 136600 681700 136840 681940
rect 136930 681700 137170 681940
rect 137260 681700 137500 681940
rect 137590 681700 137830 681940
rect 137940 681700 138180 681940
rect 138270 681700 138510 681940
rect 138600 681700 138840 681940
rect 138930 681700 139170 681940
rect 139280 681700 139520 681940
rect 139610 681700 139850 681940
rect 139940 681700 140180 681940
rect 140270 681700 140510 681940
rect 140620 681700 140860 681940
rect 140950 681700 141190 681940
rect 141280 681700 141520 681940
rect 141610 681700 141850 681940
rect 141960 681700 142200 681940
rect 142290 681700 142530 681940
rect 142620 681700 142860 681940
rect 142950 681700 143190 681940
rect 143300 681700 143540 681940
rect 143630 681700 143870 681940
rect 143960 681700 144200 681940
rect 144290 681700 144530 681940
rect 133570 681370 133810 681610
rect 133920 681370 134160 681610
rect 134250 681370 134490 681610
rect 134580 681370 134820 681610
rect 134910 681370 135150 681610
rect 135260 681370 135500 681610
rect 135590 681370 135830 681610
rect 135920 681370 136160 681610
rect 136250 681370 136490 681610
rect 136600 681370 136840 681610
rect 136930 681370 137170 681610
rect 137260 681370 137500 681610
rect 137590 681370 137830 681610
rect 137940 681370 138180 681610
rect 138270 681370 138510 681610
rect 138600 681370 138840 681610
rect 138930 681370 139170 681610
rect 139280 681370 139520 681610
rect 139610 681370 139850 681610
rect 139940 681370 140180 681610
rect 140270 681370 140510 681610
rect 140620 681370 140860 681610
rect 140950 681370 141190 681610
rect 141280 681370 141520 681610
rect 141610 681370 141850 681610
rect 141960 681370 142200 681610
rect 142290 681370 142530 681610
rect 142620 681370 142860 681610
rect 142950 681370 143190 681610
rect 143300 681370 143540 681610
rect 143630 681370 143870 681610
rect 143960 681370 144200 681610
rect 144290 681370 144530 681610
rect 133570 681040 133810 681280
rect 133920 681040 134160 681280
rect 134250 681040 134490 681280
rect 134580 681040 134820 681280
rect 134910 681040 135150 681280
rect 135260 681040 135500 681280
rect 135590 681040 135830 681280
rect 135920 681040 136160 681280
rect 136250 681040 136490 681280
rect 136600 681040 136840 681280
rect 136930 681040 137170 681280
rect 137260 681040 137500 681280
rect 137590 681040 137830 681280
rect 137940 681040 138180 681280
rect 138270 681040 138510 681280
rect 138600 681040 138840 681280
rect 138930 681040 139170 681280
rect 139280 681040 139520 681280
rect 139610 681040 139850 681280
rect 139940 681040 140180 681280
rect 140270 681040 140510 681280
rect 140620 681040 140860 681280
rect 140950 681040 141190 681280
rect 141280 681040 141520 681280
rect 141610 681040 141850 681280
rect 141960 681040 142200 681280
rect 142290 681040 142530 681280
rect 142620 681040 142860 681280
rect 142950 681040 143190 681280
rect 143300 681040 143540 681280
rect 143630 681040 143870 681280
rect 143960 681040 144200 681280
rect 144290 681040 144530 681280
rect 133570 680710 133810 680950
rect 133920 680710 134160 680950
rect 134250 680710 134490 680950
rect 134580 680710 134820 680950
rect 134910 680710 135150 680950
rect 135260 680710 135500 680950
rect 135590 680710 135830 680950
rect 135920 680710 136160 680950
rect 136250 680710 136490 680950
rect 136600 680710 136840 680950
rect 136930 680710 137170 680950
rect 137260 680710 137500 680950
rect 137590 680710 137830 680950
rect 137940 680710 138180 680950
rect 138270 680710 138510 680950
rect 138600 680710 138840 680950
rect 138930 680710 139170 680950
rect 139280 680710 139520 680950
rect 139610 680710 139850 680950
rect 139940 680710 140180 680950
rect 140270 680710 140510 680950
rect 140620 680710 140860 680950
rect 140950 680710 141190 680950
rect 141280 680710 141520 680950
rect 141610 680710 141850 680950
rect 141960 680710 142200 680950
rect 142290 680710 142530 680950
rect 142620 680710 142860 680950
rect 142950 680710 143190 680950
rect 143300 680710 143540 680950
rect 143630 680710 143870 680950
rect 143960 680710 144200 680950
rect 144290 680710 144530 680950
rect 133570 680360 133810 680600
rect 133920 680360 134160 680600
rect 134250 680360 134490 680600
rect 134580 680360 134820 680600
rect 134910 680360 135150 680600
rect 135260 680360 135500 680600
rect 135590 680360 135830 680600
rect 135920 680360 136160 680600
rect 136250 680360 136490 680600
rect 136600 680360 136840 680600
rect 136930 680360 137170 680600
rect 137260 680360 137500 680600
rect 137590 680360 137830 680600
rect 137940 680360 138180 680600
rect 138270 680360 138510 680600
rect 138600 680360 138840 680600
rect 138930 680360 139170 680600
rect 139280 680360 139520 680600
rect 139610 680360 139850 680600
rect 139940 680360 140180 680600
rect 140270 680360 140510 680600
rect 140620 680360 140860 680600
rect 140950 680360 141190 680600
rect 141280 680360 141520 680600
rect 141610 680360 141850 680600
rect 141960 680360 142200 680600
rect 142290 680360 142530 680600
rect 142620 680360 142860 680600
rect 142950 680360 143190 680600
rect 143300 680360 143540 680600
rect 143630 680360 143870 680600
rect 143960 680360 144200 680600
rect 144290 680360 144530 680600
rect 133570 680030 133810 680270
rect 133920 680030 134160 680270
rect 134250 680030 134490 680270
rect 134580 680030 134820 680270
rect 134910 680030 135150 680270
rect 135260 680030 135500 680270
rect 135590 680030 135830 680270
rect 135920 680030 136160 680270
rect 136250 680030 136490 680270
rect 136600 680030 136840 680270
rect 136930 680030 137170 680270
rect 137260 680030 137500 680270
rect 137590 680030 137830 680270
rect 137940 680030 138180 680270
rect 138270 680030 138510 680270
rect 138600 680030 138840 680270
rect 138930 680030 139170 680270
rect 139280 680030 139520 680270
rect 139610 680030 139850 680270
rect 139940 680030 140180 680270
rect 140270 680030 140510 680270
rect 140620 680030 140860 680270
rect 140950 680030 141190 680270
rect 141280 680030 141520 680270
rect 141610 680030 141850 680270
rect 141960 680030 142200 680270
rect 142290 680030 142530 680270
rect 142620 680030 142860 680270
rect 142950 680030 143190 680270
rect 143300 680030 143540 680270
rect 143630 680030 143870 680270
rect 143960 680030 144200 680270
rect 144290 680030 144530 680270
rect 133570 679700 133810 679940
rect 133920 679700 134160 679940
rect 134250 679700 134490 679940
rect 134580 679700 134820 679940
rect 134910 679700 135150 679940
rect 135260 679700 135500 679940
rect 135590 679700 135830 679940
rect 135920 679700 136160 679940
rect 136250 679700 136490 679940
rect 136600 679700 136840 679940
rect 136930 679700 137170 679940
rect 137260 679700 137500 679940
rect 137590 679700 137830 679940
rect 137940 679700 138180 679940
rect 138270 679700 138510 679940
rect 138600 679700 138840 679940
rect 138930 679700 139170 679940
rect 139280 679700 139520 679940
rect 139610 679700 139850 679940
rect 139940 679700 140180 679940
rect 140270 679700 140510 679940
rect 140620 679700 140860 679940
rect 140950 679700 141190 679940
rect 141280 679700 141520 679940
rect 141610 679700 141850 679940
rect 141960 679700 142200 679940
rect 142290 679700 142530 679940
rect 142620 679700 142860 679940
rect 142950 679700 143190 679940
rect 143300 679700 143540 679940
rect 143630 679700 143870 679940
rect 143960 679700 144200 679940
rect 144290 679700 144530 679940
rect 133570 679370 133810 679610
rect 133920 679370 134160 679610
rect 134250 679370 134490 679610
rect 134580 679370 134820 679610
rect 134910 679370 135150 679610
rect 135260 679370 135500 679610
rect 135590 679370 135830 679610
rect 135920 679370 136160 679610
rect 136250 679370 136490 679610
rect 136600 679370 136840 679610
rect 136930 679370 137170 679610
rect 137260 679370 137500 679610
rect 137590 679370 137830 679610
rect 137940 679370 138180 679610
rect 138270 679370 138510 679610
rect 138600 679370 138840 679610
rect 138930 679370 139170 679610
rect 139280 679370 139520 679610
rect 139610 679370 139850 679610
rect 139940 679370 140180 679610
rect 140270 679370 140510 679610
rect 140620 679370 140860 679610
rect 140950 679370 141190 679610
rect 141280 679370 141520 679610
rect 141610 679370 141850 679610
rect 141960 679370 142200 679610
rect 142290 679370 142530 679610
rect 142620 679370 142860 679610
rect 142950 679370 143190 679610
rect 143300 679370 143540 679610
rect 143630 679370 143870 679610
rect 143960 679370 144200 679610
rect 144290 679370 144530 679610
rect 133570 679020 133810 679260
rect 133920 679020 134160 679260
rect 134250 679020 134490 679260
rect 134580 679020 134820 679260
rect 134910 679020 135150 679260
rect 135260 679020 135500 679260
rect 135590 679020 135830 679260
rect 135920 679020 136160 679260
rect 136250 679020 136490 679260
rect 136600 679020 136840 679260
rect 136930 679020 137170 679260
rect 137260 679020 137500 679260
rect 137590 679020 137830 679260
rect 137940 679020 138180 679260
rect 138270 679020 138510 679260
rect 138600 679020 138840 679260
rect 138930 679020 139170 679260
rect 139280 679020 139520 679260
rect 139610 679020 139850 679260
rect 139940 679020 140180 679260
rect 140270 679020 140510 679260
rect 140620 679020 140860 679260
rect 140950 679020 141190 679260
rect 141280 679020 141520 679260
rect 141610 679020 141850 679260
rect 141960 679020 142200 679260
rect 142290 679020 142530 679260
rect 142620 679020 142860 679260
rect 142950 679020 143190 679260
rect 143300 679020 143540 679260
rect 143630 679020 143870 679260
rect 143960 679020 144200 679260
rect 144290 679020 144530 679260
rect 133570 678690 133810 678930
rect 133920 678690 134160 678930
rect 134250 678690 134490 678930
rect 134580 678690 134820 678930
rect 134910 678690 135150 678930
rect 135260 678690 135500 678930
rect 135590 678690 135830 678930
rect 135920 678690 136160 678930
rect 136250 678690 136490 678930
rect 136600 678690 136840 678930
rect 136930 678690 137170 678930
rect 137260 678690 137500 678930
rect 137590 678690 137830 678930
rect 137940 678690 138180 678930
rect 138270 678690 138510 678930
rect 138600 678690 138840 678930
rect 138930 678690 139170 678930
rect 139280 678690 139520 678930
rect 139610 678690 139850 678930
rect 139940 678690 140180 678930
rect 140270 678690 140510 678930
rect 140620 678690 140860 678930
rect 140950 678690 141190 678930
rect 141280 678690 141520 678930
rect 141610 678690 141850 678930
rect 141960 678690 142200 678930
rect 142290 678690 142530 678930
rect 142620 678690 142860 678930
rect 142950 678690 143190 678930
rect 143300 678690 143540 678930
rect 143630 678690 143870 678930
rect 143960 678690 144200 678930
rect 144290 678690 144530 678930
rect 133570 678360 133810 678600
rect 133920 678360 134160 678600
rect 134250 678360 134490 678600
rect 134580 678360 134820 678600
rect 134910 678360 135150 678600
rect 135260 678360 135500 678600
rect 135590 678360 135830 678600
rect 135920 678360 136160 678600
rect 136250 678360 136490 678600
rect 136600 678360 136840 678600
rect 136930 678360 137170 678600
rect 137260 678360 137500 678600
rect 137590 678360 137830 678600
rect 137940 678360 138180 678600
rect 138270 678360 138510 678600
rect 138600 678360 138840 678600
rect 138930 678360 139170 678600
rect 139280 678360 139520 678600
rect 139610 678360 139850 678600
rect 139940 678360 140180 678600
rect 140270 678360 140510 678600
rect 140620 678360 140860 678600
rect 140950 678360 141190 678600
rect 141280 678360 141520 678600
rect 141610 678360 141850 678600
rect 141960 678360 142200 678600
rect 142290 678360 142530 678600
rect 142620 678360 142860 678600
rect 142950 678360 143190 678600
rect 143300 678360 143540 678600
rect 143630 678360 143870 678600
rect 143960 678360 144200 678600
rect 144290 678360 144530 678600
rect 133570 678030 133810 678270
rect 133920 678030 134160 678270
rect 134250 678030 134490 678270
rect 134580 678030 134820 678270
rect 134910 678030 135150 678270
rect 135260 678030 135500 678270
rect 135590 678030 135830 678270
rect 135920 678030 136160 678270
rect 136250 678030 136490 678270
rect 136600 678030 136840 678270
rect 136930 678030 137170 678270
rect 137260 678030 137500 678270
rect 137590 678030 137830 678270
rect 137940 678030 138180 678270
rect 138270 678030 138510 678270
rect 138600 678030 138840 678270
rect 138930 678030 139170 678270
rect 139280 678030 139520 678270
rect 139610 678030 139850 678270
rect 139940 678030 140180 678270
rect 140270 678030 140510 678270
rect 140620 678030 140860 678270
rect 140950 678030 141190 678270
rect 141280 678030 141520 678270
rect 141610 678030 141850 678270
rect 141960 678030 142200 678270
rect 142290 678030 142530 678270
rect 142620 678030 142860 678270
rect 142950 678030 143190 678270
rect 143300 678030 143540 678270
rect 143630 678030 143870 678270
rect 143960 678030 144200 678270
rect 144290 678030 144530 678270
rect 133570 677680 133810 677920
rect 133920 677680 134160 677920
rect 134250 677680 134490 677920
rect 134580 677680 134820 677920
rect 134910 677680 135150 677920
rect 135260 677680 135500 677920
rect 135590 677680 135830 677920
rect 135920 677680 136160 677920
rect 136250 677680 136490 677920
rect 136600 677680 136840 677920
rect 136930 677680 137170 677920
rect 137260 677680 137500 677920
rect 137590 677680 137830 677920
rect 137940 677680 138180 677920
rect 138270 677680 138510 677920
rect 138600 677680 138840 677920
rect 138930 677680 139170 677920
rect 139280 677680 139520 677920
rect 139610 677680 139850 677920
rect 139940 677680 140180 677920
rect 140270 677680 140510 677920
rect 140620 677680 140860 677920
rect 140950 677680 141190 677920
rect 141280 677680 141520 677920
rect 141610 677680 141850 677920
rect 141960 677680 142200 677920
rect 142290 677680 142530 677920
rect 142620 677680 142860 677920
rect 142950 677680 143190 677920
rect 143300 677680 143540 677920
rect 143630 677680 143870 677920
rect 143960 677680 144200 677920
rect 144290 677680 144530 677920
rect 133570 677350 133810 677590
rect 133920 677350 134160 677590
rect 134250 677350 134490 677590
rect 134580 677350 134820 677590
rect 134910 677350 135150 677590
rect 135260 677350 135500 677590
rect 135590 677350 135830 677590
rect 135920 677350 136160 677590
rect 136250 677350 136490 677590
rect 136600 677350 136840 677590
rect 136930 677350 137170 677590
rect 137260 677350 137500 677590
rect 137590 677350 137830 677590
rect 137940 677350 138180 677590
rect 138270 677350 138510 677590
rect 138600 677350 138840 677590
rect 138930 677350 139170 677590
rect 139280 677350 139520 677590
rect 139610 677350 139850 677590
rect 139940 677350 140180 677590
rect 140270 677350 140510 677590
rect 140620 677350 140860 677590
rect 140950 677350 141190 677590
rect 141280 677350 141520 677590
rect 141610 677350 141850 677590
rect 141960 677350 142200 677590
rect 142290 677350 142530 677590
rect 142620 677350 142860 677590
rect 142950 677350 143190 677590
rect 143300 677350 143540 677590
rect 143630 677350 143870 677590
rect 143960 677350 144200 677590
rect 144290 677350 144530 677590
rect 133570 677020 133810 677260
rect 133920 677020 134160 677260
rect 134250 677020 134490 677260
rect 134580 677020 134820 677260
rect 134910 677020 135150 677260
rect 135260 677020 135500 677260
rect 135590 677020 135830 677260
rect 135920 677020 136160 677260
rect 136250 677020 136490 677260
rect 136600 677020 136840 677260
rect 136930 677020 137170 677260
rect 137260 677020 137500 677260
rect 137590 677020 137830 677260
rect 137940 677020 138180 677260
rect 138270 677020 138510 677260
rect 138600 677020 138840 677260
rect 138930 677020 139170 677260
rect 139280 677020 139520 677260
rect 139610 677020 139850 677260
rect 139940 677020 140180 677260
rect 140270 677020 140510 677260
rect 140620 677020 140860 677260
rect 140950 677020 141190 677260
rect 141280 677020 141520 677260
rect 141610 677020 141850 677260
rect 141960 677020 142200 677260
rect 142290 677020 142530 677260
rect 142620 677020 142860 677260
rect 142950 677020 143190 677260
rect 143300 677020 143540 677260
rect 143630 677020 143870 677260
rect 143960 677020 144200 677260
rect 144290 677020 144530 677260
rect 133570 676690 133810 676930
rect 133920 676690 134160 676930
rect 134250 676690 134490 676930
rect 134580 676690 134820 676930
rect 134910 676690 135150 676930
rect 135260 676690 135500 676930
rect 135590 676690 135830 676930
rect 135920 676690 136160 676930
rect 136250 676690 136490 676930
rect 136600 676690 136840 676930
rect 136930 676690 137170 676930
rect 137260 676690 137500 676930
rect 137590 676690 137830 676930
rect 137940 676690 138180 676930
rect 138270 676690 138510 676930
rect 138600 676690 138840 676930
rect 138930 676690 139170 676930
rect 139280 676690 139520 676930
rect 139610 676690 139850 676930
rect 139940 676690 140180 676930
rect 140270 676690 140510 676930
rect 140620 676690 140860 676930
rect 140950 676690 141190 676930
rect 141280 676690 141520 676930
rect 141610 676690 141850 676930
rect 141960 676690 142200 676930
rect 142290 676690 142530 676930
rect 142620 676690 142860 676930
rect 142950 676690 143190 676930
rect 143300 676690 143540 676930
rect 143630 676690 143870 676930
rect 143960 676690 144200 676930
rect 144290 676690 144530 676930
rect 133570 676340 133810 676580
rect 133920 676340 134160 676580
rect 134250 676340 134490 676580
rect 134580 676340 134820 676580
rect 134910 676340 135150 676580
rect 135260 676340 135500 676580
rect 135590 676340 135830 676580
rect 135920 676340 136160 676580
rect 136250 676340 136490 676580
rect 136600 676340 136840 676580
rect 136930 676340 137170 676580
rect 137260 676340 137500 676580
rect 137590 676340 137830 676580
rect 137940 676340 138180 676580
rect 138270 676340 138510 676580
rect 138600 676340 138840 676580
rect 138930 676340 139170 676580
rect 139280 676340 139520 676580
rect 139610 676340 139850 676580
rect 139940 676340 140180 676580
rect 140270 676340 140510 676580
rect 140620 676340 140860 676580
rect 140950 676340 141190 676580
rect 141280 676340 141520 676580
rect 141610 676340 141850 676580
rect 141960 676340 142200 676580
rect 142290 676340 142530 676580
rect 142620 676340 142860 676580
rect 142950 676340 143190 676580
rect 143300 676340 143540 676580
rect 143630 676340 143870 676580
rect 143960 676340 144200 676580
rect 144290 676340 144530 676580
rect 133570 676010 133810 676250
rect 133920 676010 134160 676250
rect 134250 676010 134490 676250
rect 134580 676010 134820 676250
rect 134910 676010 135150 676250
rect 135260 676010 135500 676250
rect 135590 676010 135830 676250
rect 135920 676010 136160 676250
rect 136250 676010 136490 676250
rect 136600 676010 136840 676250
rect 136930 676010 137170 676250
rect 137260 676010 137500 676250
rect 137590 676010 137830 676250
rect 137940 676010 138180 676250
rect 138270 676010 138510 676250
rect 138600 676010 138840 676250
rect 138930 676010 139170 676250
rect 139280 676010 139520 676250
rect 139610 676010 139850 676250
rect 139940 676010 140180 676250
rect 140270 676010 140510 676250
rect 140620 676010 140860 676250
rect 140950 676010 141190 676250
rect 141280 676010 141520 676250
rect 141610 676010 141850 676250
rect 141960 676010 142200 676250
rect 142290 676010 142530 676250
rect 142620 676010 142860 676250
rect 142950 676010 143190 676250
rect 143300 676010 143540 676250
rect 143630 676010 143870 676250
rect 143960 676010 144200 676250
rect 144290 676010 144530 676250
rect 133570 675680 133810 675920
rect 133920 675680 134160 675920
rect 134250 675680 134490 675920
rect 134580 675680 134820 675920
rect 134910 675680 135150 675920
rect 135260 675680 135500 675920
rect 135590 675680 135830 675920
rect 135920 675680 136160 675920
rect 136250 675680 136490 675920
rect 136600 675680 136840 675920
rect 136930 675680 137170 675920
rect 137260 675680 137500 675920
rect 137590 675680 137830 675920
rect 137940 675680 138180 675920
rect 138270 675680 138510 675920
rect 138600 675680 138840 675920
rect 138930 675680 139170 675920
rect 139280 675680 139520 675920
rect 139610 675680 139850 675920
rect 139940 675680 140180 675920
rect 140270 675680 140510 675920
rect 140620 675680 140860 675920
rect 140950 675680 141190 675920
rect 141280 675680 141520 675920
rect 141610 675680 141850 675920
rect 141960 675680 142200 675920
rect 142290 675680 142530 675920
rect 142620 675680 142860 675920
rect 142950 675680 143190 675920
rect 143300 675680 143540 675920
rect 143630 675680 143870 675920
rect 143960 675680 144200 675920
rect 144290 675680 144530 675920
rect 133570 675350 133810 675590
rect 133920 675350 134160 675590
rect 134250 675350 134490 675590
rect 134580 675350 134820 675590
rect 134910 675350 135150 675590
rect 135260 675350 135500 675590
rect 135590 675350 135830 675590
rect 135920 675350 136160 675590
rect 136250 675350 136490 675590
rect 136600 675350 136840 675590
rect 136930 675350 137170 675590
rect 137260 675350 137500 675590
rect 137590 675350 137830 675590
rect 137940 675350 138180 675590
rect 138270 675350 138510 675590
rect 138600 675350 138840 675590
rect 138930 675350 139170 675590
rect 139280 675350 139520 675590
rect 139610 675350 139850 675590
rect 139940 675350 140180 675590
rect 140270 675350 140510 675590
rect 140620 675350 140860 675590
rect 140950 675350 141190 675590
rect 141280 675350 141520 675590
rect 141610 675350 141850 675590
rect 141960 675350 142200 675590
rect 142290 675350 142530 675590
rect 142620 675350 142860 675590
rect 142950 675350 143190 675590
rect 143300 675350 143540 675590
rect 143630 675350 143870 675590
rect 143960 675350 144200 675590
rect 144290 675350 144530 675590
rect 133570 675000 133810 675240
rect 133920 675000 134160 675240
rect 134250 675000 134490 675240
rect 134580 675000 134820 675240
rect 134910 675000 135150 675240
rect 135260 675000 135500 675240
rect 135590 675000 135830 675240
rect 135920 675000 136160 675240
rect 136250 675000 136490 675240
rect 136600 675000 136840 675240
rect 136930 675000 137170 675240
rect 137260 675000 137500 675240
rect 137590 675000 137830 675240
rect 137940 675000 138180 675240
rect 138270 675000 138510 675240
rect 138600 675000 138840 675240
rect 138930 675000 139170 675240
rect 139280 675000 139520 675240
rect 139610 675000 139850 675240
rect 139940 675000 140180 675240
rect 140270 675000 140510 675240
rect 140620 675000 140860 675240
rect 140950 675000 141190 675240
rect 141280 675000 141520 675240
rect 141610 675000 141850 675240
rect 141960 675000 142200 675240
rect 142290 675000 142530 675240
rect 142620 675000 142860 675240
rect 142950 675000 143190 675240
rect 143300 675000 143540 675240
rect 143630 675000 143870 675240
rect 143960 675000 144200 675240
rect 144290 675000 144530 675240
rect 133570 674670 133810 674910
rect 133920 674670 134160 674910
rect 134250 674670 134490 674910
rect 134580 674670 134820 674910
rect 134910 674670 135150 674910
rect 135260 674670 135500 674910
rect 135590 674670 135830 674910
rect 135920 674670 136160 674910
rect 136250 674670 136490 674910
rect 136600 674670 136840 674910
rect 136930 674670 137170 674910
rect 137260 674670 137500 674910
rect 137590 674670 137830 674910
rect 137940 674670 138180 674910
rect 138270 674670 138510 674910
rect 138600 674670 138840 674910
rect 138930 674670 139170 674910
rect 139280 674670 139520 674910
rect 139610 674670 139850 674910
rect 139940 674670 140180 674910
rect 140270 674670 140510 674910
rect 140620 674670 140860 674910
rect 140950 674670 141190 674910
rect 141280 674670 141520 674910
rect 141610 674670 141850 674910
rect 141960 674670 142200 674910
rect 142290 674670 142530 674910
rect 142620 674670 142860 674910
rect 142950 674670 143190 674910
rect 143300 674670 143540 674910
rect 143630 674670 143870 674910
rect 143960 674670 144200 674910
rect 144290 674670 144530 674910
rect 133570 674340 133810 674580
rect 133920 674340 134160 674580
rect 134250 674340 134490 674580
rect 134580 674340 134820 674580
rect 134910 674340 135150 674580
rect 135260 674340 135500 674580
rect 135590 674340 135830 674580
rect 135920 674340 136160 674580
rect 136250 674340 136490 674580
rect 136600 674340 136840 674580
rect 136930 674340 137170 674580
rect 137260 674340 137500 674580
rect 137590 674340 137830 674580
rect 137940 674340 138180 674580
rect 138270 674340 138510 674580
rect 138600 674340 138840 674580
rect 138930 674340 139170 674580
rect 139280 674340 139520 674580
rect 139610 674340 139850 674580
rect 139940 674340 140180 674580
rect 140270 674340 140510 674580
rect 140620 674340 140860 674580
rect 140950 674340 141190 674580
rect 141280 674340 141520 674580
rect 141610 674340 141850 674580
rect 141960 674340 142200 674580
rect 142290 674340 142530 674580
rect 142620 674340 142860 674580
rect 142950 674340 143190 674580
rect 143300 674340 143540 674580
rect 143630 674340 143870 674580
rect 143960 674340 144200 674580
rect 144290 674340 144530 674580
rect 133570 674010 133810 674250
rect 133920 674010 134160 674250
rect 134250 674010 134490 674250
rect 134580 674010 134820 674250
rect 134910 674010 135150 674250
rect 135260 674010 135500 674250
rect 135590 674010 135830 674250
rect 135920 674010 136160 674250
rect 136250 674010 136490 674250
rect 136600 674010 136840 674250
rect 136930 674010 137170 674250
rect 137260 674010 137500 674250
rect 137590 674010 137830 674250
rect 137940 674010 138180 674250
rect 138270 674010 138510 674250
rect 138600 674010 138840 674250
rect 138930 674010 139170 674250
rect 139280 674010 139520 674250
rect 139610 674010 139850 674250
rect 139940 674010 140180 674250
rect 140270 674010 140510 674250
rect 140620 674010 140860 674250
rect 140950 674010 141190 674250
rect 141280 674010 141520 674250
rect 141610 674010 141850 674250
rect 141960 674010 142200 674250
rect 142290 674010 142530 674250
rect 142620 674010 142860 674250
rect 142950 674010 143190 674250
rect 143300 674010 143540 674250
rect 143630 674010 143870 674250
rect 143960 674010 144200 674250
rect 144290 674010 144530 674250
rect 133570 673660 133810 673900
rect 133920 673660 134160 673900
rect 134250 673660 134490 673900
rect 134580 673660 134820 673900
rect 134910 673660 135150 673900
rect 135260 673660 135500 673900
rect 135590 673660 135830 673900
rect 135920 673660 136160 673900
rect 136250 673660 136490 673900
rect 136600 673660 136840 673900
rect 136930 673660 137170 673900
rect 137260 673660 137500 673900
rect 137590 673660 137830 673900
rect 137940 673660 138180 673900
rect 138270 673660 138510 673900
rect 138600 673660 138840 673900
rect 138930 673660 139170 673900
rect 139280 673660 139520 673900
rect 139610 673660 139850 673900
rect 139940 673660 140180 673900
rect 140270 673660 140510 673900
rect 140620 673660 140860 673900
rect 140950 673660 141190 673900
rect 141280 673660 141520 673900
rect 141610 673660 141850 673900
rect 141960 673660 142200 673900
rect 142290 673660 142530 673900
rect 142620 673660 142860 673900
rect 142950 673660 143190 673900
rect 143300 673660 143540 673900
rect 143630 673660 143870 673900
rect 143960 673660 144200 673900
rect 144290 673660 144530 673900
rect 133570 673330 133810 673570
rect 133920 673330 134160 673570
rect 134250 673330 134490 673570
rect 134580 673330 134820 673570
rect 134910 673330 135150 673570
rect 135260 673330 135500 673570
rect 135590 673330 135830 673570
rect 135920 673330 136160 673570
rect 136250 673330 136490 673570
rect 136600 673330 136840 673570
rect 136930 673330 137170 673570
rect 137260 673330 137500 673570
rect 137590 673330 137830 673570
rect 137940 673330 138180 673570
rect 138270 673330 138510 673570
rect 138600 673330 138840 673570
rect 138930 673330 139170 673570
rect 139280 673330 139520 673570
rect 139610 673330 139850 673570
rect 139940 673330 140180 673570
rect 140270 673330 140510 673570
rect 140620 673330 140860 673570
rect 140950 673330 141190 673570
rect 141280 673330 141520 673570
rect 141610 673330 141850 673570
rect 141960 673330 142200 673570
rect 142290 673330 142530 673570
rect 142620 673330 142860 673570
rect 142950 673330 143190 673570
rect 143300 673330 143540 673570
rect 143630 673330 143870 673570
rect 143960 673330 144200 673570
rect 144290 673330 144530 673570
rect 133570 673000 133810 673240
rect 133920 673000 134160 673240
rect 134250 673000 134490 673240
rect 134580 673000 134820 673240
rect 134910 673000 135150 673240
rect 135260 673000 135500 673240
rect 135590 673000 135830 673240
rect 135920 673000 136160 673240
rect 136250 673000 136490 673240
rect 136600 673000 136840 673240
rect 136930 673000 137170 673240
rect 137260 673000 137500 673240
rect 137590 673000 137830 673240
rect 137940 673000 138180 673240
rect 138270 673000 138510 673240
rect 138600 673000 138840 673240
rect 138930 673000 139170 673240
rect 139280 673000 139520 673240
rect 139610 673000 139850 673240
rect 139940 673000 140180 673240
rect 140270 673000 140510 673240
rect 140620 673000 140860 673240
rect 140950 673000 141190 673240
rect 141280 673000 141520 673240
rect 141610 673000 141850 673240
rect 141960 673000 142200 673240
rect 142290 673000 142530 673240
rect 142620 673000 142860 673240
rect 142950 673000 143190 673240
rect 143300 673000 143540 673240
rect 143630 673000 143870 673240
rect 143960 673000 144200 673240
rect 144290 673000 144530 673240
rect 133570 672670 133810 672910
rect 133920 672670 134160 672910
rect 134250 672670 134490 672910
rect 134580 672670 134820 672910
rect 134910 672670 135150 672910
rect 135260 672670 135500 672910
rect 135590 672670 135830 672910
rect 135920 672670 136160 672910
rect 136250 672670 136490 672910
rect 136600 672670 136840 672910
rect 136930 672670 137170 672910
rect 137260 672670 137500 672910
rect 137590 672670 137830 672910
rect 137940 672670 138180 672910
rect 138270 672670 138510 672910
rect 138600 672670 138840 672910
rect 138930 672670 139170 672910
rect 139280 672670 139520 672910
rect 139610 672670 139850 672910
rect 139940 672670 140180 672910
rect 140270 672670 140510 672910
rect 140620 672670 140860 672910
rect 140950 672670 141190 672910
rect 141280 672670 141520 672910
rect 141610 672670 141850 672910
rect 141960 672670 142200 672910
rect 142290 672670 142530 672910
rect 142620 672670 142860 672910
rect 142950 672670 143190 672910
rect 143300 672670 143540 672910
rect 143630 672670 143870 672910
rect 143960 672670 144200 672910
rect 144290 672670 144530 672910
rect 133570 672320 133810 672560
rect 133920 672320 134160 672560
rect 134250 672320 134490 672560
rect 134580 672320 134820 672560
rect 134910 672320 135150 672560
rect 135260 672320 135500 672560
rect 135590 672320 135830 672560
rect 135920 672320 136160 672560
rect 136250 672320 136490 672560
rect 136600 672320 136840 672560
rect 136930 672320 137170 672560
rect 137260 672320 137500 672560
rect 137590 672320 137830 672560
rect 137940 672320 138180 672560
rect 138270 672320 138510 672560
rect 138600 672320 138840 672560
rect 138930 672320 139170 672560
rect 139280 672320 139520 672560
rect 139610 672320 139850 672560
rect 139940 672320 140180 672560
rect 140270 672320 140510 672560
rect 140620 672320 140860 672560
rect 140950 672320 141190 672560
rect 141280 672320 141520 672560
rect 141610 672320 141850 672560
rect 141960 672320 142200 672560
rect 142290 672320 142530 672560
rect 142620 672320 142860 672560
rect 142950 672320 143190 672560
rect 143300 672320 143540 672560
rect 143630 672320 143870 672560
rect 143960 672320 144200 672560
rect 144290 672320 144530 672560
rect 144950 683040 145190 683280
rect 145300 683040 145540 683280
rect 145630 683040 145870 683280
rect 145960 683040 146200 683280
rect 146290 683040 146530 683280
rect 146640 683040 146880 683280
rect 146970 683040 147210 683280
rect 147300 683040 147540 683280
rect 147630 683040 147870 683280
rect 147980 683040 148220 683280
rect 148310 683040 148550 683280
rect 148640 683040 148880 683280
rect 148970 683040 149210 683280
rect 149320 683040 149560 683280
rect 149650 683040 149890 683280
rect 149980 683040 150220 683280
rect 150310 683040 150550 683280
rect 150660 683040 150900 683280
rect 150990 683040 151230 683280
rect 151320 683040 151560 683280
rect 151650 683040 151890 683280
rect 152000 683040 152240 683280
rect 152330 683040 152570 683280
rect 152660 683040 152900 683280
rect 152990 683040 153230 683280
rect 153340 683040 153580 683280
rect 153670 683040 153910 683280
rect 154000 683040 154240 683280
rect 154330 683040 154570 683280
rect 154680 683040 154920 683280
rect 155010 683040 155250 683280
rect 155340 683040 155580 683280
rect 155670 683040 155910 683280
rect 144950 682710 145190 682950
rect 145300 682710 145540 682950
rect 145630 682710 145870 682950
rect 145960 682710 146200 682950
rect 146290 682710 146530 682950
rect 146640 682710 146880 682950
rect 146970 682710 147210 682950
rect 147300 682710 147540 682950
rect 147630 682710 147870 682950
rect 147980 682710 148220 682950
rect 148310 682710 148550 682950
rect 148640 682710 148880 682950
rect 148970 682710 149210 682950
rect 149320 682710 149560 682950
rect 149650 682710 149890 682950
rect 149980 682710 150220 682950
rect 150310 682710 150550 682950
rect 150660 682710 150900 682950
rect 150990 682710 151230 682950
rect 151320 682710 151560 682950
rect 151650 682710 151890 682950
rect 152000 682710 152240 682950
rect 152330 682710 152570 682950
rect 152660 682710 152900 682950
rect 152990 682710 153230 682950
rect 153340 682710 153580 682950
rect 153670 682710 153910 682950
rect 154000 682710 154240 682950
rect 154330 682710 154570 682950
rect 154680 682710 154920 682950
rect 155010 682710 155250 682950
rect 155340 682710 155580 682950
rect 155670 682710 155910 682950
rect 144950 682380 145190 682620
rect 145300 682380 145540 682620
rect 145630 682380 145870 682620
rect 145960 682380 146200 682620
rect 146290 682380 146530 682620
rect 146640 682380 146880 682620
rect 146970 682380 147210 682620
rect 147300 682380 147540 682620
rect 147630 682380 147870 682620
rect 147980 682380 148220 682620
rect 148310 682380 148550 682620
rect 148640 682380 148880 682620
rect 148970 682380 149210 682620
rect 149320 682380 149560 682620
rect 149650 682380 149890 682620
rect 149980 682380 150220 682620
rect 150310 682380 150550 682620
rect 150660 682380 150900 682620
rect 150990 682380 151230 682620
rect 151320 682380 151560 682620
rect 151650 682380 151890 682620
rect 152000 682380 152240 682620
rect 152330 682380 152570 682620
rect 152660 682380 152900 682620
rect 152990 682380 153230 682620
rect 153340 682380 153580 682620
rect 153670 682380 153910 682620
rect 154000 682380 154240 682620
rect 154330 682380 154570 682620
rect 154680 682380 154920 682620
rect 155010 682380 155250 682620
rect 155340 682380 155580 682620
rect 155670 682380 155910 682620
rect 144950 682050 145190 682290
rect 145300 682050 145540 682290
rect 145630 682050 145870 682290
rect 145960 682050 146200 682290
rect 146290 682050 146530 682290
rect 146640 682050 146880 682290
rect 146970 682050 147210 682290
rect 147300 682050 147540 682290
rect 147630 682050 147870 682290
rect 147980 682050 148220 682290
rect 148310 682050 148550 682290
rect 148640 682050 148880 682290
rect 148970 682050 149210 682290
rect 149320 682050 149560 682290
rect 149650 682050 149890 682290
rect 149980 682050 150220 682290
rect 150310 682050 150550 682290
rect 150660 682050 150900 682290
rect 150990 682050 151230 682290
rect 151320 682050 151560 682290
rect 151650 682050 151890 682290
rect 152000 682050 152240 682290
rect 152330 682050 152570 682290
rect 152660 682050 152900 682290
rect 152990 682050 153230 682290
rect 153340 682050 153580 682290
rect 153670 682050 153910 682290
rect 154000 682050 154240 682290
rect 154330 682050 154570 682290
rect 154680 682050 154920 682290
rect 155010 682050 155250 682290
rect 155340 682050 155580 682290
rect 155670 682050 155910 682290
rect 144950 681700 145190 681940
rect 145300 681700 145540 681940
rect 145630 681700 145870 681940
rect 145960 681700 146200 681940
rect 146290 681700 146530 681940
rect 146640 681700 146880 681940
rect 146970 681700 147210 681940
rect 147300 681700 147540 681940
rect 147630 681700 147870 681940
rect 147980 681700 148220 681940
rect 148310 681700 148550 681940
rect 148640 681700 148880 681940
rect 148970 681700 149210 681940
rect 149320 681700 149560 681940
rect 149650 681700 149890 681940
rect 149980 681700 150220 681940
rect 150310 681700 150550 681940
rect 150660 681700 150900 681940
rect 150990 681700 151230 681940
rect 151320 681700 151560 681940
rect 151650 681700 151890 681940
rect 152000 681700 152240 681940
rect 152330 681700 152570 681940
rect 152660 681700 152900 681940
rect 152990 681700 153230 681940
rect 153340 681700 153580 681940
rect 153670 681700 153910 681940
rect 154000 681700 154240 681940
rect 154330 681700 154570 681940
rect 154680 681700 154920 681940
rect 155010 681700 155250 681940
rect 155340 681700 155580 681940
rect 155670 681700 155910 681940
rect 144950 681370 145190 681610
rect 145300 681370 145540 681610
rect 145630 681370 145870 681610
rect 145960 681370 146200 681610
rect 146290 681370 146530 681610
rect 146640 681370 146880 681610
rect 146970 681370 147210 681610
rect 147300 681370 147540 681610
rect 147630 681370 147870 681610
rect 147980 681370 148220 681610
rect 148310 681370 148550 681610
rect 148640 681370 148880 681610
rect 148970 681370 149210 681610
rect 149320 681370 149560 681610
rect 149650 681370 149890 681610
rect 149980 681370 150220 681610
rect 150310 681370 150550 681610
rect 150660 681370 150900 681610
rect 150990 681370 151230 681610
rect 151320 681370 151560 681610
rect 151650 681370 151890 681610
rect 152000 681370 152240 681610
rect 152330 681370 152570 681610
rect 152660 681370 152900 681610
rect 152990 681370 153230 681610
rect 153340 681370 153580 681610
rect 153670 681370 153910 681610
rect 154000 681370 154240 681610
rect 154330 681370 154570 681610
rect 154680 681370 154920 681610
rect 155010 681370 155250 681610
rect 155340 681370 155580 681610
rect 155670 681370 155910 681610
rect 144950 681040 145190 681280
rect 145300 681040 145540 681280
rect 145630 681040 145870 681280
rect 145960 681040 146200 681280
rect 146290 681040 146530 681280
rect 146640 681040 146880 681280
rect 146970 681040 147210 681280
rect 147300 681040 147540 681280
rect 147630 681040 147870 681280
rect 147980 681040 148220 681280
rect 148310 681040 148550 681280
rect 148640 681040 148880 681280
rect 148970 681040 149210 681280
rect 149320 681040 149560 681280
rect 149650 681040 149890 681280
rect 149980 681040 150220 681280
rect 150310 681040 150550 681280
rect 150660 681040 150900 681280
rect 150990 681040 151230 681280
rect 151320 681040 151560 681280
rect 151650 681040 151890 681280
rect 152000 681040 152240 681280
rect 152330 681040 152570 681280
rect 152660 681040 152900 681280
rect 152990 681040 153230 681280
rect 153340 681040 153580 681280
rect 153670 681040 153910 681280
rect 154000 681040 154240 681280
rect 154330 681040 154570 681280
rect 154680 681040 154920 681280
rect 155010 681040 155250 681280
rect 155340 681040 155580 681280
rect 155670 681040 155910 681280
rect 144950 680710 145190 680950
rect 145300 680710 145540 680950
rect 145630 680710 145870 680950
rect 145960 680710 146200 680950
rect 146290 680710 146530 680950
rect 146640 680710 146880 680950
rect 146970 680710 147210 680950
rect 147300 680710 147540 680950
rect 147630 680710 147870 680950
rect 147980 680710 148220 680950
rect 148310 680710 148550 680950
rect 148640 680710 148880 680950
rect 148970 680710 149210 680950
rect 149320 680710 149560 680950
rect 149650 680710 149890 680950
rect 149980 680710 150220 680950
rect 150310 680710 150550 680950
rect 150660 680710 150900 680950
rect 150990 680710 151230 680950
rect 151320 680710 151560 680950
rect 151650 680710 151890 680950
rect 152000 680710 152240 680950
rect 152330 680710 152570 680950
rect 152660 680710 152900 680950
rect 152990 680710 153230 680950
rect 153340 680710 153580 680950
rect 153670 680710 153910 680950
rect 154000 680710 154240 680950
rect 154330 680710 154570 680950
rect 154680 680710 154920 680950
rect 155010 680710 155250 680950
rect 155340 680710 155580 680950
rect 155670 680710 155910 680950
rect 144950 680360 145190 680600
rect 145300 680360 145540 680600
rect 145630 680360 145870 680600
rect 145960 680360 146200 680600
rect 146290 680360 146530 680600
rect 146640 680360 146880 680600
rect 146970 680360 147210 680600
rect 147300 680360 147540 680600
rect 147630 680360 147870 680600
rect 147980 680360 148220 680600
rect 148310 680360 148550 680600
rect 148640 680360 148880 680600
rect 148970 680360 149210 680600
rect 149320 680360 149560 680600
rect 149650 680360 149890 680600
rect 149980 680360 150220 680600
rect 150310 680360 150550 680600
rect 150660 680360 150900 680600
rect 150990 680360 151230 680600
rect 151320 680360 151560 680600
rect 151650 680360 151890 680600
rect 152000 680360 152240 680600
rect 152330 680360 152570 680600
rect 152660 680360 152900 680600
rect 152990 680360 153230 680600
rect 153340 680360 153580 680600
rect 153670 680360 153910 680600
rect 154000 680360 154240 680600
rect 154330 680360 154570 680600
rect 154680 680360 154920 680600
rect 155010 680360 155250 680600
rect 155340 680360 155580 680600
rect 155670 680360 155910 680600
rect 144950 680030 145190 680270
rect 145300 680030 145540 680270
rect 145630 680030 145870 680270
rect 145960 680030 146200 680270
rect 146290 680030 146530 680270
rect 146640 680030 146880 680270
rect 146970 680030 147210 680270
rect 147300 680030 147540 680270
rect 147630 680030 147870 680270
rect 147980 680030 148220 680270
rect 148310 680030 148550 680270
rect 148640 680030 148880 680270
rect 148970 680030 149210 680270
rect 149320 680030 149560 680270
rect 149650 680030 149890 680270
rect 149980 680030 150220 680270
rect 150310 680030 150550 680270
rect 150660 680030 150900 680270
rect 150990 680030 151230 680270
rect 151320 680030 151560 680270
rect 151650 680030 151890 680270
rect 152000 680030 152240 680270
rect 152330 680030 152570 680270
rect 152660 680030 152900 680270
rect 152990 680030 153230 680270
rect 153340 680030 153580 680270
rect 153670 680030 153910 680270
rect 154000 680030 154240 680270
rect 154330 680030 154570 680270
rect 154680 680030 154920 680270
rect 155010 680030 155250 680270
rect 155340 680030 155580 680270
rect 155670 680030 155910 680270
rect 144950 679700 145190 679940
rect 145300 679700 145540 679940
rect 145630 679700 145870 679940
rect 145960 679700 146200 679940
rect 146290 679700 146530 679940
rect 146640 679700 146880 679940
rect 146970 679700 147210 679940
rect 147300 679700 147540 679940
rect 147630 679700 147870 679940
rect 147980 679700 148220 679940
rect 148310 679700 148550 679940
rect 148640 679700 148880 679940
rect 148970 679700 149210 679940
rect 149320 679700 149560 679940
rect 149650 679700 149890 679940
rect 149980 679700 150220 679940
rect 150310 679700 150550 679940
rect 150660 679700 150900 679940
rect 150990 679700 151230 679940
rect 151320 679700 151560 679940
rect 151650 679700 151890 679940
rect 152000 679700 152240 679940
rect 152330 679700 152570 679940
rect 152660 679700 152900 679940
rect 152990 679700 153230 679940
rect 153340 679700 153580 679940
rect 153670 679700 153910 679940
rect 154000 679700 154240 679940
rect 154330 679700 154570 679940
rect 154680 679700 154920 679940
rect 155010 679700 155250 679940
rect 155340 679700 155580 679940
rect 155670 679700 155910 679940
rect 144950 679370 145190 679610
rect 145300 679370 145540 679610
rect 145630 679370 145870 679610
rect 145960 679370 146200 679610
rect 146290 679370 146530 679610
rect 146640 679370 146880 679610
rect 146970 679370 147210 679610
rect 147300 679370 147540 679610
rect 147630 679370 147870 679610
rect 147980 679370 148220 679610
rect 148310 679370 148550 679610
rect 148640 679370 148880 679610
rect 148970 679370 149210 679610
rect 149320 679370 149560 679610
rect 149650 679370 149890 679610
rect 149980 679370 150220 679610
rect 150310 679370 150550 679610
rect 150660 679370 150900 679610
rect 150990 679370 151230 679610
rect 151320 679370 151560 679610
rect 151650 679370 151890 679610
rect 152000 679370 152240 679610
rect 152330 679370 152570 679610
rect 152660 679370 152900 679610
rect 152990 679370 153230 679610
rect 153340 679370 153580 679610
rect 153670 679370 153910 679610
rect 154000 679370 154240 679610
rect 154330 679370 154570 679610
rect 154680 679370 154920 679610
rect 155010 679370 155250 679610
rect 155340 679370 155580 679610
rect 155670 679370 155910 679610
rect 144950 679020 145190 679260
rect 145300 679020 145540 679260
rect 145630 679020 145870 679260
rect 145960 679020 146200 679260
rect 146290 679020 146530 679260
rect 146640 679020 146880 679260
rect 146970 679020 147210 679260
rect 147300 679020 147540 679260
rect 147630 679020 147870 679260
rect 147980 679020 148220 679260
rect 148310 679020 148550 679260
rect 148640 679020 148880 679260
rect 148970 679020 149210 679260
rect 149320 679020 149560 679260
rect 149650 679020 149890 679260
rect 149980 679020 150220 679260
rect 150310 679020 150550 679260
rect 150660 679020 150900 679260
rect 150990 679020 151230 679260
rect 151320 679020 151560 679260
rect 151650 679020 151890 679260
rect 152000 679020 152240 679260
rect 152330 679020 152570 679260
rect 152660 679020 152900 679260
rect 152990 679020 153230 679260
rect 153340 679020 153580 679260
rect 153670 679020 153910 679260
rect 154000 679020 154240 679260
rect 154330 679020 154570 679260
rect 154680 679020 154920 679260
rect 155010 679020 155250 679260
rect 155340 679020 155580 679260
rect 155670 679020 155910 679260
rect 144950 678690 145190 678930
rect 145300 678690 145540 678930
rect 145630 678690 145870 678930
rect 145960 678690 146200 678930
rect 146290 678690 146530 678930
rect 146640 678690 146880 678930
rect 146970 678690 147210 678930
rect 147300 678690 147540 678930
rect 147630 678690 147870 678930
rect 147980 678690 148220 678930
rect 148310 678690 148550 678930
rect 148640 678690 148880 678930
rect 148970 678690 149210 678930
rect 149320 678690 149560 678930
rect 149650 678690 149890 678930
rect 149980 678690 150220 678930
rect 150310 678690 150550 678930
rect 150660 678690 150900 678930
rect 150990 678690 151230 678930
rect 151320 678690 151560 678930
rect 151650 678690 151890 678930
rect 152000 678690 152240 678930
rect 152330 678690 152570 678930
rect 152660 678690 152900 678930
rect 152990 678690 153230 678930
rect 153340 678690 153580 678930
rect 153670 678690 153910 678930
rect 154000 678690 154240 678930
rect 154330 678690 154570 678930
rect 154680 678690 154920 678930
rect 155010 678690 155250 678930
rect 155340 678690 155580 678930
rect 155670 678690 155910 678930
rect 144950 678360 145190 678600
rect 145300 678360 145540 678600
rect 145630 678360 145870 678600
rect 145960 678360 146200 678600
rect 146290 678360 146530 678600
rect 146640 678360 146880 678600
rect 146970 678360 147210 678600
rect 147300 678360 147540 678600
rect 147630 678360 147870 678600
rect 147980 678360 148220 678600
rect 148310 678360 148550 678600
rect 148640 678360 148880 678600
rect 148970 678360 149210 678600
rect 149320 678360 149560 678600
rect 149650 678360 149890 678600
rect 149980 678360 150220 678600
rect 150310 678360 150550 678600
rect 150660 678360 150900 678600
rect 150990 678360 151230 678600
rect 151320 678360 151560 678600
rect 151650 678360 151890 678600
rect 152000 678360 152240 678600
rect 152330 678360 152570 678600
rect 152660 678360 152900 678600
rect 152990 678360 153230 678600
rect 153340 678360 153580 678600
rect 153670 678360 153910 678600
rect 154000 678360 154240 678600
rect 154330 678360 154570 678600
rect 154680 678360 154920 678600
rect 155010 678360 155250 678600
rect 155340 678360 155580 678600
rect 155670 678360 155910 678600
rect 144950 678030 145190 678270
rect 145300 678030 145540 678270
rect 145630 678030 145870 678270
rect 145960 678030 146200 678270
rect 146290 678030 146530 678270
rect 146640 678030 146880 678270
rect 146970 678030 147210 678270
rect 147300 678030 147540 678270
rect 147630 678030 147870 678270
rect 147980 678030 148220 678270
rect 148310 678030 148550 678270
rect 148640 678030 148880 678270
rect 148970 678030 149210 678270
rect 149320 678030 149560 678270
rect 149650 678030 149890 678270
rect 149980 678030 150220 678270
rect 150310 678030 150550 678270
rect 150660 678030 150900 678270
rect 150990 678030 151230 678270
rect 151320 678030 151560 678270
rect 151650 678030 151890 678270
rect 152000 678030 152240 678270
rect 152330 678030 152570 678270
rect 152660 678030 152900 678270
rect 152990 678030 153230 678270
rect 153340 678030 153580 678270
rect 153670 678030 153910 678270
rect 154000 678030 154240 678270
rect 154330 678030 154570 678270
rect 154680 678030 154920 678270
rect 155010 678030 155250 678270
rect 155340 678030 155580 678270
rect 155670 678030 155910 678270
rect 144950 677680 145190 677920
rect 145300 677680 145540 677920
rect 145630 677680 145870 677920
rect 145960 677680 146200 677920
rect 146290 677680 146530 677920
rect 146640 677680 146880 677920
rect 146970 677680 147210 677920
rect 147300 677680 147540 677920
rect 147630 677680 147870 677920
rect 147980 677680 148220 677920
rect 148310 677680 148550 677920
rect 148640 677680 148880 677920
rect 148970 677680 149210 677920
rect 149320 677680 149560 677920
rect 149650 677680 149890 677920
rect 149980 677680 150220 677920
rect 150310 677680 150550 677920
rect 150660 677680 150900 677920
rect 150990 677680 151230 677920
rect 151320 677680 151560 677920
rect 151650 677680 151890 677920
rect 152000 677680 152240 677920
rect 152330 677680 152570 677920
rect 152660 677680 152900 677920
rect 152990 677680 153230 677920
rect 153340 677680 153580 677920
rect 153670 677680 153910 677920
rect 154000 677680 154240 677920
rect 154330 677680 154570 677920
rect 154680 677680 154920 677920
rect 155010 677680 155250 677920
rect 155340 677680 155580 677920
rect 155670 677680 155910 677920
rect 144950 677350 145190 677590
rect 145300 677350 145540 677590
rect 145630 677350 145870 677590
rect 145960 677350 146200 677590
rect 146290 677350 146530 677590
rect 146640 677350 146880 677590
rect 146970 677350 147210 677590
rect 147300 677350 147540 677590
rect 147630 677350 147870 677590
rect 147980 677350 148220 677590
rect 148310 677350 148550 677590
rect 148640 677350 148880 677590
rect 148970 677350 149210 677590
rect 149320 677350 149560 677590
rect 149650 677350 149890 677590
rect 149980 677350 150220 677590
rect 150310 677350 150550 677590
rect 150660 677350 150900 677590
rect 150990 677350 151230 677590
rect 151320 677350 151560 677590
rect 151650 677350 151890 677590
rect 152000 677350 152240 677590
rect 152330 677350 152570 677590
rect 152660 677350 152900 677590
rect 152990 677350 153230 677590
rect 153340 677350 153580 677590
rect 153670 677350 153910 677590
rect 154000 677350 154240 677590
rect 154330 677350 154570 677590
rect 154680 677350 154920 677590
rect 155010 677350 155250 677590
rect 155340 677350 155580 677590
rect 155670 677350 155910 677590
rect 144950 677020 145190 677260
rect 145300 677020 145540 677260
rect 145630 677020 145870 677260
rect 145960 677020 146200 677260
rect 146290 677020 146530 677260
rect 146640 677020 146880 677260
rect 146970 677020 147210 677260
rect 147300 677020 147540 677260
rect 147630 677020 147870 677260
rect 147980 677020 148220 677260
rect 148310 677020 148550 677260
rect 148640 677020 148880 677260
rect 148970 677020 149210 677260
rect 149320 677020 149560 677260
rect 149650 677020 149890 677260
rect 149980 677020 150220 677260
rect 150310 677020 150550 677260
rect 150660 677020 150900 677260
rect 150990 677020 151230 677260
rect 151320 677020 151560 677260
rect 151650 677020 151890 677260
rect 152000 677020 152240 677260
rect 152330 677020 152570 677260
rect 152660 677020 152900 677260
rect 152990 677020 153230 677260
rect 153340 677020 153580 677260
rect 153670 677020 153910 677260
rect 154000 677020 154240 677260
rect 154330 677020 154570 677260
rect 154680 677020 154920 677260
rect 155010 677020 155250 677260
rect 155340 677020 155580 677260
rect 155670 677020 155910 677260
rect 144950 676690 145190 676930
rect 145300 676690 145540 676930
rect 145630 676690 145870 676930
rect 145960 676690 146200 676930
rect 146290 676690 146530 676930
rect 146640 676690 146880 676930
rect 146970 676690 147210 676930
rect 147300 676690 147540 676930
rect 147630 676690 147870 676930
rect 147980 676690 148220 676930
rect 148310 676690 148550 676930
rect 148640 676690 148880 676930
rect 148970 676690 149210 676930
rect 149320 676690 149560 676930
rect 149650 676690 149890 676930
rect 149980 676690 150220 676930
rect 150310 676690 150550 676930
rect 150660 676690 150900 676930
rect 150990 676690 151230 676930
rect 151320 676690 151560 676930
rect 151650 676690 151890 676930
rect 152000 676690 152240 676930
rect 152330 676690 152570 676930
rect 152660 676690 152900 676930
rect 152990 676690 153230 676930
rect 153340 676690 153580 676930
rect 153670 676690 153910 676930
rect 154000 676690 154240 676930
rect 154330 676690 154570 676930
rect 154680 676690 154920 676930
rect 155010 676690 155250 676930
rect 155340 676690 155580 676930
rect 155670 676690 155910 676930
rect 144950 676340 145190 676580
rect 145300 676340 145540 676580
rect 145630 676340 145870 676580
rect 145960 676340 146200 676580
rect 146290 676340 146530 676580
rect 146640 676340 146880 676580
rect 146970 676340 147210 676580
rect 147300 676340 147540 676580
rect 147630 676340 147870 676580
rect 147980 676340 148220 676580
rect 148310 676340 148550 676580
rect 148640 676340 148880 676580
rect 148970 676340 149210 676580
rect 149320 676340 149560 676580
rect 149650 676340 149890 676580
rect 149980 676340 150220 676580
rect 150310 676340 150550 676580
rect 150660 676340 150900 676580
rect 150990 676340 151230 676580
rect 151320 676340 151560 676580
rect 151650 676340 151890 676580
rect 152000 676340 152240 676580
rect 152330 676340 152570 676580
rect 152660 676340 152900 676580
rect 152990 676340 153230 676580
rect 153340 676340 153580 676580
rect 153670 676340 153910 676580
rect 154000 676340 154240 676580
rect 154330 676340 154570 676580
rect 154680 676340 154920 676580
rect 155010 676340 155250 676580
rect 155340 676340 155580 676580
rect 155670 676340 155910 676580
rect 144950 676010 145190 676250
rect 145300 676010 145540 676250
rect 145630 676010 145870 676250
rect 145960 676010 146200 676250
rect 146290 676010 146530 676250
rect 146640 676010 146880 676250
rect 146970 676010 147210 676250
rect 147300 676010 147540 676250
rect 147630 676010 147870 676250
rect 147980 676010 148220 676250
rect 148310 676010 148550 676250
rect 148640 676010 148880 676250
rect 148970 676010 149210 676250
rect 149320 676010 149560 676250
rect 149650 676010 149890 676250
rect 149980 676010 150220 676250
rect 150310 676010 150550 676250
rect 150660 676010 150900 676250
rect 150990 676010 151230 676250
rect 151320 676010 151560 676250
rect 151650 676010 151890 676250
rect 152000 676010 152240 676250
rect 152330 676010 152570 676250
rect 152660 676010 152900 676250
rect 152990 676010 153230 676250
rect 153340 676010 153580 676250
rect 153670 676010 153910 676250
rect 154000 676010 154240 676250
rect 154330 676010 154570 676250
rect 154680 676010 154920 676250
rect 155010 676010 155250 676250
rect 155340 676010 155580 676250
rect 155670 676010 155910 676250
rect 144950 675680 145190 675920
rect 145300 675680 145540 675920
rect 145630 675680 145870 675920
rect 145960 675680 146200 675920
rect 146290 675680 146530 675920
rect 146640 675680 146880 675920
rect 146970 675680 147210 675920
rect 147300 675680 147540 675920
rect 147630 675680 147870 675920
rect 147980 675680 148220 675920
rect 148310 675680 148550 675920
rect 148640 675680 148880 675920
rect 148970 675680 149210 675920
rect 149320 675680 149560 675920
rect 149650 675680 149890 675920
rect 149980 675680 150220 675920
rect 150310 675680 150550 675920
rect 150660 675680 150900 675920
rect 150990 675680 151230 675920
rect 151320 675680 151560 675920
rect 151650 675680 151890 675920
rect 152000 675680 152240 675920
rect 152330 675680 152570 675920
rect 152660 675680 152900 675920
rect 152990 675680 153230 675920
rect 153340 675680 153580 675920
rect 153670 675680 153910 675920
rect 154000 675680 154240 675920
rect 154330 675680 154570 675920
rect 154680 675680 154920 675920
rect 155010 675680 155250 675920
rect 155340 675680 155580 675920
rect 155670 675680 155910 675920
rect 144950 675350 145190 675590
rect 145300 675350 145540 675590
rect 145630 675350 145870 675590
rect 145960 675350 146200 675590
rect 146290 675350 146530 675590
rect 146640 675350 146880 675590
rect 146970 675350 147210 675590
rect 147300 675350 147540 675590
rect 147630 675350 147870 675590
rect 147980 675350 148220 675590
rect 148310 675350 148550 675590
rect 148640 675350 148880 675590
rect 148970 675350 149210 675590
rect 149320 675350 149560 675590
rect 149650 675350 149890 675590
rect 149980 675350 150220 675590
rect 150310 675350 150550 675590
rect 150660 675350 150900 675590
rect 150990 675350 151230 675590
rect 151320 675350 151560 675590
rect 151650 675350 151890 675590
rect 152000 675350 152240 675590
rect 152330 675350 152570 675590
rect 152660 675350 152900 675590
rect 152990 675350 153230 675590
rect 153340 675350 153580 675590
rect 153670 675350 153910 675590
rect 154000 675350 154240 675590
rect 154330 675350 154570 675590
rect 154680 675350 154920 675590
rect 155010 675350 155250 675590
rect 155340 675350 155580 675590
rect 155670 675350 155910 675590
rect 144950 675000 145190 675240
rect 145300 675000 145540 675240
rect 145630 675000 145870 675240
rect 145960 675000 146200 675240
rect 146290 675000 146530 675240
rect 146640 675000 146880 675240
rect 146970 675000 147210 675240
rect 147300 675000 147540 675240
rect 147630 675000 147870 675240
rect 147980 675000 148220 675240
rect 148310 675000 148550 675240
rect 148640 675000 148880 675240
rect 148970 675000 149210 675240
rect 149320 675000 149560 675240
rect 149650 675000 149890 675240
rect 149980 675000 150220 675240
rect 150310 675000 150550 675240
rect 150660 675000 150900 675240
rect 150990 675000 151230 675240
rect 151320 675000 151560 675240
rect 151650 675000 151890 675240
rect 152000 675000 152240 675240
rect 152330 675000 152570 675240
rect 152660 675000 152900 675240
rect 152990 675000 153230 675240
rect 153340 675000 153580 675240
rect 153670 675000 153910 675240
rect 154000 675000 154240 675240
rect 154330 675000 154570 675240
rect 154680 675000 154920 675240
rect 155010 675000 155250 675240
rect 155340 675000 155580 675240
rect 155670 675000 155910 675240
rect 144950 674670 145190 674910
rect 145300 674670 145540 674910
rect 145630 674670 145870 674910
rect 145960 674670 146200 674910
rect 146290 674670 146530 674910
rect 146640 674670 146880 674910
rect 146970 674670 147210 674910
rect 147300 674670 147540 674910
rect 147630 674670 147870 674910
rect 147980 674670 148220 674910
rect 148310 674670 148550 674910
rect 148640 674670 148880 674910
rect 148970 674670 149210 674910
rect 149320 674670 149560 674910
rect 149650 674670 149890 674910
rect 149980 674670 150220 674910
rect 150310 674670 150550 674910
rect 150660 674670 150900 674910
rect 150990 674670 151230 674910
rect 151320 674670 151560 674910
rect 151650 674670 151890 674910
rect 152000 674670 152240 674910
rect 152330 674670 152570 674910
rect 152660 674670 152900 674910
rect 152990 674670 153230 674910
rect 153340 674670 153580 674910
rect 153670 674670 153910 674910
rect 154000 674670 154240 674910
rect 154330 674670 154570 674910
rect 154680 674670 154920 674910
rect 155010 674670 155250 674910
rect 155340 674670 155580 674910
rect 155670 674670 155910 674910
rect 144950 674340 145190 674580
rect 145300 674340 145540 674580
rect 145630 674340 145870 674580
rect 145960 674340 146200 674580
rect 146290 674340 146530 674580
rect 146640 674340 146880 674580
rect 146970 674340 147210 674580
rect 147300 674340 147540 674580
rect 147630 674340 147870 674580
rect 147980 674340 148220 674580
rect 148310 674340 148550 674580
rect 148640 674340 148880 674580
rect 148970 674340 149210 674580
rect 149320 674340 149560 674580
rect 149650 674340 149890 674580
rect 149980 674340 150220 674580
rect 150310 674340 150550 674580
rect 150660 674340 150900 674580
rect 150990 674340 151230 674580
rect 151320 674340 151560 674580
rect 151650 674340 151890 674580
rect 152000 674340 152240 674580
rect 152330 674340 152570 674580
rect 152660 674340 152900 674580
rect 152990 674340 153230 674580
rect 153340 674340 153580 674580
rect 153670 674340 153910 674580
rect 154000 674340 154240 674580
rect 154330 674340 154570 674580
rect 154680 674340 154920 674580
rect 155010 674340 155250 674580
rect 155340 674340 155580 674580
rect 155670 674340 155910 674580
rect 144950 674010 145190 674250
rect 145300 674010 145540 674250
rect 145630 674010 145870 674250
rect 145960 674010 146200 674250
rect 146290 674010 146530 674250
rect 146640 674010 146880 674250
rect 146970 674010 147210 674250
rect 147300 674010 147540 674250
rect 147630 674010 147870 674250
rect 147980 674010 148220 674250
rect 148310 674010 148550 674250
rect 148640 674010 148880 674250
rect 148970 674010 149210 674250
rect 149320 674010 149560 674250
rect 149650 674010 149890 674250
rect 149980 674010 150220 674250
rect 150310 674010 150550 674250
rect 150660 674010 150900 674250
rect 150990 674010 151230 674250
rect 151320 674010 151560 674250
rect 151650 674010 151890 674250
rect 152000 674010 152240 674250
rect 152330 674010 152570 674250
rect 152660 674010 152900 674250
rect 152990 674010 153230 674250
rect 153340 674010 153580 674250
rect 153670 674010 153910 674250
rect 154000 674010 154240 674250
rect 154330 674010 154570 674250
rect 154680 674010 154920 674250
rect 155010 674010 155250 674250
rect 155340 674010 155580 674250
rect 155670 674010 155910 674250
rect 144950 673660 145190 673900
rect 145300 673660 145540 673900
rect 145630 673660 145870 673900
rect 145960 673660 146200 673900
rect 146290 673660 146530 673900
rect 146640 673660 146880 673900
rect 146970 673660 147210 673900
rect 147300 673660 147540 673900
rect 147630 673660 147870 673900
rect 147980 673660 148220 673900
rect 148310 673660 148550 673900
rect 148640 673660 148880 673900
rect 148970 673660 149210 673900
rect 149320 673660 149560 673900
rect 149650 673660 149890 673900
rect 149980 673660 150220 673900
rect 150310 673660 150550 673900
rect 150660 673660 150900 673900
rect 150990 673660 151230 673900
rect 151320 673660 151560 673900
rect 151650 673660 151890 673900
rect 152000 673660 152240 673900
rect 152330 673660 152570 673900
rect 152660 673660 152900 673900
rect 152990 673660 153230 673900
rect 153340 673660 153580 673900
rect 153670 673660 153910 673900
rect 154000 673660 154240 673900
rect 154330 673660 154570 673900
rect 154680 673660 154920 673900
rect 155010 673660 155250 673900
rect 155340 673660 155580 673900
rect 155670 673660 155910 673900
rect 144950 673330 145190 673570
rect 145300 673330 145540 673570
rect 145630 673330 145870 673570
rect 145960 673330 146200 673570
rect 146290 673330 146530 673570
rect 146640 673330 146880 673570
rect 146970 673330 147210 673570
rect 147300 673330 147540 673570
rect 147630 673330 147870 673570
rect 147980 673330 148220 673570
rect 148310 673330 148550 673570
rect 148640 673330 148880 673570
rect 148970 673330 149210 673570
rect 149320 673330 149560 673570
rect 149650 673330 149890 673570
rect 149980 673330 150220 673570
rect 150310 673330 150550 673570
rect 150660 673330 150900 673570
rect 150990 673330 151230 673570
rect 151320 673330 151560 673570
rect 151650 673330 151890 673570
rect 152000 673330 152240 673570
rect 152330 673330 152570 673570
rect 152660 673330 152900 673570
rect 152990 673330 153230 673570
rect 153340 673330 153580 673570
rect 153670 673330 153910 673570
rect 154000 673330 154240 673570
rect 154330 673330 154570 673570
rect 154680 673330 154920 673570
rect 155010 673330 155250 673570
rect 155340 673330 155580 673570
rect 155670 673330 155910 673570
rect 144950 673000 145190 673240
rect 145300 673000 145540 673240
rect 145630 673000 145870 673240
rect 145960 673000 146200 673240
rect 146290 673000 146530 673240
rect 146640 673000 146880 673240
rect 146970 673000 147210 673240
rect 147300 673000 147540 673240
rect 147630 673000 147870 673240
rect 147980 673000 148220 673240
rect 148310 673000 148550 673240
rect 148640 673000 148880 673240
rect 148970 673000 149210 673240
rect 149320 673000 149560 673240
rect 149650 673000 149890 673240
rect 149980 673000 150220 673240
rect 150310 673000 150550 673240
rect 150660 673000 150900 673240
rect 150990 673000 151230 673240
rect 151320 673000 151560 673240
rect 151650 673000 151890 673240
rect 152000 673000 152240 673240
rect 152330 673000 152570 673240
rect 152660 673000 152900 673240
rect 152990 673000 153230 673240
rect 153340 673000 153580 673240
rect 153670 673000 153910 673240
rect 154000 673000 154240 673240
rect 154330 673000 154570 673240
rect 154680 673000 154920 673240
rect 155010 673000 155250 673240
rect 155340 673000 155580 673240
rect 155670 673000 155910 673240
rect 144950 672670 145190 672910
rect 145300 672670 145540 672910
rect 145630 672670 145870 672910
rect 145960 672670 146200 672910
rect 146290 672670 146530 672910
rect 146640 672670 146880 672910
rect 146970 672670 147210 672910
rect 147300 672670 147540 672910
rect 147630 672670 147870 672910
rect 147980 672670 148220 672910
rect 148310 672670 148550 672910
rect 148640 672670 148880 672910
rect 148970 672670 149210 672910
rect 149320 672670 149560 672910
rect 149650 672670 149890 672910
rect 149980 672670 150220 672910
rect 150310 672670 150550 672910
rect 150660 672670 150900 672910
rect 150990 672670 151230 672910
rect 151320 672670 151560 672910
rect 151650 672670 151890 672910
rect 152000 672670 152240 672910
rect 152330 672670 152570 672910
rect 152660 672670 152900 672910
rect 152990 672670 153230 672910
rect 153340 672670 153580 672910
rect 153670 672670 153910 672910
rect 154000 672670 154240 672910
rect 154330 672670 154570 672910
rect 154680 672670 154920 672910
rect 155010 672670 155250 672910
rect 155340 672670 155580 672910
rect 155670 672670 155910 672910
rect 144950 672320 145190 672560
rect 145300 672320 145540 672560
rect 145630 672320 145870 672560
rect 145960 672320 146200 672560
rect 146290 672320 146530 672560
rect 146640 672320 146880 672560
rect 146970 672320 147210 672560
rect 147300 672320 147540 672560
rect 147630 672320 147870 672560
rect 147980 672320 148220 672560
rect 148310 672320 148550 672560
rect 148640 672320 148880 672560
rect 148970 672320 149210 672560
rect 149320 672320 149560 672560
rect 149650 672320 149890 672560
rect 149980 672320 150220 672560
rect 150310 672320 150550 672560
rect 150660 672320 150900 672560
rect 150990 672320 151230 672560
rect 151320 672320 151560 672560
rect 151650 672320 151890 672560
rect 152000 672320 152240 672560
rect 152330 672320 152570 672560
rect 152660 672320 152900 672560
rect 152990 672320 153230 672560
rect 153340 672320 153580 672560
rect 153670 672320 153910 672560
rect 154000 672320 154240 672560
rect 154330 672320 154570 672560
rect 154680 672320 154920 672560
rect 155010 672320 155250 672560
rect 155340 672320 155580 672560
rect 155670 672320 155910 672560
rect 110810 671660 111050 671900
rect 111140 671660 111380 671900
rect 111470 671660 111710 671900
rect 111800 671660 112040 671900
rect 112150 671660 112390 671900
rect 112480 671660 112720 671900
rect 112810 671660 113050 671900
rect 113140 671660 113380 671900
rect 113490 671660 113730 671900
rect 113820 671660 114060 671900
rect 114150 671660 114390 671900
rect 114480 671660 114720 671900
rect 114830 671660 115070 671900
rect 115160 671660 115400 671900
rect 115490 671660 115730 671900
rect 115820 671660 116060 671900
rect 116170 671660 116410 671900
rect 116500 671660 116740 671900
rect 116830 671660 117070 671900
rect 117160 671660 117400 671900
rect 117510 671660 117750 671900
rect 117840 671660 118080 671900
rect 118170 671660 118410 671900
rect 118500 671660 118740 671900
rect 118850 671660 119090 671900
rect 119180 671660 119420 671900
rect 119510 671660 119750 671900
rect 119840 671660 120080 671900
rect 120190 671660 120430 671900
rect 120520 671660 120760 671900
rect 120850 671660 121090 671900
rect 121180 671660 121420 671900
rect 121530 671660 121770 671900
rect 110810 671310 111050 671550
rect 111140 671310 111380 671550
rect 111470 671310 111710 671550
rect 111800 671310 112040 671550
rect 112150 671310 112390 671550
rect 112480 671310 112720 671550
rect 112810 671310 113050 671550
rect 113140 671310 113380 671550
rect 113490 671310 113730 671550
rect 113820 671310 114060 671550
rect 114150 671310 114390 671550
rect 114480 671310 114720 671550
rect 114830 671310 115070 671550
rect 115160 671310 115400 671550
rect 115490 671310 115730 671550
rect 115820 671310 116060 671550
rect 116170 671310 116410 671550
rect 116500 671310 116740 671550
rect 116830 671310 117070 671550
rect 117160 671310 117400 671550
rect 117510 671310 117750 671550
rect 117840 671310 118080 671550
rect 118170 671310 118410 671550
rect 118500 671310 118740 671550
rect 118850 671310 119090 671550
rect 119180 671310 119420 671550
rect 119510 671310 119750 671550
rect 119840 671310 120080 671550
rect 120190 671310 120430 671550
rect 120520 671310 120760 671550
rect 120850 671310 121090 671550
rect 121180 671310 121420 671550
rect 121530 671310 121770 671550
rect 110810 670980 111050 671220
rect 111140 670980 111380 671220
rect 111470 670980 111710 671220
rect 111800 670980 112040 671220
rect 112150 670980 112390 671220
rect 112480 670980 112720 671220
rect 112810 670980 113050 671220
rect 113140 670980 113380 671220
rect 113490 670980 113730 671220
rect 113820 670980 114060 671220
rect 114150 670980 114390 671220
rect 114480 670980 114720 671220
rect 114830 670980 115070 671220
rect 115160 670980 115400 671220
rect 115490 670980 115730 671220
rect 115820 670980 116060 671220
rect 116170 670980 116410 671220
rect 116500 670980 116740 671220
rect 116830 670980 117070 671220
rect 117160 670980 117400 671220
rect 117510 670980 117750 671220
rect 117840 670980 118080 671220
rect 118170 670980 118410 671220
rect 118500 670980 118740 671220
rect 118850 670980 119090 671220
rect 119180 670980 119420 671220
rect 119510 670980 119750 671220
rect 119840 670980 120080 671220
rect 120190 670980 120430 671220
rect 120520 670980 120760 671220
rect 120850 670980 121090 671220
rect 121180 670980 121420 671220
rect 121530 670980 121770 671220
rect 110810 670650 111050 670890
rect 111140 670650 111380 670890
rect 111470 670650 111710 670890
rect 111800 670650 112040 670890
rect 112150 670650 112390 670890
rect 112480 670650 112720 670890
rect 112810 670650 113050 670890
rect 113140 670650 113380 670890
rect 113490 670650 113730 670890
rect 113820 670650 114060 670890
rect 114150 670650 114390 670890
rect 114480 670650 114720 670890
rect 114830 670650 115070 670890
rect 115160 670650 115400 670890
rect 115490 670650 115730 670890
rect 115820 670650 116060 670890
rect 116170 670650 116410 670890
rect 116500 670650 116740 670890
rect 116830 670650 117070 670890
rect 117160 670650 117400 670890
rect 117510 670650 117750 670890
rect 117840 670650 118080 670890
rect 118170 670650 118410 670890
rect 118500 670650 118740 670890
rect 118850 670650 119090 670890
rect 119180 670650 119420 670890
rect 119510 670650 119750 670890
rect 119840 670650 120080 670890
rect 120190 670650 120430 670890
rect 120520 670650 120760 670890
rect 120850 670650 121090 670890
rect 121180 670650 121420 670890
rect 121530 670650 121770 670890
rect 110810 670320 111050 670560
rect 111140 670320 111380 670560
rect 111470 670320 111710 670560
rect 111800 670320 112040 670560
rect 112150 670320 112390 670560
rect 112480 670320 112720 670560
rect 112810 670320 113050 670560
rect 113140 670320 113380 670560
rect 113490 670320 113730 670560
rect 113820 670320 114060 670560
rect 114150 670320 114390 670560
rect 114480 670320 114720 670560
rect 114830 670320 115070 670560
rect 115160 670320 115400 670560
rect 115490 670320 115730 670560
rect 115820 670320 116060 670560
rect 116170 670320 116410 670560
rect 116500 670320 116740 670560
rect 116830 670320 117070 670560
rect 117160 670320 117400 670560
rect 117510 670320 117750 670560
rect 117840 670320 118080 670560
rect 118170 670320 118410 670560
rect 118500 670320 118740 670560
rect 118850 670320 119090 670560
rect 119180 670320 119420 670560
rect 119510 670320 119750 670560
rect 119840 670320 120080 670560
rect 120190 670320 120430 670560
rect 120520 670320 120760 670560
rect 120850 670320 121090 670560
rect 121180 670320 121420 670560
rect 121530 670320 121770 670560
rect 110810 669970 111050 670210
rect 111140 669970 111380 670210
rect 111470 669970 111710 670210
rect 111800 669970 112040 670210
rect 112150 669970 112390 670210
rect 112480 669970 112720 670210
rect 112810 669970 113050 670210
rect 113140 669970 113380 670210
rect 113490 669970 113730 670210
rect 113820 669970 114060 670210
rect 114150 669970 114390 670210
rect 114480 669970 114720 670210
rect 114830 669970 115070 670210
rect 115160 669970 115400 670210
rect 115490 669970 115730 670210
rect 115820 669970 116060 670210
rect 116170 669970 116410 670210
rect 116500 669970 116740 670210
rect 116830 669970 117070 670210
rect 117160 669970 117400 670210
rect 117510 669970 117750 670210
rect 117840 669970 118080 670210
rect 118170 669970 118410 670210
rect 118500 669970 118740 670210
rect 118850 669970 119090 670210
rect 119180 669970 119420 670210
rect 119510 669970 119750 670210
rect 119840 669970 120080 670210
rect 120190 669970 120430 670210
rect 120520 669970 120760 670210
rect 120850 669970 121090 670210
rect 121180 669970 121420 670210
rect 121530 669970 121770 670210
rect 110810 669640 111050 669880
rect 111140 669640 111380 669880
rect 111470 669640 111710 669880
rect 111800 669640 112040 669880
rect 112150 669640 112390 669880
rect 112480 669640 112720 669880
rect 112810 669640 113050 669880
rect 113140 669640 113380 669880
rect 113490 669640 113730 669880
rect 113820 669640 114060 669880
rect 114150 669640 114390 669880
rect 114480 669640 114720 669880
rect 114830 669640 115070 669880
rect 115160 669640 115400 669880
rect 115490 669640 115730 669880
rect 115820 669640 116060 669880
rect 116170 669640 116410 669880
rect 116500 669640 116740 669880
rect 116830 669640 117070 669880
rect 117160 669640 117400 669880
rect 117510 669640 117750 669880
rect 117840 669640 118080 669880
rect 118170 669640 118410 669880
rect 118500 669640 118740 669880
rect 118850 669640 119090 669880
rect 119180 669640 119420 669880
rect 119510 669640 119750 669880
rect 119840 669640 120080 669880
rect 120190 669640 120430 669880
rect 120520 669640 120760 669880
rect 120850 669640 121090 669880
rect 121180 669640 121420 669880
rect 121530 669640 121770 669880
rect 110810 669310 111050 669550
rect 111140 669310 111380 669550
rect 111470 669310 111710 669550
rect 111800 669310 112040 669550
rect 112150 669310 112390 669550
rect 112480 669310 112720 669550
rect 112810 669310 113050 669550
rect 113140 669310 113380 669550
rect 113490 669310 113730 669550
rect 113820 669310 114060 669550
rect 114150 669310 114390 669550
rect 114480 669310 114720 669550
rect 114830 669310 115070 669550
rect 115160 669310 115400 669550
rect 115490 669310 115730 669550
rect 115820 669310 116060 669550
rect 116170 669310 116410 669550
rect 116500 669310 116740 669550
rect 116830 669310 117070 669550
rect 117160 669310 117400 669550
rect 117510 669310 117750 669550
rect 117840 669310 118080 669550
rect 118170 669310 118410 669550
rect 118500 669310 118740 669550
rect 118850 669310 119090 669550
rect 119180 669310 119420 669550
rect 119510 669310 119750 669550
rect 119840 669310 120080 669550
rect 120190 669310 120430 669550
rect 120520 669310 120760 669550
rect 120850 669310 121090 669550
rect 121180 669310 121420 669550
rect 121530 669310 121770 669550
rect 110810 668980 111050 669220
rect 111140 668980 111380 669220
rect 111470 668980 111710 669220
rect 111800 668980 112040 669220
rect 112150 668980 112390 669220
rect 112480 668980 112720 669220
rect 112810 668980 113050 669220
rect 113140 668980 113380 669220
rect 113490 668980 113730 669220
rect 113820 668980 114060 669220
rect 114150 668980 114390 669220
rect 114480 668980 114720 669220
rect 114830 668980 115070 669220
rect 115160 668980 115400 669220
rect 115490 668980 115730 669220
rect 115820 668980 116060 669220
rect 116170 668980 116410 669220
rect 116500 668980 116740 669220
rect 116830 668980 117070 669220
rect 117160 668980 117400 669220
rect 117510 668980 117750 669220
rect 117840 668980 118080 669220
rect 118170 668980 118410 669220
rect 118500 668980 118740 669220
rect 118850 668980 119090 669220
rect 119180 668980 119420 669220
rect 119510 668980 119750 669220
rect 119840 668980 120080 669220
rect 120190 668980 120430 669220
rect 120520 668980 120760 669220
rect 120850 668980 121090 669220
rect 121180 668980 121420 669220
rect 121530 668980 121770 669220
rect 110810 668630 111050 668870
rect 111140 668630 111380 668870
rect 111470 668630 111710 668870
rect 111800 668630 112040 668870
rect 112150 668630 112390 668870
rect 112480 668630 112720 668870
rect 112810 668630 113050 668870
rect 113140 668630 113380 668870
rect 113490 668630 113730 668870
rect 113820 668630 114060 668870
rect 114150 668630 114390 668870
rect 114480 668630 114720 668870
rect 114830 668630 115070 668870
rect 115160 668630 115400 668870
rect 115490 668630 115730 668870
rect 115820 668630 116060 668870
rect 116170 668630 116410 668870
rect 116500 668630 116740 668870
rect 116830 668630 117070 668870
rect 117160 668630 117400 668870
rect 117510 668630 117750 668870
rect 117840 668630 118080 668870
rect 118170 668630 118410 668870
rect 118500 668630 118740 668870
rect 118850 668630 119090 668870
rect 119180 668630 119420 668870
rect 119510 668630 119750 668870
rect 119840 668630 120080 668870
rect 120190 668630 120430 668870
rect 120520 668630 120760 668870
rect 120850 668630 121090 668870
rect 121180 668630 121420 668870
rect 121530 668630 121770 668870
rect 110810 668300 111050 668540
rect 111140 668300 111380 668540
rect 111470 668300 111710 668540
rect 111800 668300 112040 668540
rect 112150 668300 112390 668540
rect 112480 668300 112720 668540
rect 112810 668300 113050 668540
rect 113140 668300 113380 668540
rect 113490 668300 113730 668540
rect 113820 668300 114060 668540
rect 114150 668300 114390 668540
rect 114480 668300 114720 668540
rect 114830 668300 115070 668540
rect 115160 668300 115400 668540
rect 115490 668300 115730 668540
rect 115820 668300 116060 668540
rect 116170 668300 116410 668540
rect 116500 668300 116740 668540
rect 116830 668300 117070 668540
rect 117160 668300 117400 668540
rect 117510 668300 117750 668540
rect 117840 668300 118080 668540
rect 118170 668300 118410 668540
rect 118500 668300 118740 668540
rect 118850 668300 119090 668540
rect 119180 668300 119420 668540
rect 119510 668300 119750 668540
rect 119840 668300 120080 668540
rect 120190 668300 120430 668540
rect 120520 668300 120760 668540
rect 120850 668300 121090 668540
rect 121180 668300 121420 668540
rect 121530 668300 121770 668540
rect 110810 667970 111050 668210
rect 111140 667970 111380 668210
rect 111470 667970 111710 668210
rect 111800 667970 112040 668210
rect 112150 667970 112390 668210
rect 112480 667970 112720 668210
rect 112810 667970 113050 668210
rect 113140 667970 113380 668210
rect 113490 667970 113730 668210
rect 113820 667970 114060 668210
rect 114150 667970 114390 668210
rect 114480 667970 114720 668210
rect 114830 667970 115070 668210
rect 115160 667970 115400 668210
rect 115490 667970 115730 668210
rect 115820 667970 116060 668210
rect 116170 667970 116410 668210
rect 116500 667970 116740 668210
rect 116830 667970 117070 668210
rect 117160 667970 117400 668210
rect 117510 667970 117750 668210
rect 117840 667970 118080 668210
rect 118170 667970 118410 668210
rect 118500 667970 118740 668210
rect 118850 667970 119090 668210
rect 119180 667970 119420 668210
rect 119510 667970 119750 668210
rect 119840 667970 120080 668210
rect 120190 667970 120430 668210
rect 120520 667970 120760 668210
rect 120850 667970 121090 668210
rect 121180 667970 121420 668210
rect 121530 667970 121770 668210
rect 110810 667640 111050 667880
rect 111140 667640 111380 667880
rect 111470 667640 111710 667880
rect 111800 667640 112040 667880
rect 112150 667640 112390 667880
rect 112480 667640 112720 667880
rect 112810 667640 113050 667880
rect 113140 667640 113380 667880
rect 113490 667640 113730 667880
rect 113820 667640 114060 667880
rect 114150 667640 114390 667880
rect 114480 667640 114720 667880
rect 114830 667640 115070 667880
rect 115160 667640 115400 667880
rect 115490 667640 115730 667880
rect 115820 667640 116060 667880
rect 116170 667640 116410 667880
rect 116500 667640 116740 667880
rect 116830 667640 117070 667880
rect 117160 667640 117400 667880
rect 117510 667640 117750 667880
rect 117840 667640 118080 667880
rect 118170 667640 118410 667880
rect 118500 667640 118740 667880
rect 118850 667640 119090 667880
rect 119180 667640 119420 667880
rect 119510 667640 119750 667880
rect 119840 667640 120080 667880
rect 120190 667640 120430 667880
rect 120520 667640 120760 667880
rect 120850 667640 121090 667880
rect 121180 667640 121420 667880
rect 121530 667640 121770 667880
rect 110810 667290 111050 667530
rect 111140 667290 111380 667530
rect 111470 667290 111710 667530
rect 111800 667290 112040 667530
rect 112150 667290 112390 667530
rect 112480 667290 112720 667530
rect 112810 667290 113050 667530
rect 113140 667290 113380 667530
rect 113490 667290 113730 667530
rect 113820 667290 114060 667530
rect 114150 667290 114390 667530
rect 114480 667290 114720 667530
rect 114830 667290 115070 667530
rect 115160 667290 115400 667530
rect 115490 667290 115730 667530
rect 115820 667290 116060 667530
rect 116170 667290 116410 667530
rect 116500 667290 116740 667530
rect 116830 667290 117070 667530
rect 117160 667290 117400 667530
rect 117510 667290 117750 667530
rect 117840 667290 118080 667530
rect 118170 667290 118410 667530
rect 118500 667290 118740 667530
rect 118850 667290 119090 667530
rect 119180 667290 119420 667530
rect 119510 667290 119750 667530
rect 119840 667290 120080 667530
rect 120190 667290 120430 667530
rect 120520 667290 120760 667530
rect 120850 667290 121090 667530
rect 121180 667290 121420 667530
rect 121530 667290 121770 667530
rect 110810 666960 111050 667200
rect 111140 666960 111380 667200
rect 111470 666960 111710 667200
rect 111800 666960 112040 667200
rect 112150 666960 112390 667200
rect 112480 666960 112720 667200
rect 112810 666960 113050 667200
rect 113140 666960 113380 667200
rect 113490 666960 113730 667200
rect 113820 666960 114060 667200
rect 114150 666960 114390 667200
rect 114480 666960 114720 667200
rect 114830 666960 115070 667200
rect 115160 666960 115400 667200
rect 115490 666960 115730 667200
rect 115820 666960 116060 667200
rect 116170 666960 116410 667200
rect 116500 666960 116740 667200
rect 116830 666960 117070 667200
rect 117160 666960 117400 667200
rect 117510 666960 117750 667200
rect 117840 666960 118080 667200
rect 118170 666960 118410 667200
rect 118500 666960 118740 667200
rect 118850 666960 119090 667200
rect 119180 666960 119420 667200
rect 119510 666960 119750 667200
rect 119840 666960 120080 667200
rect 120190 666960 120430 667200
rect 120520 666960 120760 667200
rect 120850 666960 121090 667200
rect 121180 666960 121420 667200
rect 121530 666960 121770 667200
rect 110810 666630 111050 666870
rect 111140 666630 111380 666870
rect 111470 666630 111710 666870
rect 111800 666630 112040 666870
rect 112150 666630 112390 666870
rect 112480 666630 112720 666870
rect 112810 666630 113050 666870
rect 113140 666630 113380 666870
rect 113490 666630 113730 666870
rect 113820 666630 114060 666870
rect 114150 666630 114390 666870
rect 114480 666630 114720 666870
rect 114830 666630 115070 666870
rect 115160 666630 115400 666870
rect 115490 666630 115730 666870
rect 115820 666630 116060 666870
rect 116170 666630 116410 666870
rect 116500 666630 116740 666870
rect 116830 666630 117070 666870
rect 117160 666630 117400 666870
rect 117510 666630 117750 666870
rect 117840 666630 118080 666870
rect 118170 666630 118410 666870
rect 118500 666630 118740 666870
rect 118850 666630 119090 666870
rect 119180 666630 119420 666870
rect 119510 666630 119750 666870
rect 119840 666630 120080 666870
rect 120190 666630 120430 666870
rect 120520 666630 120760 666870
rect 120850 666630 121090 666870
rect 121180 666630 121420 666870
rect 121530 666630 121770 666870
rect 110810 666300 111050 666540
rect 111140 666300 111380 666540
rect 111470 666300 111710 666540
rect 111800 666300 112040 666540
rect 112150 666300 112390 666540
rect 112480 666300 112720 666540
rect 112810 666300 113050 666540
rect 113140 666300 113380 666540
rect 113490 666300 113730 666540
rect 113820 666300 114060 666540
rect 114150 666300 114390 666540
rect 114480 666300 114720 666540
rect 114830 666300 115070 666540
rect 115160 666300 115400 666540
rect 115490 666300 115730 666540
rect 115820 666300 116060 666540
rect 116170 666300 116410 666540
rect 116500 666300 116740 666540
rect 116830 666300 117070 666540
rect 117160 666300 117400 666540
rect 117510 666300 117750 666540
rect 117840 666300 118080 666540
rect 118170 666300 118410 666540
rect 118500 666300 118740 666540
rect 118850 666300 119090 666540
rect 119180 666300 119420 666540
rect 119510 666300 119750 666540
rect 119840 666300 120080 666540
rect 120190 666300 120430 666540
rect 120520 666300 120760 666540
rect 120850 666300 121090 666540
rect 121180 666300 121420 666540
rect 121530 666300 121770 666540
rect 110810 665950 111050 666190
rect 111140 665950 111380 666190
rect 111470 665950 111710 666190
rect 111800 665950 112040 666190
rect 112150 665950 112390 666190
rect 112480 665950 112720 666190
rect 112810 665950 113050 666190
rect 113140 665950 113380 666190
rect 113490 665950 113730 666190
rect 113820 665950 114060 666190
rect 114150 665950 114390 666190
rect 114480 665950 114720 666190
rect 114830 665950 115070 666190
rect 115160 665950 115400 666190
rect 115490 665950 115730 666190
rect 115820 665950 116060 666190
rect 116170 665950 116410 666190
rect 116500 665950 116740 666190
rect 116830 665950 117070 666190
rect 117160 665950 117400 666190
rect 117510 665950 117750 666190
rect 117840 665950 118080 666190
rect 118170 665950 118410 666190
rect 118500 665950 118740 666190
rect 118850 665950 119090 666190
rect 119180 665950 119420 666190
rect 119510 665950 119750 666190
rect 119840 665950 120080 666190
rect 120190 665950 120430 666190
rect 120520 665950 120760 666190
rect 120850 665950 121090 666190
rect 121180 665950 121420 666190
rect 121530 665950 121770 666190
rect 110810 665620 111050 665860
rect 111140 665620 111380 665860
rect 111470 665620 111710 665860
rect 111800 665620 112040 665860
rect 112150 665620 112390 665860
rect 112480 665620 112720 665860
rect 112810 665620 113050 665860
rect 113140 665620 113380 665860
rect 113490 665620 113730 665860
rect 113820 665620 114060 665860
rect 114150 665620 114390 665860
rect 114480 665620 114720 665860
rect 114830 665620 115070 665860
rect 115160 665620 115400 665860
rect 115490 665620 115730 665860
rect 115820 665620 116060 665860
rect 116170 665620 116410 665860
rect 116500 665620 116740 665860
rect 116830 665620 117070 665860
rect 117160 665620 117400 665860
rect 117510 665620 117750 665860
rect 117840 665620 118080 665860
rect 118170 665620 118410 665860
rect 118500 665620 118740 665860
rect 118850 665620 119090 665860
rect 119180 665620 119420 665860
rect 119510 665620 119750 665860
rect 119840 665620 120080 665860
rect 120190 665620 120430 665860
rect 120520 665620 120760 665860
rect 120850 665620 121090 665860
rect 121180 665620 121420 665860
rect 121530 665620 121770 665860
rect 110810 665290 111050 665530
rect 111140 665290 111380 665530
rect 111470 665290 111710 665530
rect 111800 665290 112040 665530
rect 112150 665290 112390 665530
rect 112480 665290 112720 665530
rect 112810 665290 113050 665530
rect 113140 665290 113380 665530
rect 113490 665290 113730 665530
rect 113820 665290 114060 665530
rect 114150 665290 114390 665530
rect 114480 665290 114720 665530
rect 114830 665290 115070 665530
rect 115160 665290 115400 665530
rect 115490 665290 115730 665530
rect 115820 665290 116060 665530
rect 116170 665290 116410 665530
rect 116500 665290 116740 665530
rect 116830 665290 117070 665530
rect 117160 665290 117400 665530
rect 117510 665290 117750 665530
rect 117840 665290 118080 665530
rect 118170 665290 118410 665530
rect 118500 665290 118740 665530
rect 118850 665290 119090 665530
rect 119180 665290 119420 665530
rect 119510 665290 119750 665530
rect 119840 665290 120080 665530
rect 120190 665290 120430 665530
rect 120520 665290 120760 665530
rect 120850 665290 121090 665530
rect 121180 665290 121420 665530
rect 121530 665290 121770 665530
rect 110810 664960 111050 665200
rect 111140 664960 111380 665200
rect 111470 664960 111710 665200
rect 111800 664960 112040 665200
rect 112150 664960 112390 665200
rect 112480 664960 112720 665200
rect 112810 664960 113050 665200
rect 113140 664960 113380 665200
rect 113490 664960 113730 665200
rect 113820 664960 114060 665200
rect 114150 664960 114390 665200
rect 114480 664960 114720 665200
rect 114830 664960 115070 665200
rect 115160 664960 115400 665200
rect 115490 664960 115730 665200
rect 115820 664960 116060 665200
rect 116170 664960 116410 665200
rect 116500 664960 116740 665200
rect 116830 664960 117070 665200
rect 117160 664960 117400 665200
rect 117510 664960 117750 665200
rect 117840 664960 118080 665200
rect 118170 664960 118410 665200
rect 118500 664960 118740 665200
rect 118850 664960 119090 665200
rect 119180 664960 119420 665200
rect 119510 664960 119750 665200
rect 119840 664960 120080 665200
rect 120190 664960 120430 665200
rect 120520 664960 120760 665200
rect 120850 664960 121090 665200
rect 121180 664960 121420 665200
rect 121530 664960 121770 665200
rect 110810 664610 111050 664850
rect 111140 664610 111380 664850
rect 111470 664610 111710 664850
rect 111800 664610 112040 664850
rect 112150 664610 112390 664850
rect 112480 664610 112720 664850
rect 112810 664610 113050 664850
rect 113140 664610 113380 664850
rect 113490 664610 113730 664850
rect 113820 664610 114060 664850
rect 114150 664610 114390 664850
rect 114480 664610 114720 664850
rect 114830 664610 115070 664850
rect 115160 664610 115400 664850
rect 115490 664610 115730 664850
rect 115820 664610 116060 664850
rect 116170 664610 116410 664850
rect 116500 664610 116740 664850
rect 116830 664610 117070 664850
rect 117160 664610 117400 664850
rect 117510 664610 117750 664850
rect 117840 664610 118080 664850
rect 118170 664610 118410 664850
rect 118500 664610 118740 664850
rect 118850 664610 119090 664850
rect 119180 664610 119420 664850
rect 119510 664610 119750 664850
rect 119840 664610 120080 664850
rect 120190 664610 120430 664850
rect 120520 664610 120760 664850
rect 120850 664610 121090 664850
rect 121180 664610 121420 664850
rect 121530 664610 121770 664850
rect 110810 664280 111050 664520
rect 111140 664280 111380 664520
rect 111470 664280 111710 664520
rect 111800 664280 112040 664520
rect 112150 664280 112390 664520
rect 112480 664280 112720 664520
rect 112810 664280 113050 664520
rect 113140 664280 113380 664520
rect 113490 664280 113730 664520
rect 113820 664280 114060 664520
rect 114150 664280 114390 664520
rect 114480 664280 114720 664520
rect 114830 664280 115070 664520
rect 115160 664280 115400 664520
rect 115490 664280 115730 664520
rect 115820 664280 116060 664520
rect 116170 664280 116410 664520
rect 116500 664280 116740 664520
rect 116830 664280 117070 664520
rect 117160 664280 117400 664520
rect 117510 664280 117750 664520
rect 117840 664280 118080 664520
rect 118170 664280 118410 664520
rect 118500 664280 118740 664520
rect 118850 664280 119090 664520
rect 119180 664280 119420 664520
rect 119510 664280 119750 664520
rect 119840 664280 120080 664520
rect 120190 664280 120430 664520
rect 120520 664280 120760 664520
rect 120850 664280 121090 664520
rect 121180 664280 121420 664520
rect 121530 664280 121770 664520
rect 110810 663950 111050 664190
rect 111140 663950 111380 664190
rect 111470 663950 111710 664190
rect 111800 663950 112040 664190
rect 112150 663950 112390 664190
rect 112480 663950 112720 664190
rect 112810 663950 113050 664190
rect 113140 663950 113380 664190
rect 113490 663950 113730 664190
rect 113820 663950 114060 664190
rect 114150 663950 114390 664190
rect 114480 663950 114720 664190
rect 114830 663950 115070 664190
rect 115160 663950 115400 664190
rect 115490 663950 115730 664190
rect 115820 663950 116060 664190
rect 116170 663950 116410 664190
rect 116500 663950 116740 664190
rect 116830 663950 117070 664190
rect 117160 663950 117400 664190
rect 117510 663950 117750 664190
rect 117840 663950 118080 664190
rect 118170 663950 118410 664190
rect 118500 663950 118740 664190
rect 118850 663950 119090 664190
rect 119180 663950 119420 664190
rect 119510 663950 119750 664190
rect 119840 663950 120080 664190
rect 120190 663950 120430 664190
rect 120520 663950 120760 664190
rect 120850 663950 121090 664190
rect 121180 663950 121420 664190
rect 121530 663950 121770 664190
rect 110810 663620 111050 663860
rect 111140 663620 111380 663860
rect 111470 663620 111710 663860
rect 111800 663620 112040 663860
rect 112150 663620 112390 663860
rect 112480 663620 112720 663860
rect 112810 663620 113050 663860
rect 113140 663620 113380 663860
rect 113490 663620 113730 663860
rect 113820 663620 114060 663860
rect 114150 663620 114390 663860
rect 114480 663620 114720 663860
rect 114830 663620 115070 663860
rect 115160 663620 115400 663860
rect 115490 663620 115730 663860
rect 115820 663620 116060 663860
rect 116170 663620 116410 663860
rect 116500 663620 116740 663860
rect 116830 663620 117070 663860
rect 117160 663620 117400 663860
rect 117510 663620 117750 663860
rect 117840 663620 118080 663860
rect 118170 663620 118410 663860
rect 118500 663620 118740 663860
rect 118850 663620 119090 663860
rect 119180 663620 119420 663860
rect 119510 663620 119750 663860
rect 119840 663620 120080 663860
rect 120190 663620 120430 663860
rect 120520 663620 120760 663860
rect 120850 663620 121090 663860
rect 121180 663620 121420 663860
rect 121530 663620 121770 663860
rect 110810 663270 111050 663510
rect 111140 663270 111380 663510
rect 111470 663270 111710 663510
rect 111800 663270 112040 663510
rect 112150 663270 112390 663510
rect 112480 663270 112720 663510
rect 112810 663270 113050 663510
rect 113140 663270 113380 663510
rect 113490 663270 113730 663510
rect 113820 663270 114060 663510
rect 114150 663270 114390 663510
rect 114480 663270 114720 663510
rect 114830 663270 115070 663510
rect 115160 663270 115400 663510
rect 115490 663270 115730 663510
rect 115820 663270 116060 663510
rect 116170 663270 116410 663510
rect 116500 663270 116740 663510
rect 116830 663270 117070 663510
rect 117160 663270 117400 663510
rect 117510 663270 117750 663510
rect 117840 663270 118080 663510
rect 118170 663270 118410 663510
rect 118500 663270 118740 663510
rect 118850 663270 119090 663510
rect 119180 663270 119420 663510
rect 119510 663270 119750 663510
rect 119840 663270 120080 663510
rect 120190 663270 120430 663510
rect 120520 663270 120760 663510
rect 120850 663270 121090 663510
rect 121180 663270 121420 663510
rect 121530 663270 121770 663510
rect 110810 662940 111050 663180
rect 111140 662940 111380 663180
rect 111470 662940 111710 663180
rect 111800 662940 112040 663180
rect 112150 662940 112390 663180
rect 112480 662940 112720 663180
rect 112810 662940 113050 663180
rect 113140 662940 113380 663180
rect 113490 662940 113730 663180
rect 113820 662940 114060 663180
rect 114150 662940 114390 663180
rect 114480 662940 114720 663180
rect 114830 662940 115070 663180
rect 115160 662940 115400 663180
rect 115490 662940 115730 663180
rect 115820 662940 116060 663180
rect 116170 662940 116410 663180
rect 116500 662940 116740 663180
rect 116830 662940 117070 663180
rect 117160 662940 117400 663180
rect 117510 662940 117750 663180
rect 117840 662940 118080 663180
rect 118170 662940 118410 663180
rect 118500 662940 118740 663180
rect 118850 662940 119090 663180
rect 119180 662940 119420 663180
rect 119510 662940 119750 663180
rect 119840 662940 120080 663180
rect 120190 662940 120430 663180
rect 120520 662940 120760 663180
rect 120850 662940 121090 663180
rect 121180 662940 121420 663180
rect 121530 662940 121770 663180
rect 110810 662610 111050 662850
rect 111140 662610 111380 662850
rect 111470 662610 111710 662850
rect 111800 662610 112040 662850
rect 112150 662610 112390 662850
rect 112480 662610 112720 662850
rect 112810 662610 113050 662850
rect 113140 662610 113380 662850
rect 113490 662610 113730 662850
rect 113820 662610 114060 662850
rect 114150 662610 114390 662850
rect 114480 662610 114720 662850
rect 114830 662610 115070 662850
rect 115160 662610 115400 662850
rect 115490 662610 115730 662850
rect 115820 662610 116060 662850
rect 116170 662610 116410 662850
rect 116500 662610 116740 662850
rect 116830 662610 117070 662850
rect 117160 662610 117400 662850
rect 117510 662610 117750 662850
rect 117840 662610 118080 662850
rect 118170 662610 118410 662850
rect 118500 662610 118740 662850
rect 118850 662610 119090 662850
rect 119180 662610 119420 662850
rect 119510 662610 119750 662850
rect 119840 662610 120080 662850
rect 120190 662610 120430 662850
rect 120520 662610 120760 662850
rect 120850 662610 121090 662850
rect 121180 662610 121420 662850
rect 121530 662610 121770 662850
rect 110810 662280 111050 662520
rect 111140 662280 111380 662520
rect 111470 662280 111710 662520
rect 111800 662280 112040 662520
rect 112150 662280 112390 662520
rect 112480 662280 112720 662520
rect 112810 662280 113050 662520
rect 113140 662280 113380 662520
rect 113490 662280 113730 662520
rect 113820 662280 114060 662520
rect 114150 662280 114390 662520
rect 114480 662280 114720 662520
rect 114830 662280 115070 662520
rect 115160 662280 115400 662520
rect 115490 662280 115730 662520
rect 115820 662280 116060 662520
rect 116170 662280 116410 662520
rect 116500 662280 116740 662520
rect 116830 662280 117070 662520
rect 117160 662280 117400 662520
rect 117510 662280 117750 662520
rect 117840 662280 118080 662520
rect 118170 662280 118410 662520
rect 118500 662280 118740 662520
rect 118850 662280 119090 662520
rect 119180 662280 119420 662520
rect 119510 662280 119750 662520
rect 119840 662280 120080 662520
rect 120190 662280 120430 662520
rect 120520 662280 120760 662520
rect 120850 662280 121090 662520
rect 121180 662280 121420 662520
rect 121530 662280 121770 662520
rect 110810 661930 111050 662170
rect 111140 661930 111380 662170
rect 111470 661930 111710 662170
rect 111800 661930 112040 662170
rect 112150 661930 112390 662170
rect 112480 661930 112720 662170
rect 112810 661930 113050 662170
rect 113140 661930 113380 662170
rect 113490 661930 113730 662170
rect 113820 661930 114060 662170
rect 114150 661930 114390 662170
rect 114480 661930 114720 662170
rect 114830 661930 115070 662170
rect 115160 661930 115400 662170
rect 115490 661930 115730 662170
rect 115820 661930 116060 662170
rect 116170 661930 116410 662170
rect 116500 661930 116740 662170
rect 116830 661930 117070 662170
rect 117160 661930 117400 662170
rect 117510 661930 117750 662170
rect 117840 661930 118080 662170
rect 118170 661930 118410 662170
rect 118500 661930 118740 662170
rect 118850 661930 119090 662170
rect 119180 661930 119420 662170
rect 119510 661930 119750 662170
rect 119840 661930 120080 662170
rect 120190 661930 120430 662170
rect 120520 661930 120760 662170
rect 120850 661930 121090 662170
rect 121180 661930 121420 662170
rect 121530 661930 121770 662170
rect 110810 661600 111050 661840
rect 111140 661600 111380 661840
rect 111470 661600 111710 661840
rect 111800 661600 112040 661840
rect 112150 661600 112390 661840
rect 112480 661600 112720 661840
rect 112810 661600 113050 661840
rect 113140 661600 113380 661840
rect 113490 661600 113730 661840
rect 113820 661600 114060 661840
rect 114150 661600 114390 661840
rect 114480 661600 114720 661840
rect 114830 661600 115070 661840
rect 115160 661600 115400 661840
rect 115490 661600 115730 661840
rect 115820 661600 116060 661840
rect 116170 661600 116410 661840
rect 116500 661600 116740 661840
rect 116830 661600 117070 661840
rect 117160 661600 117400 661840
rect 117510 661600 117750 661840
rect 117840 661600 118080 661840
rect 118170 661600 118410 661840
rect 118500 661600 118740 661840
rect 118850 661600 119090 661840
rect 119180 661600 119420 661840
rect 119510 661600 119750 661840
rect 119840 661600 120080 661840
rect 120190 661600 120430 661840
rect 120520 661600 120760 661840
rect 120850 661600 121090 661840
rect 121180 661600 121420 661840
rect 121530 661600 121770 661840
rect 110810 661270 111050 661510
rect 111140 661270 111380 661510
rect 111470 661270 111710 661510
rect 111800 661270 112040 661510
rect 112150 661270 112390 661510
rect 112480 661270 112720 661510
rect 112810 661270 113050 661510
rect 113140 661270 113380 661510
rect 113490 661270 113730 661510
rect 113820 661270 114060 661510
rect 114150 661270 114390 661510
rect 114480 661270 114720 661510
rect 114830 661270 115070 661510
rect 115160 661270 115400 661510
rect 115490 661270 115730 661510
rect 115820 661270 116060 661510
rect 116170 661270 116410 661510
rect 116500 661270 116740 661510
rect 116830 661270 117070 661510
rect 117160 661270 117400 661510
rect 117510 661270 117750 661510
rect 117840 661270 118080 661510
rect 118170 661270 118410 661510
rect 118500 661270 118740 661510
rect 118850 661270 119090 661510
rect 119180 661270 119420 661510
rect 119510 661270 119750 661510
rect 119840 661270 120080 661510
rect 120190 661270 120430 661510
rect 120520 661270 120760 661510
rect 120850 661270 121090 661510
rect 121180 661270 121420 661510
rect 121530 661270 121770 661510
rect 110810 660940 111050 661180
rect 111140 660940 111380 661180
rect 111470 660940 111710 661180
rect 111800 660940 112040 661180
rect 112150 660940 112390 661180
rect 112480 660940 112720 661180
rect 112810 660940 113050 661180
rect 113140 660940 113380 661180
rect 113490 660940 113730 661180
rect 113820 660940 114060 661180
rect 114150 660940 114390 661180
rect 114480 660940 114720 661180
rect 114830 660940 115070 661180
rect 115160 660940 115400 661180
rect 115490 660940 115730 661180
rect 115820 660940 116060 661180
rect 116170 660940 116410 661180
rect 116500 660940 116740 661180
rect 116830 660940 117070 661180
rect 117160 660940 117400 661180
rect 117510 660940 117750 661180
rect 117840 660940 118080 661180
rect 118170 660940 118410 661180
rect 118500 660940 118740 661180
rect 118850 660940 119090 661180
rect 119180 660940 119420 661180
rect 119510 660940 119750 661180
rect 119840 660940 120080 661180
rect 120190 660940 120430 661180
rect 120520 660940 120760 661180
rect 120850 660940 121090 661180
rect 121180 660940 121420 661180
rect 121530 660940 121770 661180
rect 122190 671660 122430 671900
rect 122520 671660 122760 671900
rect 122850 671660 123090 671900
rect 123180 671660 123420 671900
rect 123530 671660 123770 671900
rect 123860 671660 124100 671900
rect 124190 671660 124430 671900
rect 124520 671660 124760 671900
rect 124870 671660 125110 671900
rect 125200 671660 125440 671900
rect 125530 671660 125770 671900
rect 125860 671660 126100 671900
rect 126210 671660 126450 671900
rect 126540 671660 126780 671900
rect 126870 671660 127110 671900
rect 127200 671660 127440 671900
rect 127550 671660 127790 671900
rect 127880 671660 128120 671900
rect 128210 671660 128450 671900
rect 128540 671660 128780 671900
rect 128890 671660 129130 671900
rect 129220 671660 129460 671900
rect 129550 671660 129790 671900
rect 129880 671660 130120 671900
rect 130230 671660 130470 671900
rect 130560 671660 130800 671900
rect 130890 671660 131130 671900
rect 131220 671660 131460 671900
rect 131570 671660 131810 671900
rect 131900 671660 132140 671900
rect 132230 671660 132470 671900
rect 132560 671660 132800 671900
rect 132910 671660 133150 671900
rect 122190 671310 122430 671550
rect 122520 671310 122760 671550
rect 122850 671310 123090 671550
rect 123180 671310 123420 671550
rect 123530 671310 123770 671550
rect 123860 671310 124100 671550
rect 124190 671310 124430 671550
rect 124520 671310 124760 671550
rect 124870 671310 125110 671550
rect 125200 671310 125440 671550
rect 125530 671310 125770 671550
rect 125860 671310 126100 671550
rect 126210 671310 126450 671550
rect 126540 671310 126780 671550
rect 126870 671310 127110 671550
rect 127200 671310 127440 671550
rect 127550 671310 127790 671550
rect 127880 671310 128120 671550
rect 128210 671310 128450 671550
rect 128540 671310 128780 671550
rect 128890 671310 129130 671550
rect 129220 671310 129460 671550
rect 129550 671310 129790 671550
rect 129880 671310 130120 671550
rect 130230 671310 130470 671550
rect 130560 671310 130800 671550
rect 130890 671310 131130 671550
rect 131220 671310 131460 671550
rect 131570 671310 131810 671550
rect 131900 671310 132140 671550
rect 132230 671310 132470 671550
rect 132560 671310 132800 671550
rect 132910 671310 133150 671550
rect 122190 670980 122430 671220
rect 122520 670980 122760 671220
rect 122850 670980 123090 671220
rect 123180 670980 123420 671220
rect 123530 670980 123770 671220
rect 123860 670980 124100 671220
rect 124190 670980 124430 671220
rect 124520 670980 124760 671220
rect 124870 670980 125110 671220
rect 125200 670980 125440 671220
rect 125530 670980 125770 671220
rect 125860 670980 126100 671220
rect 126210 670980 126450 671220
rect 126540 670980 126780 671220
rect 126870 670980 127110 671220
rect 127200 670980 127440 671220
rect 127550 670980 127790 671220
rect 127880 670980 128120 671220
rect 128210 670980 128450 671220
rect 128540 670980 128780 671220
rect 128890 670980 129130 671220
rect 129220 670980 129460 671220
rect 129550 670980 129790 671220
rect 129880 670980 130120 671220
rect 130230 670980 130470 671220
rect 130560 670980 130800 671220
rect 130890 670980 131130 671220
rect 131220 670980 131460 671220
rect 131570 670980 131810 671220
rect 131900 670980 132140 671220
rect 132230 670980 132470 671220
rect 132560 670980 132800 671220
rect 132910 670980 133150 671220
rect 122190 670650 122430 670890
rect 122520 670650 122760 670890
rect 122850 670650 123090 670890
rect 123180 670650 123420 670890
rect 123530 670650 123770 670890
rect 123860 670650 124100 670890
rect 124190 670650 124430 670890
rect 124520 670650 124760 670890
rect 124870 670650 125110 670890
rect 125200 670650 125440 670890
rect 125530 670650 125770 670890
rect 125860 670650 126100 670890
rect 126210 670650 126450 670890
rect 126540 670650 126780 670890
rect 126870 670650 127110 670890
rect 127200 670650 127440 670890
rect 127550 670650 127790 670890
rect 127880 670650 128120 670890
rect 128210 670650 128450 670890
rect 128540 670650 128780 670890
rect 128890 670650 129130 670890
rect 129220 670650 129460 670890
rect 129550 670650 129790 670890
rect 129880 670650 130120 670890
rect 130230 670650 130470 670890
rect 130560 670650 130800 670890
rect 130890 670650 131130 670890
rect 131220 670650 131460 670890
rect 131570 670650 131810 670890
rect 131900 670650 132140 670890
rect 132230 670650 132470 670890
rect 132560 670650 132800 670890
rect 132910 670650 133150 670890
rect 122190 670320 122430 670560
rect 122520 670320 122760 670560
rect 122850 670320 123090 670560
rect 123180 670320 123420 670560
rect 123530 670320 123770 670560
rect 123860 670320 124100 670560
rect 124190 670320 124430 670560
rect 124520 670320 124760 670560
rect 124870 670320 125110 670560
rect 125200 670320 125440 670560
rect 125530 670320 125770 670560
rect 125860 670320 126100 670560
rect 126210 670320 126450 670560
rect 126540 670320 126780 670560
rect 126870 670320 127110 670560
rect 127200 670320 127440 670560
rect 127550 670320 127790 670560
rect 127880 670320 128120 670560
rect 128210 670320 128450 670560
rect 128540 670320 128780 670560
rect 128890 670320 129130 670560
rect 129220 670320 129460 670560
rect 129550 670320 129790 670560
rect 129880 670320 130120 670560
rect 130230 670320 130470 670560
rect 130560 670320 130800 670560
rect 130890 670320 131130 670560
rect 131220 670320 131460 670560
rect 131570 670320 131810 670560
rect 131900 670320 132140 670560
rect 132230 670320 132470 670560
rect 132560 670320 132800 670560
rect 132910 670320 133150 670560
rect 122190 669970 122430 670210
rect 122520 669970 122760 670210
rect 122850 669970 123090 670210
rect 123180 669970 123420 670210
rect 123530 669970 123770 670210
rect 123860 669970 124100 670210
rect 124190 669970 124430 670210
rect 124520 669970 124760 670210
rect 124870 669970 125110 670210
rect 125200 669970 125440 670210
rect 125530 669970 125770 670210
rect 125860 669970 126100 670210
rect 126210 669970 126450 670210
rect 126540 669970 126780 670210
rect 126870 669970 127110 670210
rect 127200 669970 127440 670210
rect 127550 669970 127790 670210
rect 127880 669970 128120 670210
rect 128210 669970 128450 670210
rect 128540 669970 128780 670210
rect 128890 669970 129130 670210
rect 129220 669970 129460 670210
rect 129550 669970 129790 670210
rect 129880 669970 130120 670210
rect 130230 669970 130470 670210
rect 130560 669970 130800 670210
rect 130890 669970 131130 670210
rect 131220 669970 131460 670210
rect 131570 669970 131810 670210
rect 131900 669970 132140 670210
rect 132230 669970 132470 670210
rect 132560 669970 132800 670210
rect 132910 669970 133150 670210
rect 122190 669640 122430 669880
rect 122520 669640 122760 669880
rect 122850 669640 123090 669880
rect 123180 669640 123420 669880
rect 123530 669640 123770 669880
rect 123860 669640 124100 669880
rect 124190 669640 124430 669880
rect 124520 669640 124760 669880
rect 124870 669640 125110 669880
rect 125200 669640 125440 669880
rect 125530 669640 125770 669880
rect 125860 669640 126100 669880
rect 126210 669640 126450 669880
rect 126540 669640 126780 669880
rect 126870 669640 127110 669880
rect 127200 669640 127440 669880
rect 127550 669640 127790 669880
rect 127880 669640 128120 669880
rect 128210 669640 128450 669880
rect 128540 669640 128780 669880
rect 128890 669640 129130 669880
rect 129220 669640 129460 669880
rect 129550 669640 129790 669880
rect 129880 669640 130120 669880
rect 130230 669640 130470 669880
rect 130560 669640 130800 669880
rect 130890 669640 131130 669880
rect 131220 669640 131460 669880
rect 131570 669640 131810 669880
rect 131900 669640 132140 669880
rect 132230 669640 132470 669880
rect 132560 669640 132800 669880
rect 132910 669640 133150 669880
rect 122190 669310 122430 669550
rect 122520 669310 122760 669550
rect 122850 669310 123090 669550
rect 123180 669310 123420 669550
rect 123530 669310 123770 669550
rect 123860 669310 124100 669550
rect 124190 669310 124430 669550
rect 124520 669310 124760 669550
rect 124870 669310 125110 669550
rect 125200 669310 125440 669550
rect 125530 669310 125770 669550
rect 125860 669310 126100 669550
rect 126210 669310 126450 669550
rect 126540 669310 126780 669550
rect 126870 669310 127110 669550
rect 127200 669310 127440 669550
rect 127550 669310 127790 669550
rect 127880 669310 128120 669550
rect 128210 669310 128450 669550
rect 128540 669310 128780 669550
rect 128890 669310 129130 669550
rect 129220 669310 129460 669550
rect 129550 669310 129790 669550
rect 129880 669310 130120 669550
rect 130230 669310 130470 669550
rect 130560 669310 130800 669550
rect 130890 669310 131130 669550
rect 131220 669310 131460 669550
rect 131570 669310 131810 669550
rect 131900 669310 132140 669550
rect 132230 669310 132470 669550
rect 132560 669310 132800 669550
rect 132910 669310 133150 669550
rect 122190 668980 122430 669220
rect 122520 668980 122760 669220
rect 122850 668980 123090 669220
rect 123180 668980 123420 669220
rect 123530 668980 123770 669220
rect 123860 668980 124100 669220
rect 124190 668980 124430 669220
rect 124520 668980 124760 669220
rect 124870 668980 125110 669220
rect 125200 668980 125440 669220
rect 125530 668980 125770 669220
rect 125860 668980 126100 669220
rect 126210 668980 126450 669220
rect 126540 668980 126780 669220
rect 126870 668980 127110 669220
rect 127200 668980 127440 669220
rect 127550 668980 127790 669220
rect 127880 668980 128120 669220
rect 128210 668980 128450 669220
rect 128540 668980 128780 669220
rect 128890 668980 129130 669220
rect 129220 668980 129460 669220
rect 129550 668980 129790 669220
rect 129880 668980 130120 669220
rect 130230 668980 130470 669220
rect 130560 668980 130800 669220
rect 130890 668980 131130 669220
rect 131220 668980 131460 669220
rect 131570 668980 131810 669220
rect 131900 668980 132140 669220
rect 132230 668980 132470 669220
rect 132560 668980 132800 669220
rect 132910 668980 133150 669220
rect 122190 668630 122430 668870
rect 122520 668630 122760 668870
rect 122850 668630 123090 668870
rect 123180 668630 123420 668870
rect 123530 668630 123770 668870
rect 123860 668630 124100 668870
rect 124190 668630 124430 668870
rect 124520 668630 124760 668870
rect 124870 668630 125110 668870
rect 125200 668630 125440 668870
rect 125530 668630 125770 668870
rect 125860 668630 126100 668870
rect 126210 668630 126450 668870
rect 126540 668630 126780 668870
rect 126870 668630 127110 668870
rect 127200 668630 127440 668870
rect 127550 668630 127790 668870
rect 127880 668630 128120 668870
rect 128210 668630 128450 668870
rect 128540 668630 128780 668870
rect 128890 668630 129130 668870
rect 129220 668630 129460 668870
rect 129550 668630 129790 668870
rect 129880 668630 130120 668870
rect 130230 668630 130470 668870
rect 130560 668630 130800 668870
rect 130890 668630 131130 668870
rect 131220 668630 131460 668870
rect 131570 668630 131810 668870
rect 131900 668630 132140 668870
rect 132230 668630 132470 668870
rect 132560 668630 132800 668870
rect 132910 668630 133150 668870
rect 122190 668300 122430 668540
rect 122520 668300 122760 668540
rect 122850 668300 123090 668540
rect 123180 668300 123420 668540
rect 123530 668300 123770 668540
rect 123860 668300 124100 668540
rect 124190 668300 124430 668540
rect 124520 668300 124760 668540
rect 124870 668300 125110 668540
rect 125200 668300 125440 668540
rect 125530 668300 125770 668540
rect 125860 668300 126100 668540
rect 126210 668300 126450 668540
rect 126540 668300 126780 668540
rect 126870 668300 127110 668540
rect 127200 668300 127440 668540
rect 127550 668300 127790 668540
rect 127880 668300 128120 668540
rect 128210 668300 128450 668540
rect 128540 668300 128780 668540
rect 128890 668300 129130 668540
rect 129220 668300 129460 668540
rect 129550 668300 129790 668540
rect 129880 668300 130120 668540
rect 130230 668300 130470 668540
rect 130560 668300 130800 668540
rect 130890 668300 131130 668540
rect 131220 668300 131460 668540
rect 131570 668300 131810 668540
rect 131900 668300 132140 668540
rect 132230 668300 132470 668540
rect 132560 668300 132800 668540
rect 132910 668300 133150 668540
rect 122190 667970 122430 668210
rect 122520 667970 122760 668210
rect 122850 667970 123090 668210
rect 123180 667970 123420 668210
rect 123530 667970 123770 668210
rect 123860 667970 124100 668210
rect 124190 667970 124430 668210
rect 124520 667970 124760 668210
rect 124870 667970 125110 668210
rect 125200 667970 125440 668210
rect 125530 667970 125770 668210
rect 125860 667970 126100 668210
rect 126210 667970 126450 668210
rect 126540 667970 126780 668210
rect 126870 667970 127110 668210
rect 127200 667970 127440 668210
rect 127550 667970 127790 668210
rect 127880 667970 128120 668210
rect 128210 667970 128450 668210
rect 128540 667970 128780 668210
rect 128890 667970 129130 668210
rect 129220 667970 129460 668210
rect 129550 667970 129790 668210
rect 129880 667970 130120 668210
rect 130230 667970 130470 668210
rect 130560 667970 130800 668210
rect 130890 667970 131130 668210
rect 131220 667970 131460 668210
rect 131570 667970 131810 668210
rect 131900 667970 132140 668210
rect 132230 667970 132470 668210
rect 132560 667970 132800 668210
rect 132910 667970 133150 668210
rect 122190 667640 122430 667880
rect 122520 667640 122760 667880
rect 122850 667640 123090 667880
rect 123180 667640 123420 667880
rect 123530 667640 123770 667880
rect 123860 667640 124100 667880
rect 124190 667640 124430 667880
rect 124520 667640 124760 667880
rect 124870 667640 125110 667880
rect 125200 667640 125440 667880
rect 125530 667640 125770 667880
rect 125860 667640 126100 667880
rect 126210 667640 126450 667880
rect 126540 667640 126780 667880
rect 126870 667640 127110 667880
rect 127200 667640 127440 667880
rect 127550 667640 127790 667880
rect 127880 667640 128120 667880
rect 128210 667640 128450 667880
rect 128540 667640 128780 667880
rect 128890 667640 129130 667880
rect 129220 667640 129460 667880
rect 129550 667640 129790 667880
rect 129880 667640 130120 667880
rect 130230 667640 130470 667880
rect 130560 667640 130800 667880
rect 130890 667640 131130 667880
rect 131220 667640 131460 667880
rect 131570 667640 131810 667880
rect 131900 667640 132140 667880
rect 132230 667640 132470 667880
rect 132560 667640 132800 667880
rect 132910 667640 133150 667880
rect 122190 667290 122430 667530
rect 122520 667290 122760 667530
rect 122850 667290 123090 667530
rect 123180 667290 123420 667530
rect 123530 667290 123770 667530
rect 123860 667290 124100 667530
rect 124190 667290 124430 667530
rect 124520 667290 124760 667530
rect 124870 667290 125110 667530
rect 125200 667290 125440 667530
rect 125530 667290 125770 667530
rect 125860 667290 126100 667530
rect 126210 667290 126450 667530
rect 126540 667290 126780 667530
rect 126870 667290 127110 667530
rect 127200 667290 127440 667530
rect 127550 667290 127790 667530
rect 127880 667290 128120 667530
rect 128210 667290 128450 667530
rect 128540 667290 128780 667530
rect 128890 667290 129130 667530
rect 129220 667290 129460 667530
rect 129550 667290 129790 667530
rect 129880 667290 130120 667530
rect 130230 667290 130470 667530
rect 130560 667290 130800 667530
rect 130890 667290 131130 667530
rect 131220 667290 131460 667530
rect 131570 667290 131810 667530
rect 131900 667290 132140 667530
rect 132230 667290 132470 667530
rect 132560 667290 132800 667530
rect 132910 667290 133150 667530
rect 122190 666960 122430 667200
rect 122520 666960 122760 667200
rect 122850 666960 123090 667200
rect 123180 666960 123420 667200
rect 123530 666960 123770 667200
rect 123860 666960 124100 667200
rect 124190 666960 124430 667200
rect 124520 666960 124760 667200
rect 124870 666960 125110 667200
rect 125200 666960 125440 667200
rect 125530 666960 125770 667200
rect 125860 666960 126100 667200
rect 126210 666960 126450 667200
rect 126540 666960 126780 667200
rect 126870 666960 127110 667200
rect 127200 666960 127440 667200
rect 127550 666960 127790 667200
rect 127880 666960 128120 667200
rect 128210 666960 128450 667200
rect 128540 666960 128780 667200
rect 128890 666960 129130 667200
rect 129220 666960 129460 667200
rect 129550 666960 129790 667200
rect 129880 666960 130120 667200
rect 130230 666960 130470 667200
rect 130560 666960 130800 667200
rect 130890 666960 131130 667200
rect 131220 666960 131460 667200
rect 131570 666960 131810 667200
rect 131900 666960 132140 667200
rect 132230 666960 132470 667200
rect 132560 666960 132800 667200
rect 132910 666960 133150 667200
rect 122190 666630 122430 666870
rect 122520 666630 122760 666870
rect 122850 666630 123090 666870
rect 123180 666630 123420 666870
rect 123530 666630 123770 666870
rect 123860 666630 124100 666870
rect 124190 666630 124430 666870
rect 124520 666630 124760 666870
rect 124870 666630 125110 666870
rect 125200 666630 125440 666870
rect 125530 666630 125770 666870
rect 125860 666630 126100 666870
rect 126210 666630 126450 666870
rect 126540 666630 126780 666870
rect 126870 666630 127110 666870
rect 127200 666630 127440 666870
rect 127550 666630 127790 666870
rect 127880 666630 128120 666870
rect 128210 666630 128450 666870
rect 128540 666630 128780 666870
rect 128890 666630 129130 666870
rect 129220 666630 129460 666870
rect 129550 666630 129790 666870
rect 129880 666630 130120 666870
rect 130230 666630 130470 666870
rect 130560 666630 130800 666870
rect 130890 666630 131130 666870
rect 131220 666630 131460 666870
rect 131570 666630 131810 666870
rect 131900 666630 132140 666870
rect 132230 666630 132470 666870
rect 132560 666630 132800 666870
rect 132910 666630 133150 666870
rect 122190 666300 122430 666540
rect 122520 666300 122760 666540
rect 122850 666300 123090 666540
rect 123180 666300 123420 666540
rect 123530 666300 123770 666540
rect 123860 666300 124100 666540
rect 124190 666300 124430 666540
rect 124520 666300 124760 666540
rect 124870 666300 125110 666540
rect 125200 666300 125440 666540
rect 125530 666300 125770 666540
rect 125860 666300 126100 666540
rect 126210 666300 126450 666540
rect 126540 666300 126780 666540
rect 126870 666300 127110 666540
rect 127200 666300 127440 666540
rect 127550 666300 127790 666540
rect 127880 666300 128120 666540
rect 128210 666300 128450 666540
rect 128540 666300 128780 666540
rect 128890 666300 129130 666540
rect 129220 666300 129460 666540
rect 129550 666300 129790 666540
rect 129880 666300 130120 666540
rect 130230 666300 130470 666540
rect 130560 666300 130800 666540
rect 130890 666300 131130 666540
rect 131220 666300 131460 666540
rect 131570 666300 131810 666540
rect 131900 666300 132140 666540
rect 132230 666300 132470 666540
rect 132560 666300 132800 666540
rect 132910 666300 133150 666540
rect 122190 665950 122430 666190
rect 122520 665950 122760 666190
rect 122850 665950 123090 666190
rect 123180 665950 123420 666190
rect 123530 665950 123770 666190
rect 123860 665950 124100 666190
rect 124190 665950 124430 666190
rect 124520 665950 124760 666190
rect 124870 665950 125110 666190
rect 125200 665950 125440 666190
rect 125530 665950 125770 666190
rect 125860 665950 126100 666190
rect 126210 665950 126450 666190
rect 126540 665950 126780 666190
rect 126870 665950 127110 666190
rect 127200 665950 127440 666190
rect 127550 665950 127790 666190
rect 127880 665950 128120 666190
rect 128210 665950 128450 666190
rect 128540 665950 128780 666190
rect 128890 665950 129130 666190
rect 129220 665950 129460 666190
rect 129550 665950 129790 666190
rect 129880 665950 130120 666190
rect 130230 665950 130470 666190
rect 130560 665950 130800 666190
rect 130890 665950 131130 666190
rect 131220 665950 131460 666190
rect 131570 665950 131810 666190
rect 131900 665950 132140 666190
rect 132230 665950 132470 666190
rect 132560 665950 132800 666190
rect 132910 665950 133150 666190
rect 122190 665620 122430 665860
rect 122520 665620 122760 665860
rect 122850 665620 123090 665860
rect 123180 665620 123420 665860
rect 123530 665620 123770 665860
rect 123860 665620 124100 665860
rect 124190 665620 124430 665860
rect 124520 665620 124760 665860
rect 124870 665620 125110 665860
rect 125200 665620 125440 665860
rect 125530 665620 125770 665860
rect 125860 665620 126100 665860
rect 126210 665620 126450 665860
rect 126540 665620 126780 665860
rect 126870 665620 127110 665860
rect 127200 665620 127440 665860
rect 127550 665620 127790 665860
rect 127880 665620 128120 665860
rect 128210 665620 128450 665860
rect 128540 665620 128780 665860
rect 128890 665620 129130 665860
rect 129220 665620 129460 665860
rect 129550 665620 129790 665860
rect 129880 665620 130120 665860
rect 130230 665620 130470 665860
rect 130560 665620 130800 665860
rect 130890 665620 131130 665860
rect 131220 665620 131460 665860
rect 131570 665620 131810 665860
rect 131900 665620 132140 665860
rect 132230 665620 132470 665860
rect 132560 665620 132800 665860
rect 132910 665620 133150 665860
rect 122190 665290 122430 665530
rect 122520 665290 122760 665530
rect 122850 665290 123090 665530
rect 123180 665290 123420 665530
rect 123530 665290 123770 665530
rect 123860 665290 124100 665530
rect 124190 665290 124430 665530
rect 124520 665290 124760 665530
rect 124870 665290 125110 665530
rect 125200 665290 125440 665530
rect 125530 665290 125770 665530
rect 125860 665290 126100 665530
rect 126210 665290 126450 665530
rect 126540 665290 126780 665530
rect 126870 665290 127110 665530
rect 127200 665290 127440 665530
rect 127550 665290 127790 665530
rect 127880 665290 128120 665530
rect 128210 665290 128450 665530
rect 128540 665290 128780 665530
rect 128890 665290 129130 665530
rect 129220 665290 129460 665530
rect 129550 665290 129790 665530
rect 129880 665290 130120 665530
rect 130230 665290 130470 665530
rect 130560 665290 130800 665530
rect 130890 665290 131130 665530
rect 131220 665290 131460 665530
rect 131570 665290 131810 665530
rect 131900 665290 132140 665530
rect 132230 665290 132470 665530
rect 132560 665290 132800 665530
rect 132910 665290 133150 665530
rect 122190 664960 122430 665200
rect 122520 664960 122760 665200
rect 122850 664960 123090 665200
rect 123180 664960 123420 665200
rect 123530 664960 123770 665200
rect 123860 664960 124100 665200
rect 124190 664960 124430 665200
rect 124520 664960 124760 665200
rect 124870 664960 125110 665200
rect 125200 664960 125440 665200
rect 125530 664960 125770 665200
rect 125860 664960 126100 665200
rect 126210 664960 126450 665200
rect 126540 664960 126780 665200
rect 126870 664960 127110 665200
rect 127200 664960 127440 665200
rect 127550 664960 127790 665200
rect 127880 664960 128120 665200
rect 128210 664960 128450 665200
rect 128540 664960 128780 665200
rect 128890 664960 129130 665200
rect 129220 664960 129460 665200
rect 129550 664960 129790 665200
rect 129880 664960 130120 665200
rect 130230 664960 130470 665200
rect 130560 664960 130800 665200
rect 130890 664960 131130 665200
rect 131220 664960 131460 665200
rect 131570 664960 131810 665200
rect 131900 664960 132140 665200
rect 132230 664960 132470 665200
rect 132560 664960 132800 665200
rect 132910 664960 133150 665200
rect 122190 664610 122430 664850
rect 122520 664610 122760 664850
rect 122850 664610 123090 664850
rect 123180 664610 123420 664850
rect 123530 664610 123770 664850
rect 123860 664610 124100 664850
rect 124190 664610 124430 664850
rect 124520 664610 124760 664850
rect 124870 664610 125110 664850
rect 125200 664610 125440 664850
rect 125530 664610 125770 664850
rect 125860 664610 126100 664850
rect 126210 664610 126450 664850
rect 126540 664610 126780 664850
rect 126870 664610 127110 664850
rect 127200 664610 127440 664850
rect 127550 664610 127790 664850
rect 127880 664610 128120 664850
rect 128210 664610 128450 664850
rect 128540 664610 128780 664850
rect 128890 664610 129130 664850
rect 129220 664610 129460 664850
rect 129550 664610 129790 664850
rect 129880 664610 130120 664850
rect 130230 664610 130470 664850
rect 130560 664610 130800 664850
rect 130890 664610 131130 664850
rect 131220 664610 131460 664850
rect 131570 664610 131810 664850
rect 131900 664610 132140 664850
rect 132230 664610 132470 664850
rect 132560 664610 132800 664850
rect 132910 664610 133150 664850
rect 122190 664280 122430 664520
rect 122520 664280 122760 664520
rect 122850 664280 123090 664520
rect 123180 664280 123420 664520
rect 123530 664280 123770 664520
rect 123860 664280 124100 664520
rect 124190 664280 124430 664520
rect 124520 664280 124760 664520
rect 124870 664280 125110 664520
rect 125200 664280 125440 664520
rect 125530 664280 125770 664520
rect 125860 664280 126100 664520
rect 126210 664280 126450 664520
rect 126540 664280 126780 664520
rect 126870 664280 127110 664520
rect 127200 664280 127440 664520
rect 127550 664280 127790 664520
rect 127880 664280 128120 664520
rect 128210 664280 128450 664520
rect 128540 664280 128780 664520
rect 128890 664280 129130 664520
rect 129220 664280 129460 664520
rect 129550 664280 129790 664520
rect 129880 664280 130120 664520
rect 130230 664280 130470 664520
rect 130560 664280 130800 664520
rect 130890 664280 131130 664520
rect 131220 664280 131460 664520
rect 131570 664280 131810 664520
rect 131900 664280 132140 664520
rect 132230 664280 132470 664520
rect 132560 664280 132800 664520
rect 132910 664280 133150 664520
rect 122190 663950 122430 664190
rect 122520 663950 122760 664190
rect 122850 663950 123090 664190
rect 123180 663950 123420 664190
rect 123530 663950 123770 664190
rect 123860 663950 124100 664190
rect 124190 663950 124430 664190
rect 124520 663950 124760 664190
rect 124870 663950 125110 664190
rect 125200 663950 125440 664190
rect 125530 663950 125770 664190
rect 125860 663950 126100 664190
rect 126210 663950 126450 664190
rect 126540 663950 126780 664190
rect 126870 663950 127110 664190
rect 127200 663950 127440 664190
rect 127550 663950 127790 664190
rect 127880 663950 128120 664190
rect 128210 663950 128450 664190
rect 128540 663950 128780 664190
rect 128890 663950 129130 664190
rect 129220 663950 129460 664190
rect 129550 663950 129790 664190
rect 129880 663950 130120 664190
rect 130230 663950 130470 664190
rect 130560 663950 130800 664190
rect 130890 663950 131130 664190
rect 131220 663950 131460 664190
rect 131570 663950 131810 664190
rect 131900 663950 132140 664190
rect 132230 663950 132470 664190
rect 132560 663950 132800 664190
rect 132910 663950 133150 664190
rect 122190 663620 122430 663860
rect 122520 663620 122760 663860
rect 122850 663620 123090 663860
rect 123180 663620 123420 663860
rect 123530 663620 123770 663860
rect 123860 663620 124100 663860
rect 124190 663620 124430 663860
rect 124520 663620 124760 663860
rect 124870 663620 125110 663860
rect 125200 663620 125440 663860
rect 125530 663620 125770 663860
rect 125860 663620 126100 663860
rect 126210 663620 126450 663860
rect 126540 663620 126780 663860
rect 126870 663620 127110 663860
rect 127200 663620 127440 663860
rect 127550 663620 127790 663860
rect 127880 663620 128120 663860
rect 128210 663620 128450 663860
rect 128540 663620 128780 663860
rect 128890 663620 129130 663860
rect 129220 663620 129460 663860
rect 129550 663620 129790 663860
rect 129880 663620 130120 663860
rect 130230 663620 130470 663860
rect 130560 663620 130800 663860
rect 130890 663620 131130 663860
rect 131220 663620 131460 663860
rect 131570 663620 131810 663860
rect 131900 663620 132140 663860
rect 132230 663620 132470 663860
rect 132560 663620 132800 663860
rect 132910 663620 133150 663860
rect 122190 663270 122430 663510
rect 122520 663270 122760 663510
rect 122850 663270 123090 663510
rect 123180 663270 123420 663510
rect 123530 663270 123770 663510
rect 123860 663270 124100 663510
rect 124190 663270 124430 663510
rect 124520 663270 124760 663510
rect 124870 663270 125110 663510
rect 125200 663270 125440 663510
rect 125530 663270 125770 663510
rect 125860 663270 126100 663510
rect 126210 663270 126450 663510
rect 126540 663270 126780 663510
rect 126870 663270 127110 663510
rect 127200 663270 127440 663510
rect 127550 663270 127790 663510
rect 127880 663270 128120 663510
rect 128210 663270 128450 663510
rect 128540 663270 128780 663510
rect 128890 663270 129130 663510
rect 129220 663270 129460 663510
rect 129550 663270 129790 663510
rect 129880 663270 130120 663510
rect 130230 663270 130470 663510
rect 130560 663270 130800 663510
rect 130890 663270 131130 663510
rect 131220 663270 131460 663510
rect 131570 663270 131810 663510
rect 131900 663270 132140 663510
rect 132230 663270 132470 663510
rect 132560 663270 132800 663510
rect 132910 663270 133150 663510
rect 122190 662940 122430 663180
rect 122520 662940 122760 663180
rect 122850 662940 123090 663180
rect 123180 662940 123420 663180
rect 123530 662940 123770 663180
rect 123860 662940 124100 663180
rect 124190 662940 124430 663180
rect 124520 662940 124760 663180
rect 124870 662940 125110 663180
rect 125200 662940 125440 663180
rect 125530 662940 125770 663180
rect 125860 662940 126100 663180
rect 126210 662940 126450 663180
rect 126540 662940 126780 663180
rect 126870 662940 127110 663180
rect 127200 662940 127440 663180
rect 127550 662940 127790 663180
rect 127880 662940 128120 663180
rect 128210 662940 128450 663180
rect 128540 662940 128780 663180
rect 128890 662940 129130 663180
rect 129220 662940 129460 663180
rect 129550 662940 129790 663180
rect 129880 662940 130120 663180
rect 130230 662940 130470 663180
rect 130560 662940 130800 663180
rect 130890 662940 131130 663180
rect 131220 662940 131460 663180
rect 131570 662940 131810 663180
rect 131900 662940 132140 663180
rect 132230 662940 132470 663180
rect 132560 662940 132800 663180
rect 132910 662940 133150 663180
rect 122190 662610 122430 662850
rect 122520 662610 122760 662850
rect 122850 662610 123090 662850
rect 123180 662610 123420 662850
rect 123530 662610 123770 662850
rect 123860 662610 124100 662850
rect 124190 662610 124430 662850
rect 124520 662610 124760 662850
rect 124870 662610 125110 662850
rect 125200 662610 125440 662850
rect 125530 662610 125770 662850
rect 125860 662610 126100 662850
rect 126210 662610 126450 662850
rect 126540 662610 126780 662850
rect 126870 662610 127110 662850
rect 127200 662610 127440 662850
rect 127550 662610 127790 662850
rect 127880 662610 128120 662850
rect 128210 662610 128450 662850
rect 128540 662610 128780 662850
rect 128890 662610 129130 662850
rect 129220 662610 129460 662850
rect 129550 662610 129790 662850
rect 129880 662610 130120 662850
rect 130230 662610 130470 662850
rect 130560 662610 130800 662850
rect 130890 662610 131130 662850
rect 131220 662610 131460 662850
rect 131570 662610 131810 662850
rect 131900 662610 132140 662850
rect 132230 662610 132470 662850
rect 132560 662610 132800 662850
rect 132910 662610 133150 662850
rect 122190 662280 122430 662520
rect 122520 662280 122760 662520
rect 122850 662280 123090 662520
rect 123180 662280 123420 662520
rect 123530 662280 123770 662520
rect 123860 662280 124100 662520
rect 124190 662280 124430 662520
rect 124520 662280 124760 662520
rect 124870 662280 125110 662520
rect 125200 662280 125440 662520
rect 125530 662280 125770 662520
rect 125860 662280 126100 662520
rect 126210 662280 126450 662520
rect 126540 662280 126780 662520
rect 126870 662280 127110 662520
rect 127200 662280 127440 662520
rect 127550 662280 127790 662520
rect 127880 662280 128120 662520
rect 128210 662280 128450 662520
rect 128540 662280 128780 662520
rect 128890 662280 129130 662520
rect 129220 662280 129460 662520
rect 129550 662280 129790 662520
rect 129880 662280 130120 662520
rect 130230 662280 130470 662520
rect 130560 662280 130800 662520
rect 130890 662280 131130 662520
rect 131220 662280 131460 662520
rect 131570 662280 131810 662520
rect 131900 662280 132140 662520
rect 132230 662280 132470 662520
rect 132560 662280 132800 662520
rect 132910 662280 133150 662520
rect 122190 661930 122430 662170
rect 122520 661930 122760 662170
rect 122850 661930 123090 662170
rect 123180 661930 123420 662170
rect 123530 661930 123770 662170
rect 123860 661930 124100 662170
rect 124190 661930 124430 662170
rect 124520 661930 124760 662170
rect 124870 661930 125110 662170
rect 125200 661930 125440 662170
rect 125530 661930 125770 662170
rect 125860 661930 126100 662170
rect 126210 661930 126450 662170
rect 126540 661930 126780 662170
rect 126870 661930 127110 662170
rect 127200 661930 127440 662170
rect 127550 661930 127790 662170
rect 127880 661930 128120 662170
rect 128210 661930 128450 662170
rect 128540 661930 128780 662170
rect 128890 661930 129130 662170
rect 129220 661930 129460 662170
rect 129550 661930 129790 662170
rect 129880 661930 130120 662170
rect 130230 661930 130470 662170
rect 130560 661930 130800 662170
rect 130890 661930 131130 662170
rect 131220 661930 131460 662170
rect 131570 661930 131810 662170
rect 131900 661930 132140 662170
rect 132230 661930 132470 662170
rect 132560 661930 132800 662170
rect 132910 661930 133150 662170
rect 122190 661600 122430 661840
rect 122520 661600 122760 661840
rect 122850 661600 123090 661840
rect 123180 661600 123420 661840
rect 123530 661600 123770 661840
rect 123860 661600 124100 661840
rect 124190 661600 124430 661840
rect 124520 661600 124760 661840
rect 124870 661600 125110 661840
rect 125200 661600 125440 661840
rect 125530 661600 125770 661840
rect 125860 661600 126100 661840
rect 126210 661600 126450 661840
rect 126540 661600 126780 661840
rect 126870 661600 127110 661840
rect 127200 661600 127440 661840
rect 127550 661600 127790 661840
rect 127880 661600 128120 661840
rect 128210 661600 128450 661840
rect 128540 661600 128780 661840
rect 128890 661600 129130 661840
rect 129220 661600 129460 661840
rect 129550 661600 129790 661840
rect 129880 661600 130120 661840
rect 130230 661600 130470 661840
rect 130560 661600 130800 661840
rect 130890 661600 131130 661840
rect 131220 661600 131460 661840
rect 131570 661600 131810 661840
rect 131900 661600 132140 661840
rect 132230 661600 132470 661840
rect 132560 661600 132800 661840
rect 132910 661600 133150 661840
rect 122190 661270 122430 661510
rect 122520 661270 122760 661510
rect 122850 661270 123090 661510
rect 123180 661270 123420 661510
rect 123530 661270 123770 661510
rect 123860 661270 124100 661510
rect 124190 661270 124430 661510
rect 124520 661270 124760 661510
rect 124870 661270 125110 661510
rect 125200 661270 125440 661510
rect 125530 661270 125770 661510
rect 125860 661270 126100 661510
rect 126210 661270 126450 661510
rect 126540 661270 126780 661510
rect 126870 661270 127110 661510
rect 127200 661270 127440 661510
rect 127550 661270 127790 661510
rect 127880 661270 128120 661510
rect 128210 661270 128450 661510
rect 128540 661270 128780 661510
rect 128890 661270 129130 661510
rect 129220 661270 129460 661510
rect 129550 661270 129790 661510
rect 129880 661270 130120 661510
rect 130230 661270 130470 661510
rect 130560 661270 130800 661510
rect 130890 661270 131130 661510
rect 131220 661270 131460 661510
rect 131570 661270 131810 661510
rect 131900 661270 132140 661510
rect 132230 661270 132470 661510
rect 132560 661270 132800 661510
rect 132910 661270 133150 661510
rect 122190 660940 122430 661180
rect 122520 660940 122760 661180
rect 122850 660940 123090 661180
rect 123180 660940 123420 661180
rect 123530 660940 123770 661180
rect 123860 660940 124100 661180
rect 124190 660940 124430 661180
rect 124520 660940 124760 661180
rect 124870 660940 125110 661180
rect 125200 660940 125440 661180
rect 125530 660940 125770 661180
rect 125860 660940 126100 661180
rect 126210 660940 126450 661180
rect 126540 660940 126780 661180
rect 126870 660940 127110 661180
rect 127200 660940 127440 661180
rect 127550 660940 127790 661180
rect 127880 660940 128120 661180
rect 128210 660940 128450 661180
rect 128540 660940 128780 661180
rect 128890 660940 129130 661180
rect 129220 660940 129460 661180
rect 129550 660940 129790 661180
rect 129880 660940 130120 661180
rect 130230 660940 130470 661180
rect 130560 660940 130800 661180
rect 130890 660940 131130 661180
rect 131220 660940 131460 661180
rect 131570 660940 131810 661180
rect 131900 660940 132140 661180
rect 132230 660940 132470 661180
rect 132560 660940 132800 661180
rect 132910 660940 133150 661180
rect 133570 671660 133810 671900
rect 133900 671660 134140 671900
rect 134230 671660 134470 671900
rect 134560 671660 134800 671900
rect 134910 671660 135150 671900
rect 135240 671660 135480 671900
rect 135570 671660 135810 671900
rect 135900 671660 136140 671900
rect 136250 671660 136490 671900
rect 136580 671660 136820 671900
rect 136910 671660 137150 671900
rect 137240 671660 137480 671900
rect 137590 671660 137830 671900
rect 137920 671660 138160 671900
rect 138250 671660 138490 671900
rect 138580 671660 138820 671900
rect 138930 671660 139170 671900
rect 139260 671660 139500 671900
rect 139590 671660 139830 671900
rect 139920 671660 140160 671900
rect 140270 671660 140510 671900
rect 140600 671660 140840 671900
rect 140930 671660 141170 671900
rect 141260 671660 141500 671900
rect 141610 671660 141850 671900
rect 141940 671660 142180 671900
rect 142270 671660 142510 671900
rect 142600 671660 142840 671900
rect 142950 671660 143190 671900
rect 143280 671660 143520 671900
rect 143610 671660 143850 671900
rect 143940 671660 144180 671900
rect 144290 671660 144530 671900
rect 133570 671310 133810 671550
rect 133900 671310 134140 671550
rect 134230 671310 134470 671550
rect 134560 671310 134800 671550
rect 134910 671310 135150 671550
rect 135240 671310 135480 671550
rect 135570 671310 135810 671550
rect 135900 671310 136140 671550
rect 136250 671310 136490 671550
rect 136580 671310 136820 671550
rect 136910 671310 137150 671550
rect 137240 671310 137480 671550
rect 137590 671310 137830 671550
rect 137920 671310 138160 671550
rect 138250 671310 138490 671550
rect 138580 671310 138820 671550
rect 138930 671310 139170 671550
rect 139260 671310 139500 671550
rect 139590 671310 139830 671550
rect 139920 671310 140160 671550
rect 140270 671310 140510 671550
rect 140600 671310 140840 671550
rect 140930 671310 141170 671550
rect 141260 671310 141500 671550
rect 141610 671310 141850 671550
rect 141940 671310 142180 671550
rect 142270 671310 142510 671550
rect 142600 671310 142840 671550
rect 142950 671310 143190 671550
rect 143280 671310 143520 671550
rect 143610 671310 143850 671550
rect 143940 671310 144180 671550
rect 144290 671310 144530 671550
rect 133570 670980 133810 671220
rect 133900 670980 134140 671220
rect 134230 670980 134470 671220
rect 134560 670980 134800 671220
rect 134910 670980 135150 671220
rect 135240 670980 135480 671220
rect 135570 670980 135810 671220
rect 135900 670980 136140 671220
rect 136250 670980 136490 671220
rect 136580 670980 136820 671220
rect 136910 670980 137150 671220
rect 137240 670980 137480 671220
rect 137590 670980 137830 671220
rect 137920 670980 138160 671220
rect 138250 670980 138490 671220
rect 138580 670980 138820 671220
rect 138930 670980 139170 671220
rect 139260 670980 139500 671220
rect 139590 670980 139830 671220
rect 139920 670980 140160 671220
rect 140270 670980 140510 671220
rect 140600 670980 140840 671220
rect 140930 670980 141170 671220
rect 141260 670980 141500 671220
rect 141610 670980 141850 671220
rect 141940 670980 142180 671220
rect 142270 670980 142510 671220
rect 142600 670980 142840 671220
rect 142950 670980 143190 671220
rect 143280 670980 143520 671220
rect 143610 670980 143850 671220
rect 143940 670980 144180 671220
rect 144290 670980 144530 671220
rect 133570 670650 133810 670890
rect 133900 670650 134140 670890
rect 134230 670650 134470 670890
rect 134560 670650 134800 670890
rect 134910 670650 135150 670890
rect 135240 670650 135480 670890
rect 135570 670650 135810 670890
rect 135900 670650 136140 670890
rect 136250 670650 136490 670890
rect 136580 670650 136820 670890
rect 136910 670650 137150 670890
rect 137240 670650 137480 670890
rect 137590 670650 137830 670890
rect 137920 670650 138160 670890
rect 138250 670650 138490 670890
rect 138580 670650 138820 670890
rect 138930 670650 139170 670890
rect 139260 670650 139500 670890
rect 139590 670650 139830 670890
rect 139920 670650 140160 670890
rect 140270 670650 140510 670890
rect 140600 670650 140840 670890
rect 140930 670650 141170 670890
rect 141260 670650 141500 670890
rect 141610 670650 141850 670890
rect 141940 670650 142180 670890
rect 142270 670650 142510 670890
rect 142600 670650 142840 670890
rect 142950 670650 143190 670890
rect 143280 670650 143520 670890
rect 143610 670650 143850 670890
rect 143940 670650 144180 670890
rect 144290 670650 144530 670890
rect 133570 670320 133810 670560
rect 133900 670320 134140 670560
rect 134230 670320 134470 670560
rect 134560 670320 134800 670560
rect 134910 670320 135150 670560
rect 135240 670320 135480 670560
rect 135570 670320 135810 670560
rect 135900 670320 136140 670560
rect 136250 670320 136490 670560
rect 136580 670320 136820 670560
rect 136910 670320 137150 670560
rect 137240 670320 137480 670560
rect 137590 670320 137830 670560
rect 137920 670320 138160 670560
rect 138250 670320 138490 670560
rect 138580 670320 138820 670560
rect 138930 670320 139170 670560
rect 139260 670320 139500 670560
rect 139590 670320 139830 670560
rect 139920 670320 140160 670560
rect 140270 670320 140510 670560
rect 140600 670320 140840 670560
rect 140930 670320 141170 670560
rect 141260 670320 141500 670560
rect 141610 670320 141850 670560
rect 141940 670320 142180 670560
rect 142270 670320 142510 670560
rect 142600 670320 142840 670560
rect 142950 670320 143190 670560
rect 143280 670320 143520 670560
rect 143610 670320 143850 670560
rect 143940 670320 144180 670560
rect 144290 670320 144530 670560
rect 133570 669970 133810 670210
rect 133900 669970 134140 670210
rect 134230 669970 134470 670210
rect 134560 669970 134800 670210
rect 134910 669970 135150 670210
rect 135240 669970 135480 670210
rect 135570 669970 135810 670210
rect 135900 669970 136140 670210
rect 136250 669970 136490 670210
rect 136580 669970 136820 670210
rect 136910 669970 137150 670210
rect 137240 669970 137480 670210
rect 137590 669970 137830 670210
rect 137920 669970 138160 670210
rect 138250 669970 138490 670210
rect 138580 669970 138820 670210
rect 138930 669970 139170 670210
rect 139260 669970 139500 670210
rect 139590 669970 139830 670210
rect 139920 669970 140160 670210
rect 140270 669970 140510 670210
rect 140600 669970 140840 670210
rect 140930 669970 141170 670210
rect 141260 669970 141500 670210
rect 141610 669970 141850 670210
rect 141940 669970 142180 670210
rect 142270 669970 142510 670210
rect 142600 669970 142840 670210
rect 142950 669970 143190 670210
rect 143280 669970 143520 670210
rect 143610 669970 143850 670210
rect 143940 669970 144180 670210
rect 144290 669970 144530 670210
rect 133570 669640 133810 669880
rect 133900 669640 134140 669880
rect 134230 669640 134470 669880
rect 134560 669640 134800 669880
rect 134910 669640 135150 669880
rect 135240 669640 135480 669880
rect 135570 669640 135810 669880
rect 135900 669640 136140 669880
rect 136250 669640 136490 669880
rect 136580 669640 136820 669880
rect 136910 669640 137150 669880
rect 137240 669640 137480 669880
rect 137590 669640 137830 669880
rect 137920 669640 138160 669880
rect 138250 669640 138490 669880
rect 138580 669640 138820 669880
rect 138930 669640 139170 669880
rect 139260 669640 139500 669880
rect 139590 669640 139830 669880
rect 139920 669640 140160 669880
rect 140270 669640 140510 669880
rect 140600 669640 140840 669880
rect 140930 669640 141170 669880
rect 141260 669640 141500 669880
rect 141610 669640 141850 669880
rect 141940 669640 142180 669880
rect 142270 669640 142510 669880
rect 142600 669640 142840 669880
rect 142950 669640 143190 669880
rect 143280 669640 143520 669880
rect 143610 669640 143850 669880
rect 143940 669640 144180 669880
rect 144290 669640 144530 669880
rect 133570 669310 133810 669550
rect 133900 669310 134140 669550
rect 134230 669310 134470 669550
rect 134560 669310 134800 669550
rect 134910 669310 135150 669550
rect 135240 669310 135480 669550
rect 135570 669310 135810 669550
rect 135900 669310 136140 669550
rect 136250 669310 136490 669550
rect 136580 669310 136820 669550
rect 136910 669310 137150 669550
rect 137240 669310 137480 669550
rect 137590 669310 137830 669550
rect 137920 669310 138160 669550
rect 138250 669310 138490 669550
rect 138580 669310 138820 669550
rect 138930 669310 139170 669550
rect 139260 669310 139500 669550
rect 139590 669310 139830 669550
rect 139920 669310 140160 669550
rect 140270 669310 140510 669550
rect 140600 669310 140840 669550
rect 140930 669310 141170 669550
rect 141260 669310 141500 669550
rect 141610 669310 141850 669550
rect 141940 669310 142180 669550
rect 142270 669310 142510 669550
rect 142600 669310 142840 669550
rect 142950 669310 143190 669550
rect 143280 669310 143520 669550
rect 143610 669310 143850 669550
rect 143940 669310 144180 669550
rect 144290 669310 144530 669550
rect 133570 668980 133810 669220
rect 133900 668980 134140 669220
rect 134230 668980 134470 669220
rect 134560 668980 134800 669220
rect 134910 668980 135150 669220
rect 135240 668980 135480 669220
rect 135570 668980 135810 669220
rect 135900 668980 136140 669220
rect 136250 668980 136490 669220
rect 136580 668980 136820 669220
rect 136910 668980 137150 669220
rect 137240 668980 137480 669220
rect 137590 668980 137830 669220
rect 137920 668980 138160 669220
rect 138250 668980 138490 669220
rect 138580 668980 138820 669220
rect 138930 668980 139170 669220
rect 139260 668980 139500 669220
rect 139590 668980 139830 669220
rect 139920 668980 140160 669220
rect 140270 668980 140510 669220
rect 140600 668980 140840 669220
rect 140930 668980 141170 669220
rect 141260 668980 141500 669220
rect 141610 668980 141850 669220
rect 141940 668980 142180 669220
rect 142270 668980 142510 669220
rect 142600 668980 142840 669220
rect 142950 668980 143190 669220
rect 143280 668980 143520 669220
rect 143610 668980 143850 669220
rect 143940 668980 144180 669220
rect 144290 668980 144530 669220
rect 133570 668630 133810 668870
rect 133900 668630 134140 668870
rect 134230 668630 134470 668870
rect 134560 668630 134800 668870
rect 134910 668630 135150 668870
rect 135240 668630 135480 668870
rect 135570 668630 135810 668870
rect 135900 668630 136140 668870
rect 136250 668630 136490 668870
rect 136580 668630 136820 668870
rect 136910 668630 137150 668870
rect 137240 668630 137480 668870
rect 137590 668630 137830 668870
rect 137920 668630 138160 668870
rect 138250 668630 138490 668870
rect 138580 668630 138820 668870
rect 138930 668630 139170 668870
rect 139260 668630 139500 668870
rect 139590 668630 139830 668870
rect 139920 668630 140160 668870
rect 140270 668630 140510 668870
rect 140600 668630 140840 668870
rect 140930 668630 141170 668870
rect 141260 668630 141500 668870
rect 141610 668630 141850 668870
rect 141940 668630 142180 668870
rect 142270 668630 142510 668870
rect 142600 668630 142840 668870
rect 142950 668630 143190 668870
rect 143280 668630 143520 668870
rect 143610 668630 143850 668870
rect 143940 668630 144180 668870
rect 144290 668630 144530 668870
rect 133570 668300 133810 668540
rect 133900 668300 134140 668540
rect 134230 668300 134470 668540
rect 134560 668300 134800 668540
rect 134910 668300 135150 668540
rect 135240 668300 135480 668540
rect 135570 668300 135810 668540
rect 135900 668300 136140 668540
rect 136250 668300 136490 668540
rect 136580 668300 136820 668540
rect 136910 668300 137150 668540
rect 137240 668300 137480 668540
rect 137590 668300 137830 668540
rect 137920 668300 138160 668540
rect 138250 668300 138490 668540
rect 138580 668300 138820 668540
rect 138930 668300 139170 668540
rect 139260 668300 139500 668540
rect 139590 668300 139830 668540
rect 139920 668300 140160 668540
rect 140270 668300 140510 668540
rect 140600 668300 140840 668540
rect 140930 668300 141170 668540
rect 141260 668300 141500 668540
rect 141610 668300 141850 668540
rect 141940 668300 142180 668540
rect 142270 668300 142510 668540
rect 142600 668300 142840 668540
rect 142950 668300 143190 668540
rect 143280 668300 143520 668540
rect 143610 668300 143850 668540
rect 143940 668300 144180 668540
rect 144290 668300 144530 668540
rect 133570 667970 133810 668210
rect 133900 667970 134140 668210
rect 134230 667970 134470 668210
rect 134560 667970 134800 668210
rect 134910 667970 135150 668210
rect 135240 667970 135480 668210
rect 135570 667970 135810 668210
rect 135900 667970 136140 668210
rect 136250 667970 136490 668210
rect 136580 667970 136820 668210
rect 136910 667970 137150 668210
rect 137240 667970 137480 668210
rect 137590 667970 137830 668210
rect 137920 667970 138160 668210
rect 138250 667970 138490 668210
rect 138580 667970 138820 668210
rect 138930 667970 139170 668210
rect 139260 667970 139500 668210
rect 139590 667970 139830 668210
rect 139920 667970 140160 668210
rect 140270 667970 140510 668210
rect 140600 667970 140840 668210
rect 140930 667970 141170 668210
rect 141260 667970 141500 668210
rect 141610 667970 141850 668210
rect 141940 667970 142180 668210
rect 142270 667970 142510 668210
rect 142600 667970 142840 668210
rect 142950 667970 143190 668210
rect 143280 667970 143520 668210
rect 143610 667970 143850 668210
rect 143940 667970 144180 668210
rect 144290 667970 144530 668210
rect 133570 667640 133810 667880
rect 133900 667640 134140 667880
rect 134230 667640 134470 667880
rect 134560 667640 134800 667880
rect 134910 667640 135150 667880
rect 135240 667640 135480 667880
rect 135570 667640 135810 667880
rect 135900 667640 136140 667880
rect 136250 667640 136490 667880
rect 136580 667640 136820 667880
rect 136910 667640 137150 667880
rect 137240 667640 137480 667880
rect 137590 667640 137830 667880
rect 137920 667640 138160 667880
rect 138250 667640 138490 667880
rect 138580 667640 138820 667880
rect 138930 667640 139170 667880
rect 139260 667640 139500 667880
rect 139590 667640 139830 667880
rect 139920 667640 140160 667880
rect 140270 667640 140510 667880
rect 140600 667640 140840 667880
rect 140930 667640 141170 667880
rect 141260 667640 141500 667880
rect 141610 667640 141850 667880
rect 141940 667640 142180 667880
rect 142270 667640 142510 667880
rect 142600 667640 142840 667880
rect 142950 667640 143190 667880
rect 143280 667640 143520 667880
rect 143610 667640 143850 667880
rect 143940 667640 144180 667880
rect 144290 667640 144530 667880
rect 133570 667290 133810 667530
rect 133900 667290 134140 667530
rect 134230 667290 134470 667530
rect 134560 667290 134800 667530
rect 134910 667290 135150 667530
rect 135240 667290 135480 667530
rect 135570 667290 135810 667530
rect 135900 667290 136140 667530
rect 136250 667290 136490 667530
rect 136580 667290 136820 667530
rect 136910 667290 137150 667530
rect 137240 667290 137480 667530
rect 137590 667290 137830 667530
rect 137920 667290 138160 667530
rect 138250 667290 138490 667530
rect 138580 667290 138820 667530
rect 138930 667290 139170 667530
rect 139260 667290 139500 667530
rect 139590 667290 139830 667530
rect 139920 667290 140160 667530
rect 140270 667290 140510 667530
rect 140600 667290 140840 667530
rect 140930 667290 141170 667530
rect 141260 667290 141500 667530
rect 141610 667290 141850 667530
rect 141940 667290 142180 667530
rect 142270 667290 142510 667530
rect 142600 667290 142840 667530
rect 142950 667290 143190 667530
rect 143280 667290 143520 667530
rect 143610 667290 143850 667530
rect 143940 667290 144180 667530
rect 144290 667290 144530 667530
rect 133570 666960 133810 667200
rect 133900 666960 134140 667200
rect 134230 666960 134470 667200
rect 134560 666960 134800 667200
rect 134910 666960 135150 667200
rect 135240 666960 135480 667200
rect 135570 666960 135810 667200
rect 135900 666960 136140 667200
rect 136250 666960 136490 667200
rect 136580 666960 136820 667200
rect 136910 666960 137150 667200
rect 137240 666960 137480 667200
rect 137590 666960 137830 667200
rect 137920 666960 138160 667200
rect 138250 666960 138490 667200
rect 138580 666960 138820 667200
rect 138930 666960 139170 667200
rect 139260 666960 139500 667200
rect 139590 666960 139830 667200
rect 139920 666960 140160 667200
rect 140270 666960 140510 667200
rect 140600 666960 140840 667200
rect 140930 666960 141170 667200
rect 141260 666960 141500 667200
rect 141610 666960 141850 667200
rect 141940 666960 142180 667200
rect 142270 666960 142510 667200
rect 142600 666960 142840 667200
rect 142950 666960 143190 667200
rect 143280 666960 143520 667200
rect 143610 666960 143850 667200
rect 143940 666960 144180 667200
rect 144290 666960 144530 667200
rect 133570 666630 133810 666870
rect 133900 666630 134140 666870
rect 134230 666630 134470 666870
rect 134560 666630 134800 666870
rect 134910 666630 135150 666870
rect 135240 666630 135480 666870
rect 135570 666630 135810 666870
rect 135900 666630 136140 666870
rect 136250 666630 136490 666870
rect 136580 666630 136820 666870
rect 136910 666630 137150 666870
rect 137240 666630 137480 666870
rect 137590 666630 137830 666870
rect 137920 666630 138160 666870
rect 138250 666630 138490 666870
rect 138580 666630 138820 666870
rect 138930 666630 139170 666870
rect 139260 666630 139500 666870
rect 139590 666630 139830 666870
rect 139920 666630 140160 666870
rect 140270 666630 140510 666870
rect 140600 666630 140840 666870
rect 140930 666630 141170 666870
rect 141260 666630 141500 666870
rect 141610 666630 141850 666870
rect 141940 666630 142180 666870
rect 142270 666630 142510 666870
rect 142600 666630 142840 666870
rect 142950 666630 143190 666870
rect 143280 666630 143520 666870
rect 143610 666630 143850 666870
rect 143940 666630 144180 666870
rect 144290 666630 144530 666870
rect 133570 666300 133810 666540
rect 133900 666300 134140 666540
rect 134230 666300 134470 666540
rect 134560 666300 134800 666540
rect 134910 666300 135150 666540
rect 135240 666300 135480 666540
rect 135570 666300 135810 666540
rect 135900 666300 136140 666540
rect 136250 666300 136490 666540
rect 136580 666300 136820 666540
rect 136910 666300 137150 666540
rect 137240 666300 137480 666540
rect 137590 666300 137830 666540
rect 137920 666300 138160 666540
rect 138250 666300 138490 666540
rect 138580 666300 138820 666540
rect 138930 666300 139170 666540
rect 139260 666300 139500 666540
rect 139590 666300 139830 666540
rect 139920 666300 140160 666540
rect 140270 666300 140510 666540
rect 140600 666300 140840 666540
rect 140930 666300 141170 666540
rect 141260 666300 141500 666540
rect 141610 666300 141850 666540
rect 141940 666300 142180 666540
rect 142270 666300 142510 666540
rect 142600 666300 142840 666540
rect 142950 666300 143190 666540
rect 143280 666300 143520 666540
rect 143610 666300 143850 666540
rect 143940 666300 144180 666540
rect 144290 666300 144530 666540
rect 133570 665950 133810 666190
rect 133900 665950 134140 666190
rect 134230 665950 134470 666190
rect 134560 665950 134800 666190
rect 134910 665950 135150 666190
rect 135240 665950 135480 666190
rect 135570 665950 135810 666190
rect 135900 665950 136140 666190
rect 136250 665950 136490 666190
rect 136580 665950 136820 666190
rect 136910 665950 137150 666190
rect 137240 665950 137480 666190
rect 137590 665950 137830 666190
rect 137920 665950 138160 666190
rect 138250 665950 138490 666190
rect 138580 665950 138820 666190
rect 138930 665950 139170 666190
rect 139260 665950 139500 666190
rect 139590 665950 139830 666190
rect 139920 665950 140160 666190
rect 140270 665950 140510 666190
rect 140600 665950 140840 666190
rect 140930 665950 141170 666190
rect 141260 665950 141500 666190
rect 141610 665950 141850 666190
rect 141940 665950 142180 666190
rect 142270 665950 142510 666190
rect 142600 665950 142840 666190
rect 142950 665950 143190 666190
rect 143280 665950 143520 666190
rect 143610 665950 143850 666190
rect 143940 665950 144180 666190
rect 144290 665950 144530 666190
rect 133570 665620 133810 665860
rect 133900 665620 134140 665860
rect 134230 665620 134470 665860
rect 134560 665620 134800 665860
rect 134910 665620 135150 665860
rect 135240 665620 135480 665860
rect 135570 665620 135810 665860
rect 135900 665620 136140 665860
rect 136250 665620 136490 665860
rect 136580 665620 136820 665860
rect 136910 665620 137150 665860
rect 137240 665620 137480 665860
rect 137590 665620 137830 665860
rect 137920 665620 138160 665860
rect 138250 665620 138490 665860
rect 138580 665620 138820 665860
rect 138930 665620 139170 665860
rect 139260 665620 139500 665860
rect 139590 665620 139830 665860
rect 139920 665620 140160 665860
rect 140270 665620 140510 665860
rect 140600 665620 140840 665860
rect 140930 665620 141170 665860
rect 141260 665620 141500 665860
rect 141610 665620 141850 665860
rect 141940 665620 142180 665860
rect 142270 665620 142510 665860
rect 142600 665620 142840 665860
rect 142950 665620 143190 665860
rect 143280 665620 143520 665860
rect 143610 665620 143850 665860
rect 143940 665620 144180 665860
rect 144290 665620 144530 665860
rect 133570 665290 133810 665530
rect 133900 665290 134140 665530
rect 134230 665290 134470 665530
rect 134560 665290 134800 665530
rect 134910 665290 135150 665530
rect 135240 665290 135480 665530
rect 135570 665290 135810 665530
rect 135900 665290 136140 665530
rect 136250 665290 136490 665530
rect 136580 665290 136820 665530
rect 136910 665290 137150 665530
rect 137240 665290 137480 665530
rect 137590 665290 137830 665530
rect 137920 665290 138160 665530
rect 138250 665290 138490 665530
rect 138580 665290 138820 665530
rect 138930 665290 139170 665530
rect 139260 665290 139500 665530
rect 139590 665290 139830 665530
rect 139920 665290 140160 665530
rect 140270 665290 140510 665530
rect 140600 665290 140840 665530
rect 140930 665290 141170 665530
rect 141260 665290 141500 665530
rect 141610 665290 141850 665530
rect 141940 665290 142180 665530
rect 142270 665290 142510 665530
rect 142600 665290 142840 665530
rect 142950 665290 143190 665530
rect 143280 665290 143520 665530
rect 143610 665290 143850 665530
rect 143940 665290 144180 665530
rect 144290 665290 144530 665530
rect 133570 664960 133810 665200
rect 133900 664960 134140 665200
rect 134230 664960 134470 665200
rect 134560 664960 134800 665200
rect 134910 664960 135150 665200
rect 135240 664960 135480 665200
rect 135570 664960 135810 665200
rect 135900 664960 136140 665200
rect 136250 664960 136490 665200
rect 136580 664960 136820 665200
rect 136910 664960 137150 665200
rect 137240 664960 137480 665200
rect 137590 664960 137830 665200
rect 137920 664960 138160 665200
rect 138250 664960 138490 665200
rect 138580 664960 138820 665200
rect 138930 664960 139170 665200
rect 139260 664960 139500 665200
rect 139590 664960 139830 665200
rect 139920 664960 140160 665200
rect 140270 664960 140510 665200
rect 140600 664960 140840 665200
rect 140930 664960 141170 665200
rect 141260 664960 141500 665200
rect 141610 664960 141850 665200
rect 141940 664960 142180 665200
rect 142270 664960 142510 665200
rect 142600 664960 142840 665200
rect 142950 664960 143190 665200
rect 143280 664960 143520 665200
rect 143610 664960 143850 665200
rect 143940 664960 144180 665200
rect 144290 664960 144530 665200
rect 133570 664610 133810 664850
rect 133900 664610 134140 664850
rect 134230 664610 134470 664850
rect 134560 664610 134800 664850
rect 134910 664610 135150 664850
rect 135240 664610 135480 664850
rect 135570 664610 135810 664850
rect 135900 664610 136140 664850
rect 136250 664610 136490 664850
rect 136580 664610 136820 664850
rect 136910 664610 137150 664850
rect 137240 664610 137480 664850
rect 137590 664610 137830 664850
rect 137920 664610 138160 664850
rect 138250 664610 138490 664850
rect 138580 664610 138820 664850
rect 138930 664610 139170 664850
rect 139260 664610 139500 664850
rect 139590 664610 139830 664850
rect 139920 664610 140160 664850
rect 140270 664610 140510 664850
rect 140600 664610 140840 664850
rect 140930 664610 141170 664850
rect 141260 664610 141500 664850
rect 141610 664610 141850 664850
rect 141940 664610 142180 664850
rect 142270 664610 142510 664850
rect 142600 664610 142840 664850
rect 142950 664610 143190 664850
rect 143280 664610 143520 664850
rect 143610 664610 143850 664850
rect 143940 664610 144180 664850
rect 144290 664610 144530 664850
rect 133570 664280 133810 664520
rect 133900 664280 134140 664520
rect 134230 664280 134470 664520
rect 134560 664280 134800 664520
rect 134910 664280 135150 664520
rect 135240 664280 135480 664520
rect 135570 664280 135810 664520
rect 135900 664280 136140 664520
rect 136250 664280 136490 664520
rect 136580 664280 136820 664520
rect 136910 664280 137150 664520
rect 137240 664280 137480 664520
rect 137590 664280 137830 664520
rect 137920 664280 138160 664520
rect 138250 664280 138490 664520
rect 138580 664280 138820 664520
rect 138930 664280 139170 664520
rect 139260 664280 139500 664520
rect 139590 664280 139830 664520
rect 139920 664280 140160 664520
rect 140270 664280 140510 664520
rect 140600 664280 140840 664520
rect 140930 664280 141170 664520
rect 141260 664280 141500 664520
rect 141610 664280 141850 664520
rect 141940 664280 142180 664520
rect 142270 664280 142510 664520
rect 142600 664280 142840 664520
rect 142950 664280 143190 664520
rect 143280 664280 143520 664520
rect 143610 664280 143850 664520
rect 143940 664280 144180 664520
rect 144290 664280 144530 664520
rect 133570 663950 133810 664190
rect 133900 663950 134140 664190
rect 134230 663950 134470 664190
rect 134560 663950 134800 664190
rect 134910 663950 135150 664190
rect 135240 663950 135480 664190
rect 135570 663950 135810 664190
rect 135900 663950 136140 664190
rect 136250 663950 136490 664190
rect 136580 663950 136820 664190
rect 136910 663950 137150 664190
rect 137240 663950 137480 664190
rect 137590 663950 137830 664190
rect 137920 663950 138160 664190
rect 138250 663950 138490 664190
rect 138580 663950 138820 664190
rect 138930 663950 139170 664190
rect 139260 663950 139500 664190
rect 139590 663950 139830 664190
rect 139920 663950 140160 664190
rect 140270 663950 140510 664190
rect 140600 663950 140840 664190
rect 140930 663950 141170 664190
rect 141260 663950 141500 664190
rect 141610 663950 141850 664190
rect 141940 663950 142180 664190
rect 142270 663950 142510 664190
rect 142600 663950 142840 664190
rect 142950 663950 143190 664190
rect 143280 663950 143520 664190
rect 143610 663950 143850 664190
rect 143940 663950 144180 664190
rect 144290 663950 144530 664190
rect 133570 663620 133810 663860
rect 133900 663620 134140 663860
rect 134230 663620 134470 663860
rect 134560 663620 134800 663860
rect 134910 663620 135150 663860
rect 135240 663620 135480 663860
rect 135570 663620 135810 663860
rect 135900 663620 136140 663860
rect 136250 663620 136490 663860
rect 136580 663620 136820 663860
rect 136910 663620 137150 663860
rect 137240 663620 137480 663860
rect 137590 663620 137830 663860
rect 137920 663620 138160 663860
rect 138250 663620 138490 663860
rect 138580 663620 138820 663860
rect 138930 663620 139170 663860
rect 139260 663620 139500 663860
rect 139590 663620 139830 663860
rect 139920 663620 140160 663860
rect 140270 663620 140510 663860
rect 140600 663620 140840 663860
rect 140930 663620 141170 663860
rect 141260 663620 141500 663860
rect 141610 663620 141850 663860
rect 141940 663620 142180 663860
rect 142270 663620 142510 663860
rect 142600 663620 142840 663860
rect 142950 663620 143190 663860
rect 143280 663620 143520 663860
rect 143610 663620 143850 663860
rect 143940 663620 144180 663860
rect 144290 663620 144530 663860
rect 133570 663270 133810 663510
rect 133900 663270 134140 663510
rect 134230 663270 134470 663510
rect 134560 663270 134800 663510
rect 134910 663270 135150 663510
rect 135240 663270 135480 663510
rect 135570 663270 135810 663510
rect 135900 663270 136140 663510
rect 136250 663270 136490 663510
rect 136580 663270 136820 663510
rect 136910 663270 137150 663510
rect 137240 663270 137480 663510
rect 137590 663270 137830 663510
rect 137920 663270 138160 663510
rect 138250 663270 138490 663510
rect 138580 663270 138820 663510
rect 138930 663270 139170 663510
rect 139260 663270 139500 663510
rect 139590 663270 139830 663510
rect 139920 663270 140160 663510
rect 140270 663270 140510 663510
rect 140600 663270 140840 663510
rect 140930 663270 141170 663510
rect 141260 663270 141500 663510
rect 141610 663270 141850 663510
rect 141940 663270 142180 663510
rect 142270 663270 142510 663510
rect 142600 663270 142840 663510
rect 142950 663270 143190 663510
rect 143280 663270 143520 663510
rect 143610 663270 143850 663510
rect 143940 663270 144180 663510
rect 144290 663270 144530 663510
rect 133570 662940 133810 663180
rect 133900 662940 134140 663180
rect 134230 662940 134470 663180
rect 134560 662940 134800 663180
rect 134910 662940 135150 663180
rect 135240 662940 135480 663180
rect 135570 662940 135810 663180
rect 135900 662940 136140 663180
rect 136250 662940 136490 663180
rect 136580 662940 136820 663180
rect 136910 662940 137150 663180
rect 137240 662940 137480 663180
rect 137590 662940 137830 663180
rect 137920 662940 138160 663180
rect 138250 662940 138490 663180
rect 138580 662940 138820 663180
rect 138930 662940 139170 663180
rect 139260 662940 139500 663180
rect 139590 662940 139830 663180
rect 139920 662940 140160 663180
rect 140270 662940 140510 663180
rect 140600 662940 140840 663180
rect 140930 662940 141170 663180
rect 141260 662940 141500 663180
rect 141610 662940 141850 663180
rect 141940 662940 142180 663180
rect 142270 662940 142510 663180
rect 142600 662940 142840 663180
rect 142950 662940 143190 663180
rect 143280 662940 143520 663180
rect 143610 662940 143850 663180
rect 143940 662940 144180 663180
rect 144290 662940 144530 663180
rect 133570 662610 133810 662850
rect 133900 662610 134140 662850
rect 134230 662610 134470 662850
rect 134560 662610 134800 662850
rect 134910 662610 135150 662850
rect 135240 662610 135480 662850
rect 135570 662610 135810 662850
rect 135900 662610 136140 662850
rect 136250 662610 136490 662850
rect 136580 662610 136820 662850
rect 136910 662610 137150 662850
rect 137240 662610 137480 662850
rect 137590 662610 137830 662850
rect 137920 662610 138160 662850
rect 138250 662610 138490 662850
rect 138580 662610 138820 662850
rect 138930 662610 139170 662850
rect 139260 662610 139500 662850
rect 139590 662610 139830 662850
rect 139920 662610 140160 662850
rect 140270 662610 140510 662850
rect 140600 662610 140840 662850
rect 140930 662610 141170 662850
rect 141260 662610 141500 662850
rect 141610 662610 141850 662850
rect 141940 662610 142180 662850
rect 142270 662610 142510 662850
rect 142600 662610 142840 662850
rect 142950 662610 143190 662850
rect 143280 662610 143520 662850
rect 143610 662610 143850 662850
rect 143940 662610 144180 662850
rect 144290 662610 144530 662850
rect 133570 662280 133810 662520
rect 133900 662280 134140 662520
rect 134230 662280 134470 662520
rect 134560 662280 134800 662520
rect 134910 662280 135150 662520
rect 135240 662280 135480 662520
rect 135570 662280 135810 662520
rect 135900 662280 136140 662520
rect 136250 662280 136490 662520
rect 136580 662280 136820 662520
rect 136910 662280 137150 662520
rect 137240 662280 137480 662520
rect 137590 662280 137830 662520
rect 137920 662280 138160 662520
rect 138250 662280 138490 662520
rect 138580 662280 138820 662520
rect 138930 662280 139170 662520
rect 139260 662280 139500 662520
rect 139590 662280 139830 662520
rect 139920 662280 140160 662520
rect 140270 662280 140510 662520
rect 140600 662280 140840 662520
rect 140930 662280 141170 662520
rect 141260 662280 141500 662520
rect 141610 662280 141850 662520
rect 141940 662280 142180 662520
rect 142270 662280 142510 662520
rect 142600 662280 142840 662520
rect 142950 662280 143190 662520
rect 143280 662280 143520 662520
rect 143610 662280 143850 662520
rect 143940 662280 144180 662520
rect 144290 662280 144530 662520
rect 133570 661930 133810 662170
rect 133900 661930 134140 662170
rect 134230 661930 134470 662170
rect 134560 661930 134800 662170
rect 134910 661930 135150 662170
rect 135240 661930 135480 662170
rect 135570 661930 135810 662170
rect 135900 661930 136140 662170
rect 136250 661930 136490 662170
rect 136580 661930 136820 662170
rect 136910 661930 137150 662170
rect 137240 661930 137480 662170
rect 137590 661930 137830 662170
rect 137920 661930 138160 662170
rect 138250 661930 138490 662170
rect 138580 661930 138820 662170
rect 138930 661930 139170 662170
rect 139260 661930 139500 662170
rect 139590 661930 139830 662170
rect 139920 661930 140160 662170
rect 140270 661930 140510 662170
rect 140600 661930 140840 662170
rect 140930 661930 141170 662170
rect 141260 661930 141500 662170
rect 141610 661930 141850 662170
rect 141940 661930 142180 662170
rect 142270 661930 142510 662170
rect 142600 661930 142840 662170
rect 142950 661930 143190 662170
rect 143280 661930 143520 662170
rect 143610 661930 143850 662170
rect 143940 661930 144180 662170
rect 144290 661930 144530 662170
rect 133570 661600 133810 661840
rect 133900 661600 134140 661840
rect 134230 661600 134470 661840
rect 134560 661600 134800 661840
rect 134910 661600 135150 661840
rect 135240 661600 135480 661840
rect 135570 661600 135810 661840
rect 135900 661600 136140 661840
rect 136250 661600 136490 661840
rect 136580 661600 136820 661840
rect 136910 661600 137150 661840
rect 137240 661600 137480 661840
rect 137590 661600 137830 661840
rect 137920 661600 138160 661840
rect 138250 661600 138490 661840
rect 138580 661600 138820 661840
rect 138930 661600 139170 661840
rect 139260 661600 139500 661840
rect 139590 661600 139830 661840
rect 139920 661600 140160 661840
rect 140270 661600 140510 661840
rect 140600 661600 140840 661840
rect 140930 661600 141170 661840
rect 141260 661600 141500 661840
rect 141610 661600 141850 661840
rect 141940 661600 142180 661840
rect 142270 661600 142510 661840
rect 142600 661600 142840 661840
rect 142950 661600 143190 661840
rect 143280 661600 143520 661840
rect 143610 661600 143850 661840
rect 143940 661600 144180 661840
rect 144290 661600 144530 661840
rect 133570 661270 133810 661510
rect 133900 661270 134140 661510
rect 134230 661270 134470 661510
rect 134560 661270 134800 661510
rect 134910 661270 135150 661510
rect 135240 661270 135480 661510
rect 135570 661270 135810 661510
rect 135900 661270 136140 661510
rect 136250 661270 136490 661510
rect 136580 661270 136820 661510
rect 136910 661270 137150 661510
rect 137240 661270 137480 661510
rect 137590 661270 137830 661510
rect 137920 661270 138160 661510
rect 138250 661270 138490 661510
rect 138580 661270 138820 661510
rect 138930 661270 139170 661510
rect 139260 661270 139500 661510
rect 139590 661270 139830 661510
rect 139920 661270 140160 661510
rect 140270 661270 140510 661510
rect 140600 661270 140840 661510
rect 140930 661270 141170 661510
rect 141260 661270 141500 661510
rect 141610 661270 141850 661510
rect 141940 661270 142180 661510
rect 142270 661270 142510 661510
rect 142600 661270 142840 661510
rect 142950 661270 143190 661510
rect 143280 661270 143520 661510
rect 143610 661270 143850 661510
rect 143940 661270 144180 661510
rect 144290 661270 144530 661510
rect 133570 660940 133810 661180
rect 133900 660940 134140 661180
rect 134230 660940 134470 661180
rect 134560 660940 134800 661180
rect 134910 660940 135150 661180
rect 135240 660940 135480 661180
rect 135570 660940 135810 661180
rect 135900 660940 136140 661180
rect 136250 660940 136490 661180
rect 136580 660940 136820 661180
rect 136910 660940 137150 661180
rect 137240 660940 137480 661180
rect 137590 660940 137830 661180
rect 137920 660940 138160 661180
rect 138250 660940 138490 661180
rect 138580 660940 138820 661180
rect 138930 660940 139170 661180
rect 139260 660940 139500 661180
rect 139590 660940 139830 661180
rect 139920 660940 140160 661180
rect 140270 660940 140510 661180
rect 140600 660940 140840 661180
rect 140930 660940 141170 661180
rect 141260 660940 141500 661180
rect 141610 660940 141850 661180
rect 141940 660940 142180 661180
rect 142270 660940 142510 661180
rect 142600 660940 142840 661180
rect 142950 660940 143190 661180
rect 143280 660940 143520 661180
rect 143610 660940 143850 661180
rect 143940 660940 144180 661180
rect 144290 660940 144530 661180
rect 144950 671660 145190 671900
rect 145280 671660 145520 671900
rect 145610 671660 145850 671900
rect 145940 671660 146180 671900
rect 146290 671660 146530 671900
rect 146620 671660 146860 671900
rect 146950 671660 147190 671900
rect 147280 671660 147520 671900
rect 147630 671660 147870 671900
rect 147960 671660 148200 671900
rect 148290 671660 148530 671900
rect 148620 671660 148860 671900
rect 148970 671660 149210 671900
rect 149300 671660 149540 671900
rect 149630 671660 149870 671900
rect 149960 671660 150200 671900
rect 150310 671660 150550 671900
rect 150640 671660 150880 671900
rect 150970 671660 151210 671900
rect 151300 671660 151540 671900
rect 151650 671660 151890 671900
rect 151980 671660 152220 671900
rect 152310 671660 152550 671900
rect 152640 671660 152880 671900
rect 152990 671660 153230 671900
rect 153320 671660 153560 671900
rect 153650 671660 153890 671900
rect 153980 671660 154220 671900
rect 154330 671660 154570 671900
rect 154660 671660 154900 671900
rect 154990 671660 155230 671900
rect 155320 671660 155560 671900
rect 155670 671660 155910 671900
rect 144950 671310 145190 671550
rect 145280 671310 145520 671550
rect 145610 671310 145850 671550
rect 145940 671310 146180 671550
rect 146290 671310 146530 671550
rect 146620 671310 146860 671550
rect 146950 671310 147190 671550
rect 147280 671310 147520 671550
rect 147630 671310 147870 671550
rect 147960 671310 148200 671550
rect 148290 671310 148530 671550
rect 148620 671310 148860 671550
rect 148970 671310 149210 671550
rect 149300 671310 149540 671550
rect 149630 671310 149870 671550
rect 149960 671310 150200 671550
rect 150310 671310 150550 671550
rect 150640 671310 150880 671550
rect 150970 671310 151210 671550
rect 151300 671310 151540 671550
rect 151650 671310 151890 671550
rect 151980 671310 152220 671550
rect 152310 671310 152550 671550
rect 152640 671310 152880 671550
rect 152990 671310 153230 671550
rect 153320 671310 153560 671550
rect 153650 671310 153890 671550
rect 153980 671310 154220 671550
rect 154330 671310 154570 671550
rect 154660 671310 154900 671550
rect 154990 671310 155230 671550
rect 155320 671310 155560 671550
rect 155670 671310 155910 671550
rect 144950 670980 145190 671220
rect 145280 670980 145520 671220
rect 145610 670980 145850 671220
rect 145940 670980 146180 671220
rect 146290 670980 146530 671220
rect 146620 670980 146860 671220
rect 146950 670980 147190 671220
rect 147280 670980 147520 671220
rect 147630 670980 147870 671220
rect 147960 670980 148200 671220
rect 148290 670980 148530 671220
rect 148620 670980 148860 671220
rect 148970 670980 149210 671220
rect 149300 670980 149540 671220
rect 149630 670980 149870 671220
rect 149960 670980 150200 671220
rect 150310 670980 150550 671220
rect 150640 670980 150880 671220
rect 150970 670980 151210 671220
rect 151300 670980 151540 671220
rect 151650 670980 151890 671220
rect 151980 670980 152220 671220
rect 152310 670980 152550 671220
rect 152640 670980 152880 671220
rect 152990 670980 153230 671220
rect 153320 670980 153560 671220
rect 153650 670980 153890 671220
rect 153980 670980 154220 671220
rect 154330 670980 154570 671220
rect 154660 670980 154900 671220
rect 154990 670980 155230 671220
rect 155320 670980 155560 671220
rect 155670 670980 155910 671220
rect 144950 670650 145190 670890
rect 145280 670650 145520 670890
rect 145610 670650 145850 670890
rect 145940 670650 146180 670890
rect 146290 670650 146530 670890
rect 146620 670650 146860 670890
rect 146950 670650 147190 670890
rect 147280 670650 147520 670890
rect 147630 670650 147870 670890
rect 147960 670650 148200 670890
rect 148290 670650 148530 670890
rect 148620 670650 148860 670890
rect 148970 670650 149210 670890
rect 149300 670650 149540 670890
rect 149630 670650 149870 670890
rect 149960 670650 150200 670890
rect 150310 670650 150550 670890
rect 150640 670650 150880 670890
rect 150970 670650 151210 670890
rect 151300 670650 151540 670890
rect 151650 670650 151890 670890
rect 151980 670650 152220 670890
rect 152310 670650 152550 670890
rect 152640 670650 152880 670890
rect 152990 670650 153230 670890
rect 153320 670650 153560 670890
rect 153650 670650 153890 670890
rect 153980 670650 154220 670890
rect 154330 670650 154570 670890
rect 154660 670650 154900 670890
rect 154990 670650 155230 670890
rect 155320 670650 155560 670890
rect 155670 670650 155910 670890
rect 144950 670320 145190 670560
rect 145280 670320 145520 670560
rect 145610 670320 145850 670560
rect 145940 670320 146180 670560
rect 146290 670320 146530 670560
rect 146620 670320 146860 670560
rect 146950 670320 147190 670560
rect 147280 670320 147520 670560
rect 147630 670320 147870 670560
rect 147960 670320 148200 670560
rect 148290 670320 148530 670560
rect 148620 670320 148860 670560
rect 148970 670320 149210 670560
rect 149300 670320 149540 670560
rect 149630 670320 149870 670560
rect 149960 670320 150200 670560
rect 150310 670320 150550 670560
rect 150640 670320 150880 670560
rect 150970 670320 151210 670560
rect 151300 670320 151540 670560
rect 151650 670320 151890 670560
rect 151980 670320 152220 670560
rect 152310 670320 152550 670560
rect 152640 670320 152880 670560
rect 152990 670320 153230 670560
rect 153320 670320 153560 670560
rect 153650 670320 153890 670560
rect 153980 670320 154220 670560
rect 154330 670320 154570 670560
rect 154660 670320 154900 670560
rect 154990 670320 155230 670560
rect 155320 670320 155560 670560
rect 155670 670320 155910 670560
rect 144950 669970 145190 670210
rect 145280 669970 145520 670210
rect 145610 669970 145850 670210
rect 145940 669970 146180 670210
rect 146290 669970 146530 670210
rect 146620 669970 146860 670210
rect 146950 669970 147190 670210
rect 147280 669970 147520 670210
rect 147630 669970 147870 670210
rect 147960 669970 148200 670210
rect 148290 669970 148530 670210
rect 148620 669970 148860 670210
rect 148970 669970 149210 670210
rect 149300 669970 149540 670210
rect 149630 669970 149870 670210
rect 149960 669970 150200 670210
rect 150310 669970 150550 670210
rect 150640 669970 150880 670210
rect 150970 669970 151210 670210
rect 151300 669970 151540 670210
rect 151650 669970 151890 670210
rect 151980 669970 152220 670210
rect 152310 669970 152550 670210
rect 152640 669970 152880 670210
rect 152990 669970 153230 670210
rect 153320 669970 153560 670210
rect 153650 669970 153890 670210
rect 153980 669970 154220 670210
rect 154330 669970 154570 670210
rect 154660 669970 154900 670210
rect 154990 669970 155230 670210
rect 155320 669970 155560 670210
rect 155670 669970 155910 670210
rect 144950 669640 145190 669880
rect 145280 669640 145520 669880
rect 145610 669640 145850 669880
rect 145940 669640 146180 669880
rect 146290 669640 146530 669880
rect 146620 669640 146860 669880
rect 146950 669640 147190 669880
rect 147280 669640 147520 669880
rect 147630 669640 147870 669880
rect 147960 669640 148200 669880
rect 148290 669640 148530 669880
rect 148620 669640 148860 669880
rect 148970 669640 149210 669880
rect 149300 669640 149540 669880
rect 149630 669640 149870 669880
rect 149960 669640 150200 669880
rect 150310 669640 150550 669880
rect 150640 669640 150880 669880
rect 150970 669640 151210 669880
rect 151300 669640 151540 669880
rect 151650 669640 151890 669880
rect 151980 669640 152220 669880
rect 152310 669640 152550 669880
rect 152640 669640 152880 669880
rect 152990 669640 153230 669880
rect 153320 669640 153560 669880
rect 153650 669640 153890 669880
rect 153980 669640 154220 669880
rect 154330 669640 154570 669880
rect 154660 669640 154900 669880
rect 154990 669640 155230 669880
rect 155320 669640 155560 669880
rect 155670 669640 155910 669880
rect 144950 669310 145190 669550
rect 145280 669310 145520 669550
rect 145610 669310 145850 669550
rect 145940 669310 146180 669550
rect 146290 669310 146530 669550
rect 146620 669310 146860 669550
rect 146950 669310 147190 669550
rect 147280 669310 147520 669550
rect 147630 669310 147870 669550
rect 147960 669310 148200 669550
rect 148290 669310 148530 669550
rect 148620 669310 148860 669550
rect 148970 669310 149210 669550
rect 149300 669310 149540 669550
rect 149630 669310 149870 669550
rect 149960 669310 150200 669550
rect 150310 669310 150550 669550
rect 150640 669310 150880 669550
rect 150970 669310 151210 669550
rect 151300 669310 151540 669550
rect 151650 669310 151890 669550
rect 151980 669310 152220 669550
rect 152310 669310 152550 669550
rect 152640 669310 152880 669550
rect 152990 669310 153230 669550
rect 153320 669310 153560 669550
rect 153650 669310 153890 669550
rect 153980 669310 154220 669550
rect 154330 669310 154570 669550
rect 154660 669310 154900 669550
rect 154990 669310 155230 669550
rect 155320 669310 155560 669550
rect 155670 669310 155910 669550
rect 144950 668980 145190 669220
rect 145280 668980 145520 669220
rect 145610 668980 145850 669220
rect 145940 668980 146180 669220
rect 146290 668980 146530 669220
rect 146620 668980 146860 669220
rect 146950 668980 147190 669220
rect 147280 668980 147520 669220
rect 147630 668980 147870 669220
rect 147960 668980 148200 669220
rect 148290 668980 148530 669220
rect 148620 668980 148860 669220
rect 148970 668980 149210 669220
rect 149300 668980 149540 669220
rect 149630 668980 149870 669220
rect 149960 668980 150200 669220
rect 150310 668980 150550 669220
rect 150640 668980 150880 669220
rect 150970 668980 151210 669220
rect 151300 668980 151540 669220
rect 151650 668980 151890 669220
rect 151980 668980 152220 669220
rect 152310 668980 152550 669220
rect 152640 668980 152880 669220
rect 152990 668980 153230 669220
rect 153320 668980 153560 669220
rect 153650 668980 153890 669220
rect 153980 668980 154220 669220
rect 154330 668980 154570 669220
rect 154660 668980 154900 669220
rect 154990 668980 155230 669220
rect 155320 668980 155560 669220
rect 155670 668980 155910 669220
rect 144950 668630 145190 668870
rect 145280 668630 145520 668870
rect 145610 668630 145850 668870
rect 145940 668630 146180 668870
rect 146290 668630 146530 668870
rect 146620 668630 146860 668870
rect 146950 668630 147190 668870
rect 147280 668630 147520 668870
rect 147630 668630 147870 668870
rect 147960 668630 148200 668870
rect 148290 668630 148530 668870
rect 148620 668630 148860 668870
rect 148970 668630 149210 668870
rect 149300 668630 149540 668870
rect 149630 668630 149870 668870
rect 149960 668630 150200 668870
rect 150310 668630 150550 668870
rect 150640 668630 150880 668870
rect 150970 668630 151210 668870
rect 151300 668630 151540 668870
rect 151650 668630 151890 668870
rect 151980 668630 152220 668870
rect 152310 668630 152550 668870
rect 152640 668630 152880 668870
rect 152990 668630 153230 668870
rect 153320 668630 153560 668870
rect 153650 668630 153890 668870
rect 153980 668630 154220 668870
rect 154330 668630 154570 668870
rect 154660 668630 154900 668870
rect 154990 668630 155230 668870
rect 155320 668630 155560 668870
rect 155670 668630 155910 668870
rect 144950 668300 145190 668540
rect 145280 668300 145520 668540
rect 145610 668300 145850 668540
rect 145940 668300 146180 668540
rect 146290 668300 146530 668540
rect 146620 668300 146860 668540
rect 146950 668300 147190 668540
rect 147280 668300 147520 668540
rect 147630 668300 147870 668540
rect 147960 668300 148200 668540
rect 148290 668300 148530 668540
rect 148620 668300 148860 668540
rect 148970 668300 149210 668540
rect 149300 668300 149540 668540
rect 149630 668300 149870 668540
rect 149960 668300 150200 668540
rect 150310 668300 150550 668540
rect 150640 668300 150880 668540
rect 150970 668300 151210 668540
rect 151300 668300 151540 668540
rect 151650 668300 151890 668540
rect 151980 668300 152220 668540
rect 152310 668300 152550 668540
rect 152640 668300 152880 668540
rect 152990 668300 153230 668540
rect 153320 668300 153560 668540
rect 153650 668300 153890 668540
rect 153980 668300 154220 668540
rect 154330 668300 154570 668540
rect 154660 668300 154900 668540
rect 154990 668300 155230 668540
rect 155320 668300 155560 668540
rect 155670 668300 155910 668540
rect 144950 667970 145190 668210
rect 145280 667970 145520 668210
rect 145610 667970 145850 668210
rect 145940 667970 146180 668210
rect 146290 667970 146530 668210
rect 146620 667970 146860 668210
rect 146950 667970 147190 668210
rect 147280 667970 147520 668210
rect 147630 667970 147870 668210
rect 147960 667970 148200 668210
rect 148290 667970 148530 668210
rect 148620 667970 148860 668210
rect 148970 667970 149210 668210
rect 149300 667970 149540 668210
rect 149630 667970 149870 668210
rect 149960 667970 150200 668210
rect 150310 667970 150550 668210
rect 150640 667970 150880 668210
rect 150970 667970 151210 668210
rect 151300 667970 151540 668210
rect 151650 667970 151890 668210
rect 151980 667970 152220 668210
rect 152310 667970 152550 668210
rect 152640 667970 152880 668210
rect 152990 667970 153230 668210
rect 153320 667970 153560 668210
rect 153650 667970 153890 668210
rect 153980 667970 154220 668210
rect 154330 667970 154570 668210
rect 154660 667970 154900 668210
rect 154990 667970 155230 668210
rect 155320 667970 155560 668210
rect 155670 667970 155910 668210
rect 144950 667640 145190 667880
rect 145280 667640 145520 667880
rect 145610 667640 145850 667880
rect 145940 667640 146180 667880
rect 146290 667640 146530 667880
rect 146620 667640 146860 667880
rect 146950 667640 147190 667880
rect 147280 667640 147520 667880
rect 147630 667640 147870 667880
rect 147960 667640 148200 667880
rect 148290 667640 148530 667880
rect 148620 667640 148860 667880
rect 148970 667640 149210 667880
rect 149300 667640 149540 667880
rect 149630 667640 149870 667880
rect 149960 667640 150200 667880
rect 150310 667640 150550 667880
rect 150640 667640 150880 667880
rect 150970 667640 151210 667880
rect 151300 667640 151540 667880
rect 151650 667640 151890 667880
rect 151980 667640 152220 667880
rect 152310 667640 152550 667880
rect 152640 667640 152880 667880
rect 152990 667640 153230 667880
rect 153320 667640 153560 667880
rect 153650 667640 153890 667880
rect 153980 667640 154220 667880
rect 154330 667640 154570 667880
rect 154660 667640 154900 667880
rect 154990 667640 155230 667880
rect 155320 667640 155560 667880
rect 155670 667640 155910 667880
rect 144950 667290 145190 667530
rect 145280 667290 145520 667530
rect 145610 667290 145850 667530
rect 145940 667290 146180 667530
rect 146290 667290 146530 667530
rect 146620 667290 146860 667530
rect 146950 667290 147190 667530
rect 147280 667290 147520 667530
rect 147630 667290 147870 667530
rect 147960 667290 148200 667530
rect 148290 667290 148530 667530
rect 148620 667290 148860 667530
rect 148970 667290 149210 667530
rect 149300 667290 149540 667530
rect 149630 667290 149870 667530
rect 149960 667290 150200 667530
rect 150310 667290 150550 667530
rect 150640 667290 150880 667530
rect 150970 667290 151210 667530
rect 151300 667290 151540 667530
rect 151650 667290 151890 667530
rect 151980 667290 152220 667530
rect 152310 667290 152550 667530
rect 152640 667290 152880 667530
rect 152990 667290 153230 667530
rect 153320 667290 153560 667530
rect 153650 667290 153890 667530
rect 153980 667290 154220 667530
rect 154330 667290 154570 667530
rect 154660 667290 154900 667530
rect 154990 667290 155230 667530
rect 155320 667290 155560 667530
rect 155670 667290 155910 667530
rect 144950 666960 145190 667200
rect 145280 666960 145520 667200
rect 145610 666960 145850 667200
rect 145940 666960 146180 667200
rect 146290 666960 146530 667200
rect 146620 666960 146860 667200
rect 146950 666960 147190 667200
rect 147280 666960 147520 667200
rect 147630 666960 147870 667200
rect 147960 666960 148200 667200
rect 148290 666960 148530 667200
rect 148620 666960 148860 667200
rect 148970 666960 149210 667200
rect 149300 666960 149540 667200
rect 149630 666960 149870 667200
rect 149960 666960 150200 667200
rect 150310 666960 150550 667200
rect 150640 666960 150880 667200
rect 150970 666960 151210 667200
rect 151300 666960 151540 667200
rect 151650 666960 151890 667200
rect 151980 666960 152220 667200
rect 152310 666960 152550 667200
rect 152640 666960 152880 667200
rect 152990 666960 153230 667200
rect 153320 666960 153560 667200
rect 153650 666960 153890 667200
rect 153980 666960 154220 667200
rect 154330 666960 154570 667200
rect 154660 666960 154900 667200
rect 154990 666960 155230 667200
rect 155320 666960 155560 667200
rect 155670 666960 155910 667200
rect 144950 666630 145190 666870
rect 145280 666630 145520 666870
rect 145610 666630 145850 666870
rect 145940 666630 146180 666870
rect 146290 666630 146530 666870
rect 146620 666630 146860 666870
rect 146950 666630 147190 666870
rect 147280 666630 147520 666870
rect 147630 666630 147870 666870
rect 147960 666630 148200 666870
rect 148290 666630 148530 666870
rect 148620 666630 148860 666870
rect 148970 666630 149210 666870
rect 149300 666630 149540 666870
rect 149630 666630 149870 666870
rect 149960 666630 150200 666870
rect 150310 666630 150550 666870
rect 150640 666630 150880 666870
rect 150970 666630 151210 666870
rect 151300 666630 151540 666870
rect 151650 666630 151890 666870
rect 151980 666630 152220 666870
rect 152310 666630 152550 666870
rect 152640 666630 152880 666870
rect 152990 666630 153230 666870
rect 153320 666630 153560 666870
rect 153650 666630 153890 666870
rect 153980 666630 154220 666870
rect 154330 666630 154570 666870
rect 154660 666630 154900 666870
rect 154990 666630 155230 666870
rect 155320 666630 155560 666870
rect 155670 666630 155910 666870
rect 144950 666300 145190 666540
rect 145280 666300 145520 666540
rect 145610 666300 145850 666540
rect 145940 666300 146180 666540
rect 146290 666300 146530 666540
rect 146620 666300 146860 666540
rect 146950 666300 147190 666540
rect 147280 666300 147520 666540
rect 147630 666300 147870 666540
rect 147960 666300 148200 666540
rect 148290 666300 148530 666540
rect 148620 666300 148860 666540
rect 148970 666300 149210 666540
rect 149300 666300 149540 666540
rect 149630 666300 149870 666540
rect 149960 666300 150200 666540
rect 150310 666300 150550 666540
rect 150640 666300 150880 666540
rect 150970 666300 151210 666540
rect 151300 666300 151540 666540
rect 151650 666300 151890 666540
rect 151980 666300 152220 666540
rect 152310 666300 152550 666540
rect 152640 666300 152880 666540
rect 152990 666300 153230 666540
rect 153320 666300 153560 666540
rect 153650 666300 153890 666540
rect 153980 666300 154220 666540
rect 154330 666300 154570 666540
rect 154660 666300 154900 666540
rect 154990 666300 155230 666540
rect 155320 666300 155560 666540
rect 155670 666300 155910 666540
rect 144950 665950 145190 666190
rect 145280 665950 145520 666190
rect 145610 665950 145850 666190
rect 145940 665950 146180 666190
rect 146290 665950 146530 666190
rect 146620 665950 146860 666190
rect 146950 665950 147190 666190
rect 147280 665950 147520 666190
rect 147630 665950 147870 666190
rect 147960 665950 148200 666190
rect 148290 665950 148530 666190
rect 148620 665950 148860 666190
rect 148970 665950 149210 666190
rect 149300 665950 149540 666190
rect 149630 665950 149870 666190
rect 149960 665950 150200 666190
rect 150310 665950 150550 666190
rect 150640 665950 150880 666190
rect 150970 665950 151210 666190
rect 151300 665950 151540 666190
rect 151650 665950 151890 666190
rect 151980 665950 152220 666190
rect 152310 665950 152550 666190
rect 152640 665950 152880 666190
rect 152990 665950 153230 666190
rect 153320 665950 153560 666190
rect 153650 665950 153890 666190
rect 153980 665950 154220 666190
rect 154330 665950 154570 666190
rect 154660 665950 154900 666190
rect 154990 665950 155230 666190
rect 155320 665950 155560 666190
rect 155670 665950 155910 666190
rect 144950 665620 145190 665860
rect 145280 665620 145520 665860
rect 145610 665620 145850 665860
rect 145940 665620 146180 665860
rect 146290 665620 146530 665860
rect 146620 665620 146860 665860
rect 146950 665620 147190 665860
rect 147280 665620 147520 665860
rect 147630 665620 147870 665860
rect 147960 665620 148200 665860
rect 148290 665620 148530 665860
rect 148620 665620 148860 665860
rect 148970 665620 149210 665860
rect 149300 665620 149540 665860
rect 149630 665620 149870 665860
rect 149960 665620 150200 665860
rect 150310 665620 150550 665860
rect 150640 665620 150880 665860
rect 150970 665620 151210 665860
rect 151300 665620 151540 665860
rect 151650 665620 151890 665860
rect 151980 665620 152220 665860
rect 152310 665620 152550 665860
rect 152640 665620 152880 665860
rect 152990 665620 153230 665860
rect 153320 665620 153560 665860
rect 153650 665620 153890 665860
rect 153980 665620 154220 665860
rect 154330 665620 154570 665860
rect 154660 665620 154900 665860
rect 154990 665620 155230 665860
rect 155320 665620 155560 665860
rect 155670 665620 155910 665860
rect 144950 665290 145190 665530
rect 145280 665290 145520 665530
rect 145610 665290 145850 665530
rect 145940 665290 146180 665530
rect 146290 665290 146530 665530
rect 146620 665290 146860 665530
rect 146950 665290 147190 665530
rect 147280 665290 147520 665530
rect 147630 665290 147870 665530
rect 147960 665290 148200 665530
rect 148290 665290 148530 665530
rect 148620 665290 148860 665530
rect 148970 665290 149210 665530
rect 149300 665290 149540 665530
rect 149630 665290 149870 665530
rect 149960 665290 150200 665530
rect 150310 665290 150550 665530
rect 150640 665290 150880 665530
rect 150970 665290 151210 665530
rect 151300 665290 151540 665530
rect 151650 665290 151890 665530
rect 151980 665290 152220 665530
rect 152310 665290 152550 665530
rect 152640 665290 152880 665530
rect 152990 665290 153230 665530
rect 153320 665290 153560 665530
rect 153650 665290 153890 665530
rect 153980 665290 154220 665530
rect 154330 665290 154570 665530
rect 154660 665290 154900 665530
rect 154990 665290 155230 665530
rect 155320 665290 155560 665530
rect 155670 665290 155910 665530
rect 144950 664960 145190 665200
rect 145280 664960 145520 665200
rect 145610 664960 145850 665200
rect 145940 664960 146180 665200
rect 146290 664960 146530 665200
rect 146620 664960 146860 665200
rect 146950 664960 147190 665200
rect 147280 664960 147520 665200
rect 147630 664960 147870 665200
rect 147960 664960 148200 665200
rect 148290 664960 148530 665200
rect 148620 664960 148860 665200
rect 148970 664960 149210 665200
rect 149300 664960 149540 665200
rect 149630 664960 149870 665200
rect 149960 664960 150200 665200
rect 150310 664960 150550 665200
rect 150640 664960 150880 665200
rect 150970 664960 151210 665200
rect 151300 664960 151540 665200
rect 151650 664960 151890 665200
rect 151980 664960 152220 665200
rect 152310 664960 152550 665200
rect 152640 664960 152880 665200
rect 152990 664960 153230 665200
rect 153320 664960 153560 665200
rect 153650 664960 153890 665200
rect 153980 664960 154220 665200
rect 154330 664960 154570 665200
rect 154660 664960 154900 665200
rect 154990 664960 155230 665200
rect 155320 664960 155560 665200
rect 155670 664960 155910 665200
rect 144950 664610 145190 664850
rect 145280 664610 145520 664850
rect 145610 664610 145850 664850
rect 145940 664610 146180 664850
rect 146290 664610 146530 664850
rect 146620 664610 146860 664850
rect 146950 664610 147190 664850
rect 147280 664610 147520 664850
rect 147630 664610 147870 664850
rect 147960 664610 148200 664850
rect 148290 664610 148530 664850
rect 148620 664610 148860 664850
rect 148970 664610 149210 664850
rect 149300 664610 149540 664850
rect 149630 664610 149870 664850
rect 149960 664610 150200 664850
rect 150310 664610 150550 664850
rect 150640 664610 150880 664850
rect 150970 664610 151210 664850
rect 151300 664610 151540 664850
rect 151650 664610 151890 664850
rect 151980 664610 152220 664850
rect 152310 664610 152550 664850
rect 152640 664610 152880 664850
rect 152990 664610 153230 664850
rect 153320 664610 153560 664850
rect 153650 664610 153890 664850
rect 153980 664610 154220 664850
rect 154330 664610 154570 664850
rect 154660 664610 154900 664850
rect 154990 664610 155230 664850
rect 155320 664610 155560 664850
rect 155670 664610 155910 664850
rect 144950 664280 145190 664520
rect 145280 664280 145520 664520
rect 145610 664280 145850 664520
rect 145940 664280 146180 664520
rect 146290 664280 146530 664520
rect 146620 664280 146860 664520
rect 146950 664280 147190 664520
rect 147280 664280 147520 664520
rect 147630 664280 147870 664520
rect 147960 664280 148200 664520
rect 148290 664280 148530 664520
rect 148620 664280 148860 664520
rect 148970 664280 149210 664520
rect 149300 664280 149540 664520
rect 149630 664280 149870 664520
rect 149960 664280 150200 664520
rect 150310 664280 150550 664520
rect 150640 664280 150880 664520
rect 150970 664280 151210 664520
rect 151300 664280 151540 664520
rect 151650 664280 151890 664520
rect 151980 664280 152220 664520
rect 152310 664280 152550 664520
rect 152640 664280 152880 664520
rect 152990 664280 153230 664520
rect 153320 664280 153560 664520
rect 153650 664280 153890 664520
rect 153980 664280 154220 664520
rect 154330 664280 154570 664520
rect 154660 664280 154900 664520
rect 154990 664280 155230 664520
rect 155320 664280 155560 664520
rect 155670 664280 155910 664520
rect 144950 663950 145190 664190
rect 145280 663950 145520 664190
rect 145610 663950 145850 664190
rect 145940 663950 146180 664190
rect 146290 663950 146530 664190
rect 146620 663950 146860 664190
rect 146950 663950 147190 664190
rect 147280 663950 147520 664190
rect 147630 663950 147870 664190
rect 147960 663950 148200 664190
rect 148290 663950 148530 664190
rect 148620 663950 148860 664190
rect 148970 663950 149210 664190
rect 149300 663950 149540 664190
rect 149630 663950 149870 664190
rect 149960 663950 150200 664190
rect 150310 663950 150550 664190
rect 150640 663950 150880 664190
rect 150970 663950 151210 664190
rect 151300 663950 151540 664190
rect 151650 663950 151890 664190
rect 151980 663950 152220 664190
rect 152310 663950 152550 664190
rect 152640 663950 152880 664190
rect 152990 663950 153230 664190
rect 153320 663950 153560 664190
rect 153650 663950 153890 664190
rect 153980 663950 154220 664190
rect 154330 663950 154570 664190
rect 154660 663950 154900 664190
rect 154990 663950 155230 664190
rect 155320 663950 155560 664190
rect 155670 663950 155910 664190
rect 144950 663620 145190 663860
rect 145280 663620 145520 663860
rect 145610 663620 145850 663860
rect 145940 663620 146180 663860
rect 146290 663620 146530 663860
rect 146620 663620 146860 663860
rect 146950 663620 147190 663860
rect 147280 663620 147520 663860
rect 147630 663620 147870 663860
rect 147960 663620 148200 663860
rect 148290 663620 148530 663860
rect 148620 663620 148860 663860
rect 148970 663620 149210 663860
rect 149300 663620 149540 663860
rect 149630 663620 149870 663860
rect 149960 663620 150200 663860
rect 150310 663620 150550 663860
rect 150640 663620 150880 663860
rect 150970 663620 151210 663860
rect 151300 663620 151540 663860
rect 151650 663620 151890 663860
rect 151980 663620 152220 663860
rect 152310 663620 152550 663860
rect 152640 663620 152880 663860
rect 152990 663620 153230 663860
rect 153320 663620 153560 663860
rect 153650 663620 153890 663860
rect 153980 663620 154220 663860
rect 154330 663620 154570 663860
rect 154660 663620 154900 663860
rect 154990 663620 155230 663860
rect 155320 663620 155560 663860
rect 155670 663620 155910 663860
rect 144950 663270 145190 663510
rect 145280 663270 145520 663510
rect 145610 663270 145850 663510
rect 145940 663270 146180 663510
rect 146290 663270 146530 663510
rect 146620 663270 146860 663510
rect 146950 663270 147190 663510
rect 147280 663270 147520 663510
rect 147630 663270 147870 663510
rect 147960 663270 148200 663510
rect 148290 663270 148530 663510
rect 148620 663270 148860 663510
rect 148970 663270 149210 663510
rect 149300 663270 149540 663510
rect 149630 663270 149870 663510
rect 149960 663270 150200 663510
rect 150310 663270 150550 663510
rect 150640 663270 150880 663510
rect 150970 663270 151210 663510
rect 151300 663270 151540 663510
rect 151650 663270 151890 663510
rect 151980 663270 152220 663510
rect 152310 663270 152550 663510
rect 152640 663270 152880 663510
rect 152990 663270 153230 663510
rect 153320 663270 153560 663510
rect 153650 663270 153890 663510
rect 153980 663270 154220 663510
rect 154330 663270 154570 663510
rect 154660 663270 154900 663510
rect 154990 663270 155230 663510
rect 155320 663270 155560 663510
rect 155670 663270 155910 663510
rect 144950 662940 145190 663180
rect 145280 662940 145520 663180
rect 145610 662940 145850 663180
rect 145940 662940 146180 663180
rect 146290 662940 146530 663180
rect 146620 662940 146860 663180
rect 146950 662940 147190 663180
rect 147280 662940 147520 663180
rect 147630 662940 147870 663180
rect 147960 662940 148200 663180
rect 148290 662940 148530 663180
rect 148620 662940 148860 663180
rect 148970 662940 149210 663180
rect 149300 662940 149540 663180
rect 149630 662940 149870 663180
rect 149960 662940 150200 663180
rect 150310 662940 150550 663180
rect 150640 662940 150880 663180
rect 150970 662940 151210 663180
rect 151300 662940 151540 663180
rect 151650 662940 151890 663180
rect 151980 662940 152220 663180
rect 152310 662940 152550 663180
rect 152640 662940 152880 663180
rect 152990 662940 153230 663180
rect 153320 662940 153560 663180
rect 153650 662940 153890 663180
rect 153980 662940 154220 663180
rect 154330 662940 154570 663180
rect 154660 662940 154900 663180
rect 154990 662940 155230 663180
rect 155320 662940 155560 663180
rect 155670 662940 155910 663180
rect 144950 662610 145190 662850
rect 145280 662610 145520 662850
rect 145610 662610 145850 662850
rect 145940 662610 146180 662850
rect 146290 662610 146530 662850
rect 146620 662610 146860 662850
rect 146950 662610 147190 662850
rect 147280 662610 147520 662850
rect 147630 662610 147870 662850
rect 147960 662610 148200 662850
rect 148290 662610 148530 662850
rect 148620 662610 148860 662850
rect 148970 662610 149210 662850
rect 149300 662610 149540 662850
rect 149630 662610 149870 662850
rect 149960 662610 150200 662850
rect 150310 662610 150550 662850
rect 150640 662610 150880 662850
rect 150970 662610 151210 662850
rect 151300 662610 151540 662850
rect 151650 662610 151890 662850
rect 151980 662610 152220 662850
rect 152310 662610 152550 662850
rect 152640 662610 152880 662850
rect 152990 662610 153230 662850
rect 153320 662610 153560 662850
rect 153650 662610 153890 662850
rect 153980 662610 154220 662850
rect 154330 662610 154570 662850
rect 154660 662610 154900 662850
rect 154990 662610 155230 662850
rect 155320 662610 155560 662850
rect 155670 662610 155910 662850
rect 144950 662280 145190 662520
rect 145280 662280 145520 662520
rect 145610 662280 145850 662520
rect 145940 662280 146180 662520
rect 146290 662280 146530 662520
rect 146620 662280 146860 662520
rect 146950 662280 147190 662520
rect 147280 662280 147520 662520
rect 147630 662280 147870 662520
rect 147960 662280 148200 662520
rect 148290 662280 148530 662520
rect 148620 662280 148860 662520
rect 148970 662280 149210 662520
rect 149300 662280 149540 662520
rect 149630 662280 149870 662520
rect 149960 662280 150200 662520
rect 150310 662280 150550 662520
rect 150640 662280 150880 662520
rect 150970 662280 151210 662520
rect 151300 662280 151540 662520
rect 151650 662280 151890 662520
rect 151980 662280 152220 662520
rect 152310 662280 152550 662520
rect 152640 662280 152880 662520
rect 152990 662280 153230 662520
rect 153320 662280 153560 662520
rect 153650 662280 153890 662520
rect 153980 662280 154220 662520
rect 154330 662280 154570 662520
rect 154660 662280 154900 662520
rect 154990 662280 155230 662520
rect 155320 662280 155560 662520
rect 155670 662280 155910 662520
rect 144950 661930 145190 662170
rect 145280 661930 145520 662170
rect 145610 661930 145850 662170
rect 145940 661930 146180 662170
rect 146290 661930 146530 662170
rect 146620 661930 146860 662170
rect 146950 661930 147190 662170
rect 147280 661930 147520 662170
rect 147630 661930 147870 662170
rect 147960 661930 148200 662170
rect 148290 661930 148530 662170
rect 148620 661930 148860 662170
rect 148970 661930 149210 662170
rect 149300 661930 149540 662170
rect 149630 661930 149870 662170
rect 149960 661930 150200 662170
rect 150310 661930 150550 662170
rect 150640 661930 150880 662170
rect 150970 661930 151210 662170
rect 151300 661930 151540 662170
rect 151650 661930 151890 662170
rect 151980 661930 152220 662170
rect 152310 661930 152550 662170
rect 152640 661930 152880 662170
rect 152990 661930 153230 662170
rect 153320 661930 153560 662170
rect 153650 661930 153890 662170
rect 153980 661930 154220 662170
rect 154330 661930 154570 662170
rect 154660 661930 154900 662170
rect 154990 661930 155230 662170
rect 155320 661930 155560 662170
rect 155670 661930 155910 662170
rect 144950 661600 145190 661840
rect 145280 661600 145520 661840
rect 145610 661600 145850 661840
rect 145940 661600 146180 661840
rect 146290 661600 146530 661840
rect 146620 661600 146860 661840
rect 146950 661600 147190 661840
rect 147280 661600 147520 661840
rect 147630 661600 147870 661840
rect 147960 661600 148200 661840
rect 148290 661600 148530 661840
rect 148620 661600 148860 661840
rect 148970 661600 149210 661840
rect 149300 661600 149540 661840
rect 149630 661600 149870 661840
rect 149960 661600 150200 661840
rect 150310 661600 150550 661840
rect 150640 661600 150880 661840
rect 150970 661600 151210 661840
rect 151300 661600 151540 661840
rect 151650 661600 151890 661840
rect 151980 661600 152220 661840
rect 152310 661600 152550 661840
rect 152640 661600 152880 661840
rect 152990 661600 153230 661840
rect 153320 661600 153560 661840
rect 153650 661600 153890 661840
rect 153980 661600 154220 661840
rect 154330 661600 154570 661840
rect 154660 661600 154900 661840
rect 154990 661600 155230 661840
rect 155320 661600 155560 661840
rect 155670 661600 155910 661840
rect 144950 661270 145190 661510
rect 145280 661270 145520 661510
rect 145610 661270 145850 661510
rect 145940 661270 146180 661510
rect 146290 661270 146530 661510
rect 146620 661270 146860 661510
rect 146950 661270 147190 661510
rect 147280 661270 147520 661510
rect 147630 661270 147870 661510
rect 147960 661270 148200 661510
rect 148290 661270 148530 661510
rect 148620 661270 148860 661510
rect 148970 661270 149210 661510
rect 149300 661270 149540 661510
rect 149630 661270 149870 661510
rect 149960 661270 150200 661510
rect 150310 661270 150550 661510
rect 150640 661270 150880 661510
rect 150970 661270 151210 661510
rect 151300 661270 151540 661510
rect 151650 661270 151890 661510
rect 151980 661270 152220 661510
rect 152310 661270 152550 661510
rect 152640 661270 152880 661510
rect 152990 661270 153230 661510
rect 153320 661270 153560 661510
rect 153650 661270 153890 661510
rect 153980 661270 154220 661510
rect 154330 661270 154570 661510
rect 154660 661270 154900 661510
rect 154990 661270 155230 661510
rect 155320 661270 155560 661510
rect 155670 661270 155910 661510
rect 144950 660940 145190 661180
rect 145280 660940 145520 661180
rect 145610 660940 145850 661180
rect 145940 660940 146180 661180
rect 146290 660940 146530 661180
rect 146620 660940 146860 661180
rect 146950 660940 147190 661180
rect 147280 660940 147520 661180
rect 147630 660940 147870 661180
rect 147960 660940 148200 661180
rect 148290 660940 148530 661180
rect 148620 660940 148860 661180
rect 148970 660940 149210 661180
rect 149300 660940 149540 661180
rect 149630 660940 149870 661180
rect 149960 660940 150200 661180
rect 150310 660940 150550 661180
rect 150640 660940 150880 661180
rect 150970 660940 151210 661180
rect 151300 660940 151540 661180
rect 151650 660940 151890 661180
rect 151980 660940 152220 661180
rect 152310 660940 152550 661180
rect 152640 660940 152880 661180
rect 152990 660940 153230 661180
rect 153320 660940 153560 661180
rect 153650 660940 153890 661180
rect 153980 660940 154220 661180
rect 154330 660940 154570 661180
rect 154660 660940 154900 661180
rect 154990 660940 155230 661180
rect 155320 660940 155560 661180
rect 155670 660940 155910 661180
rect 110810 660100 111050 660340
rect 111160 660100 111400 660340
rect 111490 660100 111730 660340
rect 111820 660100 112060 660340
rect 112150 660100 112390 660340
rect 112500 660100 112740 660340
rect 112830 660100 113070 660340
rect 113160 660100 113400 660340
rect 113490 660100 113730 660340
rect 113840 660100 114080 660340
rect 114170 660100 114410 660340
rect 114500 660100 114740 660340
rect 114830 660100 115070 660340
rect 115180 660100 115420 660340
rect 115510 660100 115750 660340
rect 115840 660100 116080 660340
rect 116170 660100 116410 660340
rect 116520 660100 116760 660340
rect 116850 660100 117090 660340
rect 117180 660100 117420 660340
rect 117510 660100 117750 660340
rect 117860 660100 118100 660340
rect 118190 660100 118430 660340
rect 118520 660100 118760 660340
rect 118850 660100 119090 660340
rect 119200 660100 119440 660340
rect 119530 660100 119770 660340
rect 119860 660100 120100 660340
rect 120190 660100 120430 660340
rect 120540 660100 120780 660340
rect 120870 660100 121110 660340
rect 121200 660100 121440 660340
rect 121530 660100 121770 660340
rect 110810 659770 111050 660010
rect 111160 659770 111400 660010
rect 111490 659770 111730 660010
rect 111820 659770 112060 660010
rect 112150 659770 112390 660010
rect 112500 659770 112740 660010
rect 112830 659770 113070 660010
rect 113160 659770 113400 660010
rect 113490 659770 113730 660010
rect 113840 659770 114080 660010
rect 114170 659770 114410 660010
rect 114500 659770 114740 660010
rect 114830 659770 115070 660010
rect 115180 659770 115420 660010
rect 115510 659770 115750 660010
rect 115840 659770 116080 660010
rect 116170 659770 116410 660010
rect 116520 659770 116760 660010
rect 116850 659770 117090 660010
rect 117180 659770 117420 660010
rect 117510 659770 117750 660010
rect 117860 659770 118100 660010
rect 118190 659770 118430 660010
rect 118520 659770 118760 660010
rect 118850 659770 119090 660010
rect 119200 659770 119440 660010
rect 119530 659770 119770 660010
rect 119860 659770 120100 660010
rect 120190 659770 120430 660010
rect 120540 659770 120780 660010
rect 120870 659770 121110 660010
rect 121200 659770 121440 660010
rect 121530 659770 121770 660010
rect 110810 659440 111050 659680
rect 111160 659440 111400 659680
rect 111490 659440 111730 659680
rect 111820 659440 112060 659680
rect 112150 659440 112390 659680
rect 112500 659440 112740 659680
rect 112830 659440 113070 659680
rect 113160 659440 113400 659680
rect 113490 659440 113730 659680
rect 113840 659440 114080 659680
rect 114170 659440 114410 659680
rect 114500 659440 114740 659680
rect 114830 659440 115070 659680
rect 115180 659440 115420 659680
rect 115510 659440 115750 659680
rect 115840 659440 116080 659680
rect 116170 659440 116410 659680
rect 116520 659440 116760 659680
rect 116850 659440 117090 659680
rect 117180 659440 117420 659680
rect 117510 659440 117750 659680
rect 117860 659440 118100 659680
rect 118190 659440 118430 659680
rect 118520 659440 118760 659680
rect 118850 659440 119090 659680
rect 119200 659440 119440 659680
rect 119530 659440 119770 659680
rect 119860 659440 120100 659680
rect 120190 659440 120430 659680
rect 120540 659440 120780 659680
rect 120870 659440 121110 659680
rect 121200 659440 121440 659680
rect 121530 659440 121770 659680
rect 110810 659110 111050 659350
rect 111160 659110 111400 659350
rect 111490 659110 111730 659350
rect 111820 659110 112060 659350
rect 112150 659110 112390 659350
rect 112500 659110 112740 659350
rect 112830 659110 113070 659350
rect 113160 659110 113400 659350
rect 113490 659110 113730 659350
rect 113840 659110 114080 659350
rect 114170 659110 114410 659350
rect 114500 659110 114740 659350
rect 114830 659110 115070 659350
rect 115180 659110 115420 659350
rect 115510 659110 115750 659350
rect 115840 659110 116080 659350
rect 116170 659110 116410 659350
rect 116520 659110 116760 659350
rect 116850 659110 117090 659350
rect 117180 659110 117420 659350
rect 117510 659110 117750 659350
rect 117860 659110 118100 659350
rect 118190 659110 118430 659350
rect 118520 659110 118760 659350
rect 118850 659110 119090 659350
rect 119200 659110 119440 659350
rect 119530 659110 119770 659350
rect 119860 659110 120100 659350
rect 120190 659110 120430 659350
rect 120540 659110 120780 659350
rect 120870 659110 121110 659350
rect 121200 659110 121440 659350
rect 121530 659110 121770 659350
rect 110810 658760 111050 659000
rect 111160 658760 111400 659000
rect 111490 658760 111730 659000
rect 111820 658760 112060 659000
rect 112150 658760 112390 659000
rect 112500 658760 112740 659000
rect 112830 658760 113070 659000
rect 113160 658760 113400 659000
rect 113490 658760 113730 659000
rect 113840 658760 114080 659000
rect 114170 658760 114410 659000
rect 114500 658760 114740 659000
rect 114830 658760 115070 659000
rect 115180 658760 115420 659000
rect 115510 658760 115750 659000
rect 115840 658760 116080 659000
rect 116170 658760 116410 659000
rect 116520 658760 116760 659000
rect 116850 658760 117090 659000
rect 117180 658760 117420 659000
rect 117510 658760 117750 659000
rect 117860 658760 118100 659000
rect 118190 658760 118430 659000
rect 118520 658760 118760 659000
rect 118850 658760 119090 659000
rect 119200 658760 119440 659000
rect 119530 658760 119770 659000
rect 119860 658760 120100 659000
rect 120190 658760 120430 659000
rect 120540 658760 120780 659000
rect 120870 658760 121110 659000
rect 121200 658760 121440 659000
rect 121530 658760 121770 659000
rect 110810 658430 111050 658670
rect 111160 658430 111400 658670
rect 111490 658430 111730 658670
rect 111820 658430 112060 658670
rect 112150 658430 112390 658670
rect 112500 658430 112740 658670
rect 112830 658430 113070 658670
rect 113160 658430 113400 658670
rect 113490 658430 113730 658670
rect 113840 658430 114080 658670
rect 114170 658430 114410 658670
rect 114500 658430 114740 658670
rect 114830 658430 115070 658670
rect 115180 658430 115420 658670
rect 115510 658430 115750 658670
rect 115840 658430 116080 658670
rect 116170 658430 116410 658670
rect 116520 658430 116760 658670
rect 116850 658430 117090 658670
rect 117180 658430 117420 658670
rect 117510 658430 117750 658670
rect 117860 658430 118100 658670
rect 118190 658430 118430 658670
rect 118520 658430 118760 658670
rect 118850 658430 119090 658670
rect 119200 658430 119440 658670
rect 119530 658430 119770 658670
rect 119860 658430 120100 658670
rect 120190 658430 120430 658670
rect 120540 658430 120780 658670
rect 120870 658430 121110 658670
rect 121200 658430 121440 658670
rect 121530 658430 121770 658670
rect 110810 658100 111050 658340
rect 111160 658100 111400 658340
rect 111490 658100 111730 658340
rect 111820 658100 112060 658340
rect 112150 658100 112390 658340
rect 112500 658100 112740 658340
rect 112830 658100 113070 658340
rect 113160 658100 113400 658340
rect 113490 658100 113730 658340
rect 113840 658100 114080 658340
rect 114170 658100 114410 658340
rect 114500 658100 114740 658340
rect 114830 658100 115070 658340
rect 115180 658100 115420 658340
rect 115510 658100 115750 658340
rect 115840 658100 116080 658340
rect 116170 658100 116410 658340
rect 116520 658100 116760 658340
rect 116850 658100 117090 658340
rect 117180 658100 117420 658340
rect 117510 658100 117750 658340
rect 117860 658100 118100 658340
rect 118190 658100 118430 658340
rect 118520 658100 118760 658340
rect 118850 658100 119090 658340
rect 119200 658100 119440 658340
rect 119530 658100 119770 658340
rect 119860 658100 120100 658340
rect 120190 658100 120430 658340
rect 120540 658100 120780 658340
rect 120870 658100 121110 658340
rect 121200 658100 121440 658340
rect 121530 658100 121770 658340
rect 110810 657770 111050 658010
rect 111160 657770 111400 658010
rect 111490 657770 111730 658010
rect 111820 657770 112060 658010
rect 112150 657770 112390 658010
rect 112500 657770 112740 658010
rect 112830 657770 113070 658010
rect 113160 657770 113400 658010
rect 113490 657770 113730 658010
rect 113840 657770 114080 658010
rect 114170 657770 114410 658010
rect 114500 657770 114740 658010
rect 114830 657770 115070 658010
rect 115180 657770 115420 658010
rect 115510 657770 115750 658010
rect 115840 657770 116080 658010
rect 116170 657770 116410 658010
rect 116520 657770 116760 658010
rect 116850 657770 117090 658010
rect 117180 657770 117420 658010
rect 117510 657770 117750 658010
rect 117860 657770 118100 658010
rect 118190 657770 118430 658010
rect 118520 657770 118760 658010
rect 118850 657770 119090 658010
rect 119200 657770 119440 658010
rect 119530 657770 119770 658010
rect 119860 657770 120100 658010
rect 120190 657770 120430 658010
rect 120540 657770 120780 658010
rect 120870 657770 121110 658010
rect 121200 657770 121440 658010
rect 121530 657770 121770 658010
rect 110810 657420 111050 657660
rect 111160 657420 111400 657660
rect 111490 657420 111730 657660
rect 111820 657420 112060 657660
rect 112150 657420 112390 657660
rect 112500 657420 112740 657660
rect 112830 657420 113070 657660
rect 113160 657420 113400 657660
rect 113490 657420 113730 657660
rect 113840 657420 114080 657660
rect 114170 657420 114410 657660
rect 114500 657420 114740 657660
rect 114830 657420 115070 657660
rect 115180 657420 115420 657660
rect 115510 657420 115750 657660
rect 115840 657420 116080 657660
rect 116170 657420 116410 657660
rect 116520 657420 116760 657660
rect 116850 657420 117090 657660
rect 117180 657420 117420 657660
rect 117510 657420 117750 657660
rect 117860 657420 118100 657660
rect 118190 657420 118430 657660
rect 118520 657420 118760 657660
rect 118850 657420 119090 657660
rect 119200 657420 119440 657660
rect 119530 657420 119770 657660
rect 119860 657420 120100 657660
rect 120190 657420 120430 657660
rect 120540 657420 120780 657660
rect 120870 657420 121110 657660
rect 121200 657420 121440 657660
rect 121530 657420 121770 657660
rect 110810 657090 111050 657330
rect 111160 657090 111400 657330
rect 111490 657090 111730 657330
rect 111820 657090 112060 657330
rect 112150 657090 112390 657330
rect 112500 657090 112740 657330
rect 112830 657090 113070 657330
rect 113160 657090 113400 657330
rect 113490 657090 113730 657330
rect 113840 657090 114080 657330
rect 114170 657090 114410 657330
rect 114500 657090 114740 657330
rect 114830 657090 115070 657330
rect 115180 657090 115420 657330
rect 115510 657090 115750 657330
rect 115840 657090 116080 657330
rect 116170 657090 116410 657330
rect 116520 657090 116760 657330
rect 116850 657090 117090 657330
rect 117180 657090 117420 657330
rect 117510 657090 117750 657330
rect 117860 657090 118100 657330
rect 118190 657090 118430 657330
rect 118520 657090 118760 657330
rect 118850 657090 119090 657330
rect 119200 657090 119440 657330
rect 119530 657090 119770 657330
rect 119860 657090 120100 657330
rect 120190 657090 120430 657330
rect 120540 657090 120780 657330
rect 120870 657090 121110 657330
rect 121200 657090 121440 657330
rect 121530 657090 121770 657330
rect 110810 656760 111050 657000
rect 111160 656760 111400 657000
rect 111490 656760 111730 657000
rect 111820 656760 112060 657000
rect 112150 656760 112390 657000
rect 112500 656760 112740 657000
rect 112830 656760 113070 657000
rect 113160 656760 113400 657000
rect 113490 656760 113730 657000
rect 113840 656760 114080 657000
rect 114170 656760 114410 657000
rect 114500 656760 114740 657000
rect 114830 656760 115070 657000
rect 115180 656760 115420 657000
rect 115510 656760 115750 657000
rect 115840 656760 116080 657000
rect 116170 656760 116410 657000
rect 116520 656760 116760 657000
rect 116850 656760 117090 657000
rect 117180 656760 117420 657000
rect 117510 656760 117750 657000
rect 117860 656760 118100 657000
rect 118190 656760 118430 657000
rect 118520 656760 118760 657000
rect 118850 656760 119090 657000
rect 119200 656760 119440 657000
rect 119530 656760 119770 657000
rect 119860 656760 120100 657000
rect 120190 656760 120430 657000
rect 120540 656760 120780 657000
rect 120870 656760 121110 657000
rect 121200 656760 121440 657000
rect 121530 656760 121770 657000
rect 110810 656430 111050 656670
rect 111160 656430 111400 656670
rect 111490 656430 111730 656670
rect 111820 656430 112060 656670
rect 112150 656430 112390 656670
rect 112500 656430 112740 656670
rect 112830 656430 113070 656670
rect 113160 656430 113400 656670
rect 113490 656430 113730 656670
rect 113840 656430 114080 656670
rect 114170 656430 114410 656670
rect 114500 656430 114740 656670
rect 114830 656430 115070 656670
rect 115180 656430 115420 656670
rect 115510 656430 115750 656670
rect 115840 656430 116080 656670
rect 116170 656430 116410 656670
rect 116520 656430 116760 656670
rect 116850 656430 117090 656670
rect 117180 656430 117420 656670
rect 117510 656430 117750 656670
rect 117860 656430 118100 656670
rect 118190 656430 118430 656670
rect 118520 656430 118760 656670
rect 118850 656430 119090 656670
rect 119200 656430 119440 656670
rect 119530 656430 119770 656670
rect 119860 656430 120100 656670
rect 120190 656430 120430 656670
rect 120540 656430 120780 656670
rect 120870 656430 121110 656670
rect 121200 656430 121440 656670
rect 121530 656430 121770 656670
rect 110810 656080 111050 656320
rect 111160 656080 111400 656320
rect 111490 656080 111730 656320
rect 111820 656080 112060 656320
rect 112150 656080 112390 656320
rect 112500 656080 112740 656320
rect 112830 656080 113070 656320
rect 113160 656080 113400 656320
rect 113490 656080 113730 656320
rect 113840 656080 114080 656320
rect 114170 656080 114410 656320
rect 114500 656080 114740 656320
rect 114830 656080 115070 656320
rect 115180 656080 115420 656320
rect 115510 656080 115750 656320
rect 115840 656080 116080 656320
rect 116170 656080 116410 656320
rect 116520 656080 116760 656320
rect 116850 656080 117090 656320
rect 117180 656080 117420 656320
rect 117510 656080 117750 656320
rect 117860 656080 118100 656320
rect 118190 656080 118430 656320
rect 118520 656080 118760 656320
rect 118850 656080 119090 656320
rect 119200 656080 119440 656320
rect 119530 656080 119770 656320
rect 119860 656080 120100 656320
rect 120190 656080 120430 656320
rect 120540 656080 120780 656320
rect 120870 656080 121110 656320
rect 121200 656080 121440 656320
rect 121530 656080 121770 656320
rect 110810 655750 111050 655990
rect 111160 655750 111400 655990
rect 111490 655750 111730 655990
rect 111820 655750 112060 655990
rect 112150 655750 112390 655990
rect 112500 655750 112740 655990
rect 112830 655750 113070 655990
rect 113160 655750 113400 655990
rect 113490 655750 113730 655990
rect 113840 655750 114080 655990
rect 114170 655750 114410 655990
rect 114500 655750 114740 655990
rect 114830 655750 115070 655990
rect 115180 655750 115420 655990
rect 115510 655750 115750 655990
rect 115840 655750 116080 655990
rect 116170 655750 116410 655990
rect 116520 655750 116760 655990
rect 116850 655750 117090 655990
rect 117180 655750 117420 655990
rect 117510 655750 117750 655990
rect 117860 655750 118100 655990
rect 118190 655750 118430 655990
rect 118520 655750 118760 655990
rect 118850 655750 119090 655990
rect 119200 655750 119440 655990
rect 119530 655750 119770 655990
rect 119860 655750 120100 655990
rect 120190 655750 120430 655990
rect 120540 655750 120780 655990
rect 120870 655750 121110 655990
rect 121200 655750 121440 655990
rect 121530 655750 121770 655990
rect 110810 655420 111050 655660
rect 111160 655420 111400 655660
rect 111490 655420 111730 655660
rect 111820 655420 112060 655660
rect 112150 655420 112390 655660
rect 112500 655420 112740 655660
rect 112830 655420 113070 655660
rect 113160 655420 113400 655660
rect 113490 655420 113730 655660
rect 113840 655420 114080 655660
rect 114170 655420 114410 655660
rect 114500 655420 114740 655660
rect 114830 655420 115070 655660
rect 115180 655420 115420 655660
rect 115510 655420 115750 655660
rect 115840 655420 116080 655660
rect 116170 655420 116410 655660
rect 116520 655420 116760 655660
rect 116850 655420 117090 655660
rect 117180 655420 117420 655660
rect 117510 655420 117750 655660
rect 117860 655420 118100 655660
rect 118190 655420 118430 655660
rect 118520 655420 118760 655660
rect 118850 655420 119090 655660
rect 119200 655420 119440 655660
rect 119530 655420 119770 655660
rect 119860 655420 120100 655660
rect 120190 655420 120430 655660
rect 120540 655420 120780 655660
rect 120870 655420 121110 655660
rect 121200 655420 121440 655660
rect 121530 655420 121770 655660
rect 110810 655090 111050 655330
rect 111160 655090 111400 655330
rect 111490 655090 111730 655330
rect 111820 655090 112060 655330
rect 112150 655090 112390 655330
rect 112500 655090 112740 655330
rect 112830 655090 113070 655330
rect 113160 655090 113400 655330
rect 113490 655090 113730 655330
rect 113840 655090 114080 655330
rect 114170 655090 114410 655330
rect 114500 655090 114740 655330
rect 114830 655090 115070 655330
rect 115180 655090 115420 655330
rect 115510 655090 115750 655330
rect 115840 655090 116080 655330
rect 116170 655090 116410 655330
rect 116520 655090 116760 655330
rect 116850 655090 117090 655330
rect 117180 655090 117420 655330
rect 117510 655090 117750 655330
rect 117860 655090 118100 655330
rect 118190 655090 118430 655330
rect 118520 655090 118760 655330
rect 118850 655090 119090 655330
rect 119200 655090 119440 655330
rect 119530 655090 119770 655330
rect 119860 655090 120100 655330
rect 120190 655090 120430 655330
rect 120540 655090 120780 655330
rect 120870 655090 121110 655330
rect 121200 655090 121440 655330
rect 121530 655090 121770 655330
rect 110810 654740 111050 654980
rect 111160 654740 111400 654980
rect 111490 654740 111730 654980
rect 111820 654740 112060 654980
rect 112150 654740 112390 654980
rect 112500 654740 112740 654980
rect 112830 654740 113070 654980
rect 113160 654740 113400 654980
rect 113490 654740 113730 654980
rect 113840 654740 114080 654980
rect 114170 654740 114410 654980
rect 114500 654740 114740 654980
rect 114830 654740 115070 654980
rect 115180 654740 115420 654980
rect 115510 654740 115750 654980
rect 115840 654740 116080 654980
rect 116170 654740 116410 654980
rect 116520 654740 116760 654980
rect 116850 654740 117090 654980
rect 117180 654740 117420 654980
rect 117510 654740 117750 654980
rect 117860 654740 118100 654980
rect 118190 654740 118430 654980
rect 118520 654740 118760 654980
rect 118850 654740 119090 654980
rect 119200 654740 119440 654980
rect 119530 654740 119770 654980
rect 119860 654740 120100 654980
rect 120190 654740 120430 654980
rect 120540 654740 120780 654980
rect 120870 654740 121110 654980
rect 121200 654740 121440 654980
rect 121530 654740 121770 654980
rect 110810 654410 111050 654650
rect 111160 654410 111400 654650
rect 111490 654410 111730 654650
rect 111820 654410 112060 654650
rect 112150 654410 112390 654650
rect 112500 654410 112740 654650
rect 112830 654410 113070 654650
rect 113160 654410 113400 654650
rect 113490 654410 113730 654650
rect 113840 654410 114080 654650
rect 114170 654410 114410 654650
rect 114500 654410 114740 654650
rect 114830 654410 115070 654650
rect 115180 654410 115420 654650
rect 115510 654410 115750 654650
rect 115840 654410 116080 654650
rect 116170 654410 116410 654650
rect 116520 654410 116760 654650
rect 116850 654410 117090 654650
rect 117180 654410 117420 654650
rect 117510 654410 117750 654650
rect 117860 654410 118100 654650
rect 118190 654410 118430 654650
rect 118520 654410 118760 654650
rect 118850 654410 119090 654650
rect 119200 654410 119440 654650
rect 119530 654410 119770 654650
rect 119860 654410 120100 654650
rect 120190 654410 120430 654650
rect 120540 654410 120780 654650
rect 120870 654410 121110 654650
rect 121200 654410 121440 654650
rect 121530 654410 121770 654650
rect 110810 654080 111050 654320
rect 111160 654080 111400 654320
rect 111490 654080 111730 654320
rect 111820 654080 112060 654320
rect 112150 654080 112390 654320
rect 112500 654080 112740 654320
rect 112830 654080 113070 654320
rect 113160 654080 113400 654320
rect 113490 654080 113730 654320
rect 113840 654080 114080 654320
rect 114170 654080 114410 654320
rect 114500 654080 114740 654320
rect 114830 654080 115070 654320
rect 115180 654080 115420 654320
rect 115510 654080 115750 654320
rect 115840 654080 116080 654320
rect 116170 654080 116410 654320
rect 116520 654080 116760 654320
rect 116850 654080 117090 654320
rect 117180 654080 117420 654320
rect 117510 654080 117750 654320
rect 117860 654080 118100 654320
rect 118190 654080 118430 654320
rect 118520 654080 118760 654320
rect 118850 654080 119090 654320
rect 119200 654080 119440 654320
rect 119530 654080 119770 654320
rect 119860 654080 120100 654320
rect 120190 654080 120430 654320
rect 120540 654080 120780 654320
rect 120870 654080 121110 654320
rect 121200 654080 121440 654320
rect 121530 654080 121770 654320
rect 110810 653750 111050 653990
rect 111160 653750 111400 653990
rect 111490 653750 111730 653990
rect 111820 653750 112060 653990
rect 112150 653750 112390 653990
rect 112500 653750 112740 653990
rect 112830 653750 113070 653990
rect 113160 653750 113400 653990
rect 113490 653750 113730 653990
rect 113840 653750 114080 653990
rect 114170 653750 114410 653990
rect 114500 653750 114740 653990
rect 114830 653750 115070 653990
rect 115180 653750 115420 653990
rect 115510 653750 115750 653990
rect 115840 653750 116080 653990
rect 116170 653750 116410 653990
rect 116520 653750 116760 653990
rect 116850 653750 117090 653990
rect 117180 653750 117420 653990
rect 117510 653750 117750 653990
rect 117860 653750 118100 653990
rect 118190 653750 118430 653990
rect 118520 653750 118760 653990
rect 118850 653750 119090 653990
rect 119200 653750 119440 653990
rect 119530 653750 119770 653990
rect 119860 653750 120100 653990
rect 120190 653750 120430 653990
rect 120540 653750 120780 653990
rect 120870 653750 121110 653990
rect 121200 653750 121440 653990
rect 121530 653750 121770 653990
rect 110810 653400 111050 653640
rect 111160 653400 111400 653640
rect 111490 653400 111730 653640
rect 111820 653400 112060 653640
rect 112150 653400 112390 653640
rect 112500 653400 112740 653640
rect 112830 653400 113070 653640
rect 113160 653400 113400 653640
rect 113490 653400 113730 653640
rect 113840 653400 114080 653640
rect 114170 653400 114410 653640
rect 114500 653400 114740 653640
rect 114830 653400 115070 653640
rect 115180 653400 115420 653640
rect 115510 653400 115750 653640
rect 115840 653400 116080 653640
rect 116170 653400 116410 653640
rect 116520 653400 116760 653640
rect 116850 653400 117090 653640
rect 117180 653400 117420 653640
rect 117510 653400 117750 653640
rect 117860 653400 118100 653640
rect 118190 653400 118430 653640
rect 118520 653400 118760 653640
rect 118850 653400 119090 653640
rect 119200 653400 119440 653640
rect 119530 653400 119770 653640
rect 119860 653400 120100 653640
rect 120190 653400 120430 653640
rect 120540 653400 120780 653640
rect 120870 653400 121110 653640
rect 121200 653400 121440 653640
rect 121530 653400 121770 653640
rect 110810 653070 111050 653310
rect 111160 653070 111400 653310
rect 111490 653070 111730 653310
rect 111820 653070 112060 653310
rect 112150 653070 112390 653310
rect 112500 653070 112740 653310
rect 112830 653070 113070 653310
rect 113160 653070 113400 653310
rect 113490 653070 113730 653310
rect 113840 653070 114080 653310
rect 114170 653070 114410 653310
rect 114500 653070 114740 653310
rect 114830 653070 115070 653310
rect 115180 653070 115420 653310
rect 115510 653070 115750 653310
rect 115840 653070 116080 653310
rect 116170 653070 116410 653310
rect 116520 653070 116760 653310
rect 116850 653070 117090 653310
rect 117180 653070 117420 653310
rect 117510 653070 117750 653310
rect 117860 653070 118100 653310
rect 118190 653070 118430 653310
rect 118520 653070 118760 653310
rect 118850 653070 119090 653310
rect 119200 653070 119440 653310
rect 119530 653070 119770 653310
rect 119860 653070 120100 653310
rect 120190 653070 120430 653310
rect 120540 653070 120780 653310
rect 120870 653070 121110 653310
rect 121200 653070 121440 653310
rect 121530 653070 121770 653310
rect 110810 652740 111050 652980
rect 111160 652740 111400 652980
rect 111490 652740 111730 652980
rect 111820 652740 112060 652980
rect 112150 652740 112390 652980
rect 112500 652740 112740 652980
rect 112830 652740 113070 652980
rect 113160 652740 113400 652980
rect 113490 652740 113730 652980
rect 113840 652740 114080 652980
rect 114170 652740 114410 652980
rect 114500 652740 114740 652980
rect 114830 652740 115070 652980
rect 115180 652740 115420 652980
rect 115510 652740 115750 652980
rect 115840 652740 116080 652980
rect 116170 652740 116410 652980
rect 116520 652740 116760 652980
rect 116850 652740 117090 652980
rect 117180 652740 117420 652980
rect 117510 652740 117750 652980
rect 117860 652740 118100 652980
rect 118190 652740 118430 652980
rect 118520 652740 118760 652980
rect 118850 652740 119090 652980
rect 119200 652740 119440 652980
rect 119530 652740 119770 652980
rect 119860 652740 120100 652980
rect 120190 652740 120430 652980
rect 120540 652740 120780 652980
rect 120870 652740 121110 652980
rect 121200 652740 121440 652980
rect 121530 652740 121770 652980
rect 110810 652410 111050 652650
rect 111160 652410 111400 652650
rect 111490 652410 111730 652650
rect 111820 652410 112060 652650
rect 112150 652410 112390 652650
rect 112500 652410 112740 652650
rect 112830 652410 113070 652650
rect 113160 652410 113400 652650
rect 113490 652410 113730 652650
rect 113840 652410 114080 652650
rect 114170 652410 114410 652650
rect 114500 652410 114740 652650
rect 114830 652410 115070 652650
rect 115180 652410 115420 652650
rect 115510 652410 115750 652650
rect 115840 652410 116080 652650
rect 116170 652410 116410 652650
rect 116520 652410 116760 652650
rect 116850 652410 117090 652650
rect 117180 652410 117420 652650
rect 117510 652410 117750 652650
rect 117860 652410 118100 652650
rect 118190 652410 118430 652650
rect 118520 652410 118760 652650
rect 118850 652410 119090 652650
rect 119200 652410 119440 652650
rect 119530 652410 119770 652650
rect 119860 652410 120100 652650
rect 120190 652410 120430 652650
rect 120540 652410 120780 652650
rect 120870 652410 121110 652650
rect 121200 652410 121440 652650
rect 121530 652410 121770 652650
rect 110810 652060 111050 652300
rect 111160 652060 111400 652300
rect 111490 652060 111730 652300
rect 111820 652060 112060 652300
rect 112150 652060 112390 652300
rect 112500 652060 112740 652300
rect 112830 652060 113070 652300
rect 113160 652060 113400 652300
rect 113490 652060 113730 652300
rect 113840 652060 114080 652300
rect 114170 652060 114410 652300
rect 114500 652060 114740 652300
rect 114830 652060 115070 652300
rect 115180 652060 115420 652300
rect 115510 652060 115750 652300
rect 115840 652060 116080 652300
rect 116170 652060 116410 652300
rect 116520 652060 116760 652300
rect 116850 652060 117090 652300
rect 117180 652060 117420 652300
rect 117510 652060 117750 652300
rect 117860 652060 118100 652300
rect 118190 652060 118430 652300
rect 118520 652060 118760 652300
rect 118850 652060 119090 652300
rect 119200 652060 119440 652300
rect 119530 652060 119770 652300
rect 119860 652060 120100 652300
rect 120190 652060 120430 652300
rect 120540 652060 120780 652300
rect 120870 652060 121110 652300
rect 121200 652060 121440 652300
rect 121530 652060 121770 652300
rect 110810 651730 111050 651970
rect 111160 651730 111400 651970
rect 111490 651730 111730 651970
rect 111820 651730 112060 651970
rect 112150 651730 112390 651970
rect 112500 651730 112740 651970
rect 112830 651730 113070 651970
rect 113160 651730 113400 651970
rect 113490 651730 113730 651970
rect 113840 651730 114080 651970
rect 114170 651730 114410 651970
rect 114500 651730 114740 651970
rect 114830 651730 115070 651970
rect 115180 651730 115420 651970
rect 115510 651730 115750 651970
rect 115840 651730 116080 651970
rect 116170 651730 116410 651970
rect 116520 651730 116760 651970
rect 116850 651730 117090 651970
rect 117180 651730 117420 651970
rect 117510 651730 117750 651970
rect 117860 651730 118100 651970
rect 118190 651730 118430 651970
rect 118520 651730 118760 651970
rect 118850 651730 119090 651970
rect 119200 651730 119440 651970
rect 119530 651730 119770 651970
rect 119860 651730 120100 651970
rect 120190 651730 120430 651970
rect 120540 651730 120780 651970
rect 120870 651730 121110 651970
rect 121200 651730 121440 651970
rect 121530 651730 121770 651970
rect 110810 651400 111050 651640
rect 111160 651400 111400 651640
rect 111490 651400 111730 651640
rect 111820 651400 112060 651640
rect 112150 651400 112390 651640
rect 112500 651400 112740 651640
rect 112830 651400 113070 651640
rect 113160 651400 113400 651640
rect 113490 651400 113730 651640
rect 113840 651400 114080 651640
rect 114170 651400 114410 651640
rect 114500 651400 114740 651640
rect 114830 651400 115070 651640
rect 115180 651400 115420 651640
rect 115510 651400 115750 651640
rect 115840 651400 116080 651640
rect 116170 651400 116410 651640
rect 116520 651400 116760 651640
rect 116850 651400 117090 651640
rect 117180 651400 117420 651640
rect 117510 651400 117750 651640
rect 117860 651400 118100 651640
rect 118190 651400 118430 651640
rect 118520 651400 118760 651640
rect 118850 651400 119090 651640
rect 119200 651400 119440 651640
rect 119530 651400 119770 651640
rect 119860 651400 120100 651640
rect 120190 651400 120430 651640
rect 120540 651400 120780 651640
rect 120870 651400 121110 651640
rect 121200 651400 121440 651640
rect 121530 651400 121770 651640
rect 110810 651070 111050 651310
rect 111160 651070 111400 651310
rect 111490 651070 111730 651310
rect 111820 651070 112060 651310
rect 112150 651070 112390 651310
rect 112500 651070 112740 651310
rect 112830 651070 113070 651310
rect 113160 651070 113400 651310
rect 113490 651070 113730 651310
rect 113840 651070 114080 651310
rect 114170 651070 114410 651310
rect 114500 651070 114740 651310
rect 114830 651070 115070 651310
rect 115180 651070 115420 651310
rect 115510 651070 115750 651310
rect 115840 651070 116080 651310
rect 116170 651070 116410 651310
rect 116520 651070 116760 651310
rect 116850 651070 117090 651310
rect 117180 651070 117420 651310
rect 117510 651070 117750 651310
rect 117860 651070 118100 651310
rect 118190 651070 118430 651310
rect 118520 651070 118760 651310
rect 118850 651070 119090 651310
rect 119200 651070 119440 651310
rect 119530 651070 119770 651310
rect 119860 651070 120100 651310
rect 120190 651070 120430 651310
rect 120540 651070 120780 651310
rect 120870 651070 121110 651310
rect 121200 651070 121440 651310
rect 121530 651070 121770 651310
rect 110810 650720 111050 650960
rect 111160 650720 111400 650960
rect 111490 650720 111730 650960
rect 111820 650720 112060 650960
rect 112150 650720 112390 650960
rect 112500 650720 112740 650960
rect 112830 650720 113070 650960
rect 113160 650720 113400 650960
rect 113490 650720 113730 650960
rect 113840 650720 114080 650960
rect 114170 650720 114410 650960
rect 114500 650720 114740 650960
rect 114830 650720 115070 650960
rect 115180 650720 115420 650960
rect 115510 650720 115750 650960
rect 115840 650720 116080 650960
rect 116170 650720 116410 650960
rect 116520 650720 116760 650960
rect 116850 650720 117090 650960
rect 117180 650720 117420 650960
rect 117510 650720 117750 650960
rect 117860 650720 118100 650960
rect 118190 650720 118430 650960
rect 118520 650720 118760 650960
rect 118850 650720 119090 650960
rect 119200 650720 119440 650960
rect 119530 650720 119770 650960
rect 119860 650720 120100 650960
rect 120190 650720 120430 650960
rect 120540 650720 120780 650960
rect 120870 650720 121110 650960
rect 121200 650720 121440 650960
rect 121530 650720 121770 650960
rect 110810 650390 111050 650630
rect 111160 650390 111400 650630
rect 111490 650390 111730 650630
rect 111820 650390 112060 650630
rect 112150 650390 112390 650630
rect 112500 650390 112740 650630
rect 112830 650390 113070 650630
rect 113160 650390 113400 650630
rect 113490 650390 113730 650630
rect 113840 650390 114080 650630
rect 114170 650390 114410 650630
rect 114500 650390 114740 650630
rect 114830 650390 115070 650630
rect 115180 650390 115420 650630
rect 115510 650390 115750 650630
rect 115840 650390 116080 650630
rect 116170 650390 116410 650630
rect 116520 650390 116760 650630
rect 116850 650390 117090 650630
rect 117180 650390 117420 650630
rect 117510 650390 117750 650630
rect 117860 650390 118100 650630
rect 118190 650390 118430 650630
rect 118520 650390 118760 650630
rect 118850 650390 119090 650630
rect 119200 650390 119440 650630
rect 119530 650390 119770 650630
rect 119860 650390 120100 650630
rect 120190 650390 120430 650630
rect 120540 650390 120780 650630
rect 120870 650390 121110 650630
rect 121200 650390 121440 650630
rect 121530 650390 121770 650630
rect 110810 650060 111050 650300
rect 111160 650060 111400 650300
rect 111490 650060 111730 650300
rect 111820 650060 112060 650300
rect 112150 650060 112390 650300
rect 112500 650060 112740 650300
rect 112830 650060 113070 650300
rect 113160 650060 113400 650300
rect 113490 650060 113730 650300
rect 113840 650060 114080 650300
rect 114170 650060 114410 650300
rect 114500 650060 114740 650300
rect 114830 650060 115070 650300
rect 115180 650060 115420 650300
rect 115510 650060 115750 650300
rect 115840 650060 116080 650300
rect 116170 650060 116410 650300
rect 116520 650060 116760 650300
rect 116850 650060 117090 650300
rect 117180 650060 117420 650300
rect 117510 650060 117750 650300
rect 117860 650060 118100 650300
rect 118190 650060 118430 650300
rect 118520 650060 118760 650300
rect 118850 650060 119090 650300
rect 119200 650060 119440 650300
rect 119530 650060 119770 650300
rect 119860 650060 120100 650300
rect 120190 650060 120430 650300
rect 120540 650060 120780 650300
rect 120870 650060 121110 650300
rect 121200 650060 121440 650300
rect 121530 650060 121770 650300
rect 110810 649730 111050 649970
rect 111160 649730 111400 649970
rect 111490 649730 111730 649970
rect 111820 649730 112060 649970
rect 112150 649730 112390 649970
rect 112500 649730 112740 649970
rect 112830 649730 113070 649970
rect 113160 649730 113400 649970
rect 113490 649730 113730 649970
rect 113840 649730 114080 649970
rect 114170 649730 114410 649970
rect 114500 649730 114740 649970
rect 114830 649730 115070 649970
rect 115180 649730 115420 649970
rect 115510 649730 115750 649970
rect 115840 649730 116080 649970
rect 116170 649730 116410 649970
rect 116520 649730 116760 649970
rect 116850 649730 117090 649970
rect 117180 649730 117420 649970
rect 117510 649730 117750 649970
rect 117860 649730 118100 649970
rect 118190 649730 118430 649970
rect 118520 649730 118760 649970
rect 118850 649730 119090 649970
rect 119200 649730 119440 649970
rect 119530 649730 119770 649970
rect 119860 649730 120100 649970
rect 120190 649730 120430 649970
rect 120540 649730 120780 649970
rect 120870 649730 121110 649970
rect 121200 649730 121440 649970
rect 121530 649730 121770 649970
rect 110810 649380 111050 649620
rect 111160 649380 111400 649620
rect 111490 649380 111730 649620
rect 111820 649380 112060 649620
rect 112150 649380 112390 649620
rect 112500 649380 112740 649620
rect 112830 649380 113070 649620
rect 113160 649380 113400 649620
rect 113490 649380 113730 649620
rect 113840 649380 114080 649620
rect 114170 649380 114410 649620
rect 114500 649380 114740 649620
rect 114830 649380 115070 649620
rect 115180 649380 115420 649620
rect 115510 649380 115750 649620
rect 115840 649380 116080 649620
rect 116170 649380 116410 649620
rect 116520 649380 116760 649620
rect 116850 649380 117090 649620
rect 117180 649380 117420 649620
rect 117510 649380 117750 649620
rect 117860 649380 118100 649620
rect 118190 649380 118430 649620
rect 118520 649380 118760 649620
rect 118850 649380 119090 649620
rect 119200 649380 119440 649620
rect 119530 649380 119770 649620
rect 119860 649380 120100 649620
rect 120190 649380 120430 649620
rect 120540 649380 120780 649620
rect 120870 649380 121110 649620
rect 121200 649380 121440 649620
rect 121530 649380 121770 649620
rect 122190 660100 122430 660340
rect 122540 660100 122780 660340
rect 122870 660100 123110 660340
rect 123200 660100 123440 660340
rect 123530 660100 123770 660340
rect 123880 660100 124120 660340
rect 124210 660100 124450 660340
rect 124540 660100 124780 660340
rect 124870 660100 125110 660340
rect 125220 660100 125460 660340
rect 125550 660100 125790 660340
rect 125880 660100 126120 660340
rect 126210 660100 126450 660340
rect 126560 660100 126800 660340
rect 126890 660100 127130 660340
rect 127220 660100 127460 660340
rect 127550 660100 127790 660340
rect 127900 660100 128140 660340
rect 128230 660100 128470 660340
rect 128560 660100 128800 660340
rect 128890 660100 129130 660340
rect 129240 660100 129480 660340
rect 129570 660100 129810 660340
rect 129900 660100 130140 660340
rect 130230 660100 130470 660340
rect 130580 660100 130820 660340
rect 130910 660100 131150 660340
rect 131240 660100 131480 660340
rect 131570 660100 131810 660340
rect 131920 660100 132160 660340
rect 132250 660100 132490 660340
rect 132580 660100 132820 660340
rect 132910 660100 133150 660340
rect 122190 659770 122430 660010
rect 122540 659770 122780 660010
rect 122870 659770 123110 660010
rect 123200 659770 123440 660010
rect 123530 659770 123770 660010
rect 123880 659770 124120 660010
rect 124210 659770 124450 660010
rect 124540 659770 124780 660010
rect 124870 659770 125110 660010
rect 125220 659770 125460 660010
rect 125550 659770 125790 660010
rect 125880 659770 126120 660010
rect 126210 659770 126450 660010
rect 126560 659770 126800 660010
rect 126890 659770 127130 660010
rect 127220 659770 127460 660010
rect 127550 659770 127790 660010
rect 127900 659770 128140 660010
rect 128230 659770 128470 660010
rect 128560 659770 128800 660010
rect 128890 659770 129130 660010
rect 129240 659770 129480 660010
rect 129570 659770 129810 660010
rect 129900 659770 130140 660010
rect 130230 659770 130470 660010
rect 130580 659770 130820 660010
rect 130910 659770 131150 660010
rect 131240 659770 131480 660010
rect 131570 659770 131810 660010
rect 131920 659770 132160 660010
rect 132250 659770 132490 660010
rect 132580 659770 132820 660010
rect 132910 659770 133150 660010
rect 122190 659440 122430 659680
rect 122540 659440 122780 659680
rect 122870 659440 123110 659680
rect 123200 659440 123440 659680
rect 123530 659440 123770 659680
rect 123880 659440 124120 659680
rect 124210 659440 124450 659680
rect 124540 659440 124780 659680
rect 124870 659440 125110 659680
rect 125220 659440 125460 659680
rect 125550 659440 125790 659680
rect 125880 659440 126120 659680
rect 126210 659440 126450 659680
rect 126560 659440 126800 659680
rect 126890 659440 127130 659680
rect 127220 659440 127460 659680
rect 127550 659440 127790 659680
rect 127900 659440 128140 659680
rect 128230 659440 128470 659680
rect 128560 659440 128800 659680
rect 128890 659440 129130 659680
rect 129240 659440 129480 659680
rect 129570 659440 129810 659680
rect 129900 659440 130140 659680
rect 130230 659440 130470 659680
rect 130580 659440 130820 659680
rect 130910 659440 131150 659680
rect 131240 659440 131480 659680
rect 131570 659440 131810 659680
rect 131920 659440 132160 659680
rect 132250 659440 132490 659680
rect 132580 659440 132820 659680
rect 132910 659440 133150 659680
rect 122190 659110 122430 659350
rect 122540 659110 122780 659350
rect 122870 659110 123110 659350
rect 123200 659110 123440 659350
rect 123530 659110 123770 659350
rect 123880 659110 124120 659350
rect 124210 659110 124450 659350
rect 124540 659110 124780 659350
rect 124870 659110 125110 659350
rect 125220 659110 125460 659350
rect 125550 659110 125790 659350
rect 125880 659110 126120 659350
rect 126210 659110 126450 659350
rect 126560 659110 126800 659350
rect 126890 659110 127130 659350
rect 127220 659110 127460 659350
rect 127550 659110 127790 659350
rect 127900 659110 128140 659350
rect 128230 659110 128470 659350
rect 128560 659110 128800 659350
rect 128890 659110 129130 659350
rect 129240 659110 129480 659350
rect 129570 659110 129810 659350
rect 129900 659110 130140 659350
rect 130230 659110 130470 659350
rect 130580 659110 130820 659350
rect 130910 659110 131150 659350
rect 131240 659110 131480 659350
rect 131570 659110 131810 659350
rect 131920 659110 132160 659350
rect 132250 659110 132490 659350
rect 132580 659110 132820 659350
rect 132910 659110 133150 659350
rect 122190 658760 122430 659000
rect 122540 658760 122780 659000
rect 122870 658760 123110 659000
rect 123200 658760 123440 659000
rect 123530 658760 123770 659000
rect 123880 658760 124120 659000
rect 124210 658760 124450 659000
rect 124540 658760 124780 659000
rect 124870 658760 125110 659000
rect 125220 658760 125460 659000
rect 125550 658760 125790 659000
rect 125880 658760 126120 659000
rect 126210 658760 126450 659000
rect 126560 658760 126800 659000
rect 126890 658760 127130 659000
rect 127220 658760 127460 659000
rect 127550 658760 127790 659000
rect 127900 658760 128140 659000
rect 128230 658760 128470 659000
rect 128560 658760 128800 659000
rect 128890 658760 129130 659000
rect 129240 658760 129480 659000
rect 129570 658760 129810 659000
rect 129900 658760 130140 659000
rect 130230 658760 130470 659000
rect 130580 658760 130820 659000
rect 130910 658760 131150 659000
rect 131240 658760 131480 659000
rect 131570 658760 131810 659000
rect 131920 658760 132160 659000
rect 132250 658760 132490 659000
rect 132580 658760 132820 659000
rect 132910 658760 133150 659000
rect 122190 658430 122430 658670
rect 122540 658430 122780 658670
rect 122870 658430 123110 658670
rect 123200 658430 123440 658670
rect 123530 658430 123770 658670
rect 123880 658430 124120 658670
rect 124210 658430 124450 658670
rect 124540 658430 124780 658670
rect 124870 658430 125110 658670
rect 125220 658430 125460 658670
rect 125550 658430 125790 658670
rect 125880 658430 126120 658670
rect 126210 658430 126450 658670
rect 126560 658430 126800 658670
rect 126890 658430 127130 658670
rect 127220 658430 127460 658670
rect 127550 658430 127790 658670
rect 127900 658430 128140 658670
rect 128230 658430 128470 658670
rect 128560 658430 128800 658670
rect 128890 658430 129130 658670
rect 129240 658430 129480 658670
rect 129570 658430 129810 658670
rect 129900 658430 130140 658670
rect 130230 658430 130470 658670
rect 130580 658430 130820 658670
rect 130910 658430 131150 658670
rect 131240 658430 131480 658670
rect 131570 658430 131810 658670
rect 131920 658430 132160 658670
rect 132250 658430 132490 658670
rect 132580 658430 132820 658670
rect 132910 658430 133150 658670
rect 122190 658100 122430 658340
rect 122540 658100 122780 658340
rect 122870 658100 123110 658340
rect 123200 658100 123440 658340
rect 123530 658100 123770 658340
rect 123880 658100 124120 658340
rect 124210 658100 124450 658340
rect 124540 658100 124780 658340
rect 124870 658100 125110 658340
rect 125220 658100 125460 658340
rect 125550 658100 125790 658340
rect 125880 658100 126120 658340
rect 126210 658100 126450 658340
rect 126560 658100 126800 658340
rect 126890 658100 127130 658340
rect 127220 658100 127460 658340
rect 127550 658100 127790 658340
rect 127900 658100 128140 658340
rect 128230 658100 128470 658340
rect 128560 658100 128800 658340
rect 128890 658100 129130 658340
rect 129240 658100 129480 658340
rect 129570 658100 129810 658340
rect 129900 658100 130140 658340
rect 130230 658100 130470 658340
rect 130580 658100 130820 658340
rect 130910 658100 131150 658340
rect 131240 658100 131480 658340
rect 131570 658100 131810 658340
rect 131920 658100 132160 658340
rect 132250 658100 132490 658340
rect 132580 658100 132820 658340
rect 132910 658100 133150 658340
rect 122190 657770 122430 658010
rect 122540 657770 122780 658010
rect 122870 657770 123110 658010
rect 123200 657770 123440 658010
rect 123530 657770 123770 658010
rect 123880 657770 124120 658010
rect 124210 657770 124450 658010
rect 124540 657770 124780 658010
rect 124870 657770 125110 658010
rect 125220 657770 125460 658010
rect 125550 657770 125790 658010
rect 125880 657770 126120 658010
rect 126210 657770 126450 658010
rect 126560 657770 126800 658010
rect 126890 657770 127130 658010
rect 127220 657770 127460 658010
rect 127550 657770 127790 658010
rect 127900 657770 128140 658010
rect 128230 657770 128470 658010
rect 128560 657770 128800 658010
rect 128890 657770 129130 658010
rect 129240 657770 129480 658010
rect 129570 657770 129810 658010
rect 129900 657770 130140 658010
rect 130230 657770 130470 658010
rect 130580 657770 130820 658010
rect 130910 657770 131150 658010
rect 131240 657770 131480 658010
rect 131570 657770 131810 658010
rect 131920 657770 132160 658010
rect 132250 657770 132490 658010
rect 132580 657770 132820 658010
rect 132910 657770 133150 658010
rect 122190 657420 122430 657660
rect 122540 657420 122780 657660
rect 122870 657420 123110 657660
rect 123200 657420 123440 657660
rect 123530 657420 123770 657660
rect 123880 657420 124120 657660
rect 124210 657420 124450 657660
rect 124540 657420 124780 657660
rect 124870 657420 125110 657660
rect 125220 657420 125460 657660
rect 125550 657420 125790 657660
rect 125880 657420 126120 657660
rect 126210 657420 126450 657660
rect 126560 657420 126800 657660
rect 126890 657420 127130 657660
rect 127220 657420 127460 657660
rect 127550 657420 127790 657660
rect 127900 657420 128140 657660
rect 128230 657420 128470 657660
rect 128560 657420 128800 657660
rect 128890 657420 129130 657660
rect 129240 657420 129480 657660
rect 129570 657420 129810 657660
rect 129900 657420 130140 657660
rect 130230 657420 130470 657660
rect 130580 657420 130820 657660
rect 130910 657420 131150 657660
rect 131240 657420 131480 657660
rect 131570 657420 131810 657660
rect 131920 657420 132160 657660
rect 132250 657420 132490 657660
rect 132580 657420 132820 657660
rect 132910 657420 133150 657660
rect 122190 657090 122430 657330
rect 122540 657090 122780 657330
rect 122870 657090 123110 657330
rect 123200 657090 123440 657330
rect 123530 657090 123770 657330
rect 123880 657090 124120 657330
rect 124210 657090 124450 657330
rect 124540 657090 124780 657330
rect 124870 657090 125110 657330
rect 125220 657090 125460 657330
rect 125550 657090 125790 657330
rect 125880 657090 126120 657330
rect 126210 657090 126450 657330
rect 126560 657090 126800 657330
rect 126890 657090 127130 657330
rect 127220 657090 127460 657330
rect 127550 657090 127790 657330
rect 127900 657090 128140 657330
rect 128230 657090 128470 657330
rect 128560 657090 128800 657330
rect 128890 657090 129130 657330
rect 129240 657090 129480 657330
rect 129570 657090 129810 657330
rect 129900 657090 130140 657330
rect 130230 657090 130470 657330
rect 130580 657090 130820 657330
rect 130910 657090 131150 657330
rect 131240 657090 131480 657330
rect 131570 657090 131810 657330
rect 131920 657090 132160 657330
rect 132250 657090 132490 657330
rect 132580 657090 132820 657330
rect 132910 657090 133150 657330
rect 122190 656760 122430 657000
rect 122540 656760 122780 657000
rect 122870 656760 123110 657000
rect 123200 656760 123440 657000
rect 123530 656760 123770 657000
rect 123880 656760 124120 657000
rect 124210 656760 124450 657000
rect 124540 656760 124780 657000
rect 124870 656760 125110 657000
rect 125220 656760 125460 657000
rect 125550 656760 125790 657000
rect 125880 656760 126120 657000
rect 126210 656760 126450 657000
rect 126560 656760 126800 657000
rect 126890 656760 127130 657000
rect 127220 656760 127460 657000
rect 127550 656760 127790 657000
rect 127900 656760 128140 657000
rect 128230 656760 128470 657000
rect 128560 656760 128800 657000
rect 128890 656760 129130 657000
rect 129240 656760 129480 657000
rect 129570 656760 129810 657000
rect 129900 656760 130140 657000
rect 130230 656760 130470 657000
rect 130580 656760 130820 657000
rect 130910 656760 131150 657000
rect 131240 656760 131480 657000
rect 131570 656760 131810 657000
rect 131920 656760 132160 657000
rect 132250 656760 132490 657000
rect 132580 656760 132820 657000
rect 132910 656760 133150 657000
rect 122190 656430 122430 656670
rect 122540 656430 122780 656670
rect 122870 656430 123110 656670
rect 123200 656430 123440 656670
rect 123530 656430 123770 656670
rect 123880 656430 124120 656670
rect 124210 656430 124450 656670
rect 124540 656430 124780 656670
rect 124870 656430 125110 656670
rect 125220 656430 125460 656670
rect 125550 656430 125790 656670
rect 125880 656430 126120 656670
rect 126210 656430 126450 656670
rect 126560 656430 126800 656670
rect 126890 656430 127130 656670
rect 127220 656430 127460 656670
rect 127550 656430 127790 656670
rect 127900 656430 128140 656670
rect 128230 656430 128470 656670
rect 128560 656430 128800 656670
rect 128890 656430 129130 656670
rect 129240 656430 129480 656670
rect 129570 656430 129810 656670
rect 129900 656430 130140 656670
rect 130230 656430 130470 656670
rect 130580 656430 130820 656670
rect 130910 656430 131150 656670
rect 131240 656430 131480 656670
rect 131570 656430 131810 656670
rect 131920 656430 132160 656670
rect 132250 656430 132490 656670
rect 132580 656430 132820 656670
rect 132910 656430 133150 656670
rect 122190 656080 122430 656320
rect 122540 656080 122780 656320
rect 122870 656080 123110 656320
rect 123200 656080 123440 656320
rect 123530 656080 123770 656320
rect 123880 656080 124120 656320
rect 124210 656080 124450 656320
rect 124540 656080 124780 656320
rect 124870 656080 125110 656320
rect 125220 656080 125460 656320
rect 125550 656080 125790 656320
rect 125880 656080 126120 656320
rect 126210 656080 126450 656320
rect 126560 656080 126800 656320
rect 126890 656080 127130 656320
rect 127220 656080 127460 656320
rect 127550 656080 127790 656320
rect 127900 656080 128140 656320
rect 128230 656080 128470 656320
rect 128560 656080 128800 656320
rect 128890 656080 129130 656320
rect 129240 656080 129480 656320
rect 129570 656080 129810 656320
rect 129900 656080 130140 656320
rect 130230 656080 130470 656320
rect 130580 656080 130820 656320
rect 130910 656080 131150 656320
rect 131240 656080 131480 656320
rect 131570 656080 131810 656320
rect 131920 656080 132160 656320
rect 132250 656080 132490 656320
rect 132580 656080 132820 656320
rect 132910 656080 133150 656320
rect 122190 655750 122430 655990
rect 122540 655750 122780 655990
rect 122870 655750 123110 655990
rect 123200 655750 123440 655990
rect 123530 655750 123770 655990
rect 123880 655750 124120 655990
rect 124210 655750 124450 655990
rect 124540 655750 124780 655990
rect 124870 655750 125110 655990
rect 125220 655750 125460 655990
rect 125550 655750 125790 655990
rect 125880 655750 126120 655990
rect 126210 655750 126450 655990
rect 126560 655750 126800 655990
rect 126890 655750 127130 655990
rect 127220 655750 127460 655990
rect 127550 655750 127790 655990
rect 127900 655750 128140 655990
rect 128230 655750 128470 655990
rect 128560 655750 128800 655990
rect 128890 655750 129130 655990
rect 129240 655750 129480 655990
rect 129570 655750 129810 655990
rect 129900 655750 130140 655990
rect 130230 655750 130470 655990
rect 130580 655750 130820 655990
rect 130910 655750 131150 655990
rect 131240 655750 131480 655990
rect 131570 655750 131810 655990
rect 131920 655750 132160 655990
rect 132250 655750 132490 655990
rect 132580 655750 132820 655990
rect 132910 655750 133150 655990
rect 122190 655420 122430 655660
rect 122540 655420 122780 655660
rect 122870 655420 123110 655660
rect 123200 655420 123440 655660
rect 123530 655420 123770 655660
rect 123880 655420 124120 655660
rect 124210 655420 124450 655660
rect 124540 655420 124780 655660
rect 124870 655420 125110 655660
rect 125220 655420 125460 655660
rect 125550 655420 125790 655660
rect 125880 655420 126120 655660
rect 126210 655420 126450 655660
rect 126560 655420 126800 655660
rect 126890 655420 127130 655660
rect 127220 655420 127460 655660
rect 127550 655420 127790 655660
rect 127900 655420 128140 655660
rect 128230 655420 128470 655660
rect 128560 655420 128800 655660
rect 128890 655420 129130 655660
rect 129240 655420 129480 655660
rect 129570 655420 129810 655660
rect 129900 655420 130140 655660
rect 130230 655420 130470 655660
rect 130580 655420 130820 655660
rect 130910 655420 131150 655660
rect 131240 655420 131480 655660
rect 131570 655420 131810 655660
rect 131920 655420 132160 655660
rect 132250 655420 132490 655660
rect 132580 655420 132820 655660
rect 132910 655420 133150 655660
rect 122190 655090 122430 655330
rect 122540 655090 122780 655330
rect 122870 655090 123110 655330
rect 123200 655090 123440 655330
rect 123530 655090 123770 655330
rect 123880 655090 124120 655330
rect 124210 655090 124450 655330
rect 124540 655090 124780 655330
rect 124870 655090 125110 655330
rect 125220 655090 125460 655330
rect 125550 655090 125790 655330
rect 125880 655090 126120 655330
rect 126210 655090 126450 655330
rect 126560 655090 126800 655330
rect 126890 655090 127130 655330
rect 127220 655090 127460 655330
rect 127550 655090 127790 655330
rect 127900 655090 128140 655330
rect 128230 655090 128470 655330
rect 128560 655090 128800 655330
rect 128890 655090 129130 655330
rect 129240 655090 129480 655330
rect 129570 655090 129810 655330
rect 129900 655090 130140 655330
rect 130230 655090 130470 655330
rect 130580 655090 130820 655330
rect 130910 655090 131150 655330
rect 131240 655090 131480 655330
rect 131570 655090 131810 655330
rect 131920 655090 132160 655330
rect 132250 655090 132490 655330
rect 132580 655090 132820 655330
rect 132910 655090 133150 655330
rect 122190 654740 122430 654980
rect 122540 654740 122780 654980
rect 122870 654740 123110 654980
rect 123200 654740 123440 654980
rect 123530 654740 123770 654980
rect 123880 654740 124120 654980
rect 124210 654740 124450 654980
rect 124540 654740 124780 654980
rect 124870 654740 125110 654980
rect 125220 654740 125460 654980
rect 125550 654740 125790 654980
rect 125880 654740 126120 654980
rect 126210 654740 126450 654980
rect 126560 654740 126800 654980
rect 126890 654740 127130 654980
rect 127220 654740 127460 654980
rect 127550 654740 127790 654980
rect 127900 654740 128140 654980
rect 128230 654740 128470 654980
rect 128560 654740 128800 654980
rect 128890 654740 129130 654980
rect 129240 654740 129480 654980
rect 129570 654740 129810 654980
rect 129900 654740 130140 654980
rect 130230 654740 130470 654980
rect 130580 654740 130820 654980
rect 130910 654740 131150 654980
rect 131240 654740 131480 654980
rect 131570 654740 131810 654980
rect 131920 654740 132160 654980
rect 132250 654740 132490 654980
rect 132580 654740 132820 654980
rect 132910 654740 133150 654980
rect 122190 654410 122430 654650
rect 122540 654410 122780 654650
rect 122870 654410 123110 654650
rect 123200 654410 123440 654650
rect 123530 654410 123770 654650
rect 123880 654410 124120 654650
rect 124210 654410 124450 654650
rect 124540 654410 124780 654650
rect 124870 654410 125110 654650
rect 125220 654410 125460 654650
rect 125550 654410 125790 654650
rect 125880 654410 126120 654650
rect 126210 654410 126450 654650
rect 126560 654410 126800 654650
rect 126890 654410 127130 654650
rect 127220 654410 127460 654650
rect 127550 654410 127790 654650
rect 127900 654410 128140 654650
rect 128230 654410 128470 654650
rect 128560 654410 128800 654650
rect 128890 654410 129130 654650
rect 129240 654410 129480 654650
rect 129570 654410 129810 654650
rect 129900 654410 130140 654650
rect 130230 654410 130470 654650
rect 130580 654410 130820 654650
rect 130910 654410 131150 654650
rect 131240 654410 131480 654650
rect 131570 654410 131810 654650
rect 131920 654410 132160 654650
rect 132250 654410 132490 654650
rect 132580 654410 132820 654650
rect 132910 654410 133150 654650
rect 122190 654080 122430 654320
rect 122540 654080 122780 654320
rect 122870 654080 123110 654320
rect 123200 654080 123440 654320
rect 123530 654080 123770 654320
rect 123880 654080 124120 654320
rect 124210 654080 124450 654320
rect 124540 654080 124780 654320
rect 124870 654080 125110 654320
rect 125220 654080 125460 654320
rect 125550 654080 125790 654320
rect 125880 654080 126120 654320
rect 126210 654080 126450 654320
rect 126560 654080 126800 654320
rect 126890 654080 127130 654320
rect 127220 654080 127460 654320
rect 127550 654080 127790 654320
rect 127900 654080 128140 654320
rect 128230 654080 128470 654320
rect 128560 654080 128800 654320
rect 128890 654080 129130 654320
rect 129240 654080 129480 654320
rect 129570 654080 129810 654320
rect 129900 654080 130140 654320
rect 130230 654080 130470 654320
rect 130580 654080 130820 654320
rect 130910 654080 131150 654320
rect 131240 654080 131480 654320
rect 131570 654080 131810 654320
rect 131920 654080 132160 654320
rect 132250 654080 132490 654320
rect 132580 654080 132820 654320
rect 132910 654080 133150 654320
rect 122190 653750 122430 653990
rect 122540 653750 122780 653990
rect 122870 653750 123110 653990
rect 123200 653750 123440 653990
rect 123530 653750 123770 653990
rect 123880 653750 124120 653990
rect 124210 653750 124450 653990
rect 124540 653750 124780 653990
rect 124870 653750 125110 653990
rect 125220 653750 125460 653990
rect 125550 653750 125790 653990
rect 125880 653750 126120 653990
rect 126210 653750 126450 653990
rect 126560 653750 126800 653990
rect 126890 653750 127130 653990
rect 127220 653750 127460 653990
rect 127550 653750 127790 653990
rect 127900 653750 128140 653990
rect 128230 653750 128470 653990
rect 128560 653750 128800 653990
rect 128890 653750 129130 653990
rect 129240 653750 129480 653990
rect 129570 653750 129810 653990
rect 129900 653750 130140 653990
rect 130230 653750 130470 653990
rect 130580 653750 130820 653990
rect 130910 653750 131150 653990
rect 131240 653750 131480 653990
rect 131570 653750 131810 653990
rect 131920 653750 132160 653990
rect 132250 653750 132490 653990
rect 132580 653750 132820 653990
rect 132910 653750 133150 653990
rect 122190 653400 122430 653640
rect 122540 653400 122780 653640
rect 122870 653400 123110 653640
rect 123200 653400 123440 653640
rect 123530 653400 123770 653640
rect 123880 653400 124120 653640
rect 124210 653400 124450 653640
rect 124540 653400 124780 653640
rect 124870 653400 125110 653640
rect 125220 653400 125460 653640
rect 125550 653400 125790 653640
rect 125880 653400 126120 653640
rect 126210 653400 126450 653640
rect 126560 653400 126800 653640
rect 126890 653400 127130 653640
rect 127220 653400 127460 653640
rect 127550 653400 127790 653640
rect 127900 653400 128140 653640
rect 128230 653400 128470 653640
rect 128560 653400 128800 653640
rect 128890 653400 129130 653640
rect 129240 653400 129480 653640
rect 129570 653400 129810 653640
rect 129900 653400 130140 653640
rect 130230 653400 130470 653640
rect 130580 653400 130820 653640
rect 130910 653400 131150 653640
rect 131240 653400 131480 653640
rect 131570 653400 131810 653640
rect 131920 653400 132160 653640
rect 132250 653400 132490 653640
rect 132580 653400 132820 653640
rect 132910 653400 133150 653640
rect 122190 653070 122430 653310
rect 122540 653070 122780 653310
rect 122870 653070 123110 653310
rect 123200 653070 123440 653310
rect 123530 653070 123770 653310
rect 123880 653070 124120 653310
rect 124210 653070 124450 653310
rect 124540 653070 124780 653310
rect 124870 653070 125110 653310
rect 125220 653070 125460 653310
rect 125550 653070 125790 653310
rect 125880 653070 126120 653310
rect 126210 653070 126450 653310
rect 126560 653070 126800 653310
rect 126890 653070 127130 653310
rect 127220 653070 127460 653310
rect 127550 653070 127790 653310
rect 127900 653070 128140 653310
rect 128230 653070 128470 653310
rect 128560 653070 128800 653310
rect 128890 653070 129130 653310
rect 129240 653070 129480 653310
rect 129570 653070 129810 653310
rect 129900 653070 130140 653310
rect 130230 653070 130470 653310
rect 130580 653070 130820 653310
rect 130910 653070 131150 653310
rect 131240 653070 131480 653310
rect 131570 653070 131810 653310
rect 131920 653070 132160 653310
rect 132250 653070 132490 653310
rect 132580 653070 132820 653310
rect 132910 653070 133150 653310
rect 122190 652740 122430 652980
rect 122540 652740 122780 652980
rect 122870 652740 123110 652980
rect 123200 652740 123440 652980
rect 123530 652740 123770 652980
rect 123880 652740 124120 652980
rect 124210 652740 124450 652980
rect 124540 652740 124780 652980
rect 124870 652740 125110 652980
rect 125220 652740 125460 652980
rect 125550 652740 125790 652980
rect 125880 652740 126120 652980
rect 126210 652740 126450 652980
rect 126560 652740 126800 652980
rect 126890 652740 127130 652980
rect 127220 652740 127460 652980
rect 127550 652740 127790 652980
rect 127900 652740 128140 652980
rect 128230 652740 128470 652980
rect 128560 652740 128800 652980
rect 128890 652740 129130 652980
rect 129240 652740 129480 652980
rect 129570 652740 129810 652980
rect 129900 652740 130140 652980
rect 130230 652740 130470 652980
rect 130580 652740 130820 652980
rect 130910 652740 131150 652980
rect 131240 652740 131480 652980
rect 131570 652740 131810 652980
rect 131920 652740 132160 652980
rect 132250 652740 132490 652980
rect 132580 652740 132820 652980
rect 132910 652740 133150 652980
rect 122190 652410 122430 652650
rect 122540 652410 122780 652650
rect 122870 652410 123110 652650
rect 123200 652410 123440 652650
rect 123530 652410 123770 652650
rect 123880 652410 124120 652650
rect 124210 652410 124450 652650
rect 124540 652410 124780 652650
rect 124870 652410 125110 652650
rect 125220 652410 125460 652650
rect 125550 652410 125790 652650
rect 125880 652410 126120 652650
rect 126210 652410 126450 652650
rect 126560 652410 126800 652650
rect 126890 652410 127130 652650
rect 127220 652410 127460 652650
rect 127550 652410 127790 652650
rect 127900 652410 128140 652650
rect 128230 652410 128470 652650
rect 128560 652410 128800 652650
rect 128890 652410 129130 652650
rect 129240 652410 129480 652650
rect 129570 652410 129810 652650
rect 129900 652410 130140 652650
rect 130230 652410 130470 652650
rect 130580 652410 130820 652650
rect 130910 652410 131150 652650
rect 131240 652410 131480 652650
rect 131570 652410 131810 652650
rect 131920 652410 132160 652650
rect 132250 652410 132490 652650
rect 132580 652410 132820 652650
rect 132910 652410 133150 652650
rect 122190 652060 122430 652300
rect 122540 652060 122780 652300
rect 122870 652060 123110 652300
rect 123200 652060 123440 652300
rect 123530 652060 123770 652300
rect 123880 652060 124120 652300
rect 124210 652060 124450 652300
rect 124540 652060 124780 652300
rect 124870 652060 125110 652300
rect 125220 652060 125460 652300
rect 125550 652060 125790 652300
rect 125880 652060 126120 652300
rect 126210 652060 126450 652300
rect 126560 652060 126800 652300
rect 126890 652060 127130 652300
rect 127220 652060 127460 652300
rect 127550 652060 127790 652300
rect 127900 652060 128140 652300
rect 128230 652060 128470 652300
rect 128560 652060 128800 652300
rect 128890 652060 129130 652300
rect 129240 652060 129480 652300
rect 129570 652060 129810 652300
rect 129900 652060 130140 652300
rect 130230 652060 130470 652300
rect 130580 652060 130820 652300
rect 130910 652060 131150 652300
rect 131240 652060 131480 652300
rect 131570 652060 131810 652300
rect 131920 652060 132160 652300
rect 132250 652060 132490 652300
rect 132580 652060 132820 652300
rect 132910 652060 133150 652300
rect 122190 651730 122430 651970
rect 122540 651730 122780 651970
rect 122870 651730 123110 651970
rect 123200 651730 123440 651970
rect 123530 651730 123770 651970
rect 123880 651730 124120 651970
rect 124210 651730 124450 651970
rect 124540 651730 124780 651970
rect 124870 651730 125110 651970
rect 125220 651730 125460 651970
rect 125550 651730 125790 651970
rect 125880 651730 126120 651970
rect 126210 651730 126450 651970
rect 126560 651730 126800 651970
rect 126890 651730 127130 651970
rect 127220 651730 127460 651970
rect 127550 651730 127790 651970
rect 127900 651730 128140 651970
rect 128230 651730 128470 651970
rect 128560 651730 128800 651970
rect 128890 651730 129130 651970
rect 129240 651730 129480 651970
rect 129570 651730 129810 651970
rect 129900 651730 130140 651970
rect 130230 651730 130470 651970
rect 130580 651730 130820 651970
rect 130910 651730 131150 651970
rect 131240 651730 131480 651970
rect 131570 651730 131810 651970
rect 131920 651730 132160 651970
rect 132250 651730 132490 651970
rect 132580 651730 132820 651970
rect 132910 651730 133150 651970
rect 122190 651400 122430 651640
rect 122540 651400 122780 651640
rect 122870 651400 123110 651640
rect 123200 651400 123440 651640
rect 123530 651400 123770 651640
rect 123880 651400 124120 651640
rect 124210 651400 124450 651640
rect 124540 651400 124780 651640
rect 124870 651400 125110 651640
rect 125220 651400 125460 651640
rect 125550 651400 125790 651640
rect 125880 651400 126120 651640
rect 126210 651400 126450 651640
rect 126560 651400 126800 651640
rect 126890 651400 127130 651640
rect 127220 651400 127460 651640
rect 127550 651400 127790 651640
rect 127900 651400 128140 651640
rect 128230 651400 128470 651640
rect 128560 651400 128800 651640
rect 128890 651400 129130 651640
rect 129240 651400 129480 651640
rect 129570 651400 129810 651640
rect 129900 651400 130140 651640
rect 130230 651400 130470 651640
rect 130580 651400 130820 651640
rect 130910 651400 131150 651640
rect 131240 651400 131480 651640
rect 131570 651400 131810 651640
rect 131920 651400 132160 651640
rect 132250 651400 132490 651640
rect 132580 651400 132820 651640
rect 132910 651400 133150 651640
rect 122190 651070 122430 651310
rect 122540 651070 122780 651310
rect 122870 651070 123110 651310
rect 123200 651070 123440 651310
rect 123530 651070 123770 651310
rect 123880 651070 124120 651310
rect 124210 651070 124450 651310
rect 124540 651070 124780 651310
rect 124870 651070 125110 651310
rect 125220 651070 125460 651310
rect 125550 651070 125790 651310
rect 125880 651070 126120 651310
rect 126210 651070 126450 651310
rect 126560 651070 126800 651310
rect 126890 651070 127130 651310
rect 127220 651070 127460 651310
rect 127550 651070 127790 651310
rect 127900 651070 128140 651310
rect 128230 651070 128470 651310
rect 128560 651070 128800 651310
rect 128890 651070 129130 651310
rect 129240 651070 129480 651310
rect 129570 651070 129810 651310
rect 129900 651070 130140 651310
rect 130230 651070 130470 651310
rect 130580 651070 130820 651310
rect 130910 651070 131150 651310
rect 131240 651070 131480 651310
rect 131570 651070 131810 651310
rect 131920 651070 132160 651310
rect 132250 651070 132490 651310
rect 132580 651070 132820 651310
rect 132910 651070 133150 651310
rect 122190 650720 122430 650960
rect 122540 650720 122780 650960
rect 122870 650720 123110 650960
rect 123200 650720 123440 650960
rect 123530 650720 123770 650960
rect 123880 650720 124120 650960
rect 124210 650720 124450 650960
rect 124540 650720 124780 650960
rect 124870 650720 125110 650960
rect 125220 650720 125460 650960
rect 125550 650720 125790 650960
rect 125880 650720 126120 650960
rect 126210 650720 126450 650960
rect 126560 650720 126800 650960
rect 126890 650720 127130 650960
rect 127220 650720 127460 650960
rect 127550 650720 127790 650960
rect 127900 650720 128140 650960
rect 128230 650720 128470 650960
rect 128560 650720 128800 650960
rect 128890 650720 129130 650960
rect 129240 650720 129480 650960
rect 129570 650720 129810 650960
rect 129900 650720 130140 650960
rect 130230 650720 130470 650960
rect 130580 650720 130820 650960
rect 130910 650720 131150 650960
rect 131240 650720 131480 650960
rect 131570 650720 131810 650960
rect 131920 650720 132160 650960
rect 132250 650720 132490 650960
rect 132580 650720 132820 650960
rect 132910 650720 133150 650960
rect 122190 650390 122430 650630
rect 122540 650390 122780 650630
rect 122870 650390 123110 650630
rect 123200 650390 123440 650630
rect 123530 650390 123770 650630
rect 123880 650390 124120 650630
rect 124210 650390 124450 650630
rect 124540 650390 124780 650630
rect 124870 650390 125110 650630
rect 125220 650390 125460 650630
rect 125550 650390 125790 650630
rect 125880 650390 126120 650630
rect 126210 650390 126450 650630
rect 126560 650390 126800 650630
rect 126890 650390 127130 650630
rect 127220 650390 127460 650630
rect 127550 650390 127790 650630
rect 127900 650390 128140 650630
rect 128230 650390 128470 650630
rect 128560 650390 128800 650630
rect 128890 650390 129130 650630
rect 129240 650390 129480 650630
rect 129570 650390 129810 650630
rect 129900 650390 130140 650630
rect 130230 650390 130470 650630
rect 130580 650390 130820 650630
rect 130910 650390 131150 650630
rect 131240 650390 131480 650630
rect 131570 650390 131810 650630
rect 131920 650390 132160 650630
rect 132250 650390 132490 650630
rect 132580 650390 132820 650630
rect 132910 650390 133150 650630
rect 122190 650060 122430 650300
rect 122540 650060 122780 650300
rect 122870 650060 123110 650300
rect 123200 650060 123440 650300
rect 123530 650060 123770 650300
rect 123880 650060 124120 650300
rect 124210 650060 124450 650300
rect 124540 650060 124780 650300
rect 124870 650060 125110 650300
rect 125220 650060 125460 650300
rect 125550 650060 125790 650300
rect 125880 650060 126120 650300
rect 126210 650060 126450 650300
rect 126560 650060 126800 650300
rect 126890 650060 127130 650300
rect 127220 650060 127460 650300
rect 127550 650060 127790 650300
rect 127900 650060 128140 650300
rect 128230 650060 128470 650300
rect 128560 650060 128800 650300
rect 128890 650060 129130 650300
rect 129240 650060 129480 650300
rect 129570 650060 129810 650300
rect 129900 650060 130140 650300
rect 130230 650060 130470 650300
rect 130580 650060 130820 650300
rect 130910 650060 131150 650300
rect 131240 650060 131480 650300
rect 131570 650060 131810 650300
rect 131920 650060 132160 650300
rect 132250 650060 132490 650300
rect 132580 650060 132820 650300
rect 132910 650060 133150 650300
rect 122190 649730 122430 649970
rect 122540 649730 122780 649970
rect 122870 649730 123110 649970
rect 123200 649730 123440 649970
rect 123530 649730 123770 649970
rect 123880 649730 124120 649970
rect 124210 649730 124450 649970
rect 124540 649730 124780 649970
rect 124870 649730 125110 649970
rect 125220 649730 125460 649970
rect 125550 649730 125790 649970
rect 125880 649730 126120 649970
rect 126210 649730 126450 649970
rect 126560 649730 126800 649970
rect 126890 649730 127130 649970
rect 127220 649730 127460 649970
rect 127550 649730 127790 649970
rect 127900 649730 128140 649970
rect 128230 649730 128470 649970
rect 128560 649730 128800 649970
rect 128890 649730 129130 649970
rect 129240 649730 129480 649970
rect 129570 649730 129810 649970
rect 129900 649730 130140 649970
rect 130230 649730 130470 649970
rect 130580 649730 130820 649970
rect 130910 649730 131150 649970
rect 131240 649730 131480 649970
rect 131570 649730 131810 649970
rect 131920 649730 132160 649970
rect 132250 649730 132490 649970
rect 132580 649730 132820 649970
rect 132910 649730 133150 649970
rect 122190 649380 122430 649620
rect 122540 649380 122780 649620
rect 122870 649380 123110 649620
rect 123200 649380 123440 649620
rect 123530 649380 123770 649620
rect 123880 649380 124120 649620
rect 124210 649380 124450 649620
rect 124540 649380 124780 649620
rect 124870 649380 125110 649620
rect 125220 649380 125460 649620
rect 125550 649380 125790 649620
rect 125880 649380 126120 649620
rect 126210 649380 126450 649620
rect 126560 649380 126800 649620
rect 126890 649380 127130 649620
rect 127220 649380 127460 649620
rect 127550 649380 127790 649620
rect 127900 649380 128140 649620
rect 128230 649380 128470 649620
rect 128560 649380 128800 649620
rect 128890 649380 129130 649620
rect 129240 649380 129480 649620
rect 129570 649380 129810 649620
rect 129900 649380 130140 649620
rect 130230 649380 130470 649620
rect 130580 649380 130820 649620
rect 130910 649380 131150 649620
rect 131240 649380 131480 649620
rect 131570 649380 131810 649620
rect 131920 649380 132160 649620
rect 132250 649380 132490 649620
rect 132580 649380 132820 649620
rect 132910 649380 133150 649620
rect 133570 660100 133810 660340
rect 133920 660100 134160 660340
rect 134250 660100 134490 660340
rect 134580 660100 134820 660340
rect 134910 660100 135150 660340
rect 135260 660100 135500 660340
rect 135590 660100 135830 660340
rect 135920 660100 136160 660340
rect 136250 660100 136490 660340
rect 136600 660100 136840 660340
rect 136930 660100 137170 660340
rect 137260 660100 137500 660340
rect 137590 660100 137830 660340
rect 137940 660100 138180 660340
rect 138270 660100 138510 660340
rect 138600 660100 138840 660340
rect 138930 660100 139170 660340
rect 139280 660100 139520 660340
rect 139610 660100 139850 660340
rect 139940 660100 140180 660340
rect 140270 660100 140510 660340
rect 140620 660100 140860 660340
rect 140950 660100 141190 660340
rect 141280 660100 141520 660340
rect 141610 660100 141850 660340
rect 141960 660100 142200 660340
rect 142290 660100 142530 660340
rect 142620 660100 142860 660340
rect 142950 660100 143190 660340
rect 143300 660100 143540 660340
rect 143630 660100 143870 660340
rect 143960 660100 144200 660340
rect 144290 660100 144530 660340
rect 133570 659770 133810 660010
rect 133920 659770 134160 660010
rect 134250 659770 134490 660010
rect 134580 659770 134820 660010
rect 134910 659770 135150 660010
rect 135260 659770 135500 660010
rect 135590 659770 135830 660010
rect 135920 659770 136160 660010
rect 136250 659770 136490 660010
rect 136600 659770 136840 660010
rect 136930 659770 137170 660010
rect 137260 659770 137500 660010
rect 137590 659770 137830 660010
rect 137940 659770 138180 660010
rect 138270 659770 138510 660010
rect 138600 659770 138840 660010
rect 138930 659770 139170 660010
rect 139280 659770 139520 660010
rect 139610 659770 139850 660010
rect 139940 659770 140180 660010
rect 140270 659770 140510 660010
rect 140620 659770 140860 660010
rect 140950 659770 141190 660010
rect 141280 659770 141520 660010
rect 141610 659770 141850 660010
rect 141960 659770 142200 660010
rect 142290 659770 142530 660010
rect 142620 659770 142860 660010
rect 142950 659770 143190 660010
rect 143300 659770 143540 660010
rect 143630 659770 143870 660010
rect 143960 659770 144200 660010
rect 144290 659770 144530 660010
rect 133570 659440 133810 659680
rect 133920 659440 134160 659680
rect 134250 659440 134490 659680
rect 134580 659440 134820 659680
rect 134910 659440 135150 659680
rect 135260 659440 135500 659680
rect 135590 659440 135830 659680
rect 135920 659440 136160 659680
rect 136250 659440 136490 659680
rect 136600 659440 136840 659680
rect 136930 659440 137170 659680
rect 137260 659440 137500 659680
rect 137590 659440 137830 659680
rect 137940 659440 138180 659680
rect 138270 659440 138510 659680
rect 138600 659440 138840 659680
rect 138930 659440 139170 659680
rect 139280 659440 139520 659680
rect 139610 659440 139850 659680
rect 139940 659440 140180 659680
rect 140270 659440 140510 659680
rect 140620 659440 140860 659680
rect 140950 659440 141190 659680
rect 141280 659440 141520 659680
rect 141610 659440 141850 659680
rect 141960 659440 142200 659680
rect 142290 659440 142530 659680
rect 142620 659440 142860 659680
rect 142950 659440 143190 659680
rect 143300 659440 143540 659680
rect 143630 659440 143870 659680
rect 143960 659440 144200 659680
rect 144290 659440 144530 659680
rect 133570 659110 133810 659350
rect 133920 659110 134160 659350
rect 134250 659110 134490 659350
rect 134580 659110 134820 659350
rect 134910 659110 135150 659350
rect 135260 659110 135500 659350
rect 135590 659110 135830 659350
rect 135920 659110 136160 659350
rect 136250 659110 136490 659350
rect 136600 659110 136840 659350
rect 136930 659110 137170 659350
rect 137260 659110 137500 659350
rect 137590 659110 137830 659350
rect 137940 659110 138180 659350
rect 138270 659110 138510 659350
rect 138600 659110 138840 659350
rect 138930 659110 139170 659350
rect 139280 659110 139520 659350
rect 139610 659110 139850 659350
rect 139940 659110 140180 659350
rect 140270 659110 140510 659350
rect 140620 659110 140860 659350
rect 140950 659110 141190 659350
rect 141280 659110 141520 659350
rect 141610 659110 141850 659350
rect 141960 659110 142200 659350
rect 142290 659110 142530 659350
rect 142620 659110 142860 659350
rect 142950 659110 143190 659350
rect 143300 659110 143540 659350
rect 143630 659110 143870 659350
rect 143960 659110 144200 659350
rect 144290 659110 144530 659350
rect 133570 658760 133810 659000
rect 133920 658760 134160 659000
rect 134250 658760 134490 659000
rect 134580 658760 134820 659000
rect 134910 658760 135150 659000
rect 135260 658760 135500 659000
rect 135590 658760 135830 659000
rect 135920 658760 136160 659000
rect 136250 658760 136490 659000
rect 136600 658760 136840 659000
rect 136930 658760 137170 659000
rect 137260 658760 137500 659000
rect 137590 658760 137830 659000
rect 137940 658760 138180 659000
rect 138270 658760 138510 659000
rect 138600 658760 138840 659000
rect 138930 658760 139170 659000
rect 139280 658760 139520 659000
rect 139610 658760 139850 659000
rect 139940 658760 140180 659000
rect 140270 658760 140510 659000
rect 140620 658760 140860 659000
rect 140950 658760 141190 659000
rect 141280 658760 141520 659000
rect 141610 658760 141850 659000
rect 141960 658760 142200 659000
rect 142290 658760 142530 659000
rect 142620 658760 142860 659000
rect 142950 658760 143190 659000
rect 143300 658760 143540 659000
rect 143630 658760 143870 659000
rect 143960 658760 144200 659000
rect 144290 658760 144530 659000
rect 133570 658430 133810 658670
rect 133920 658430 134160 658670
rect 134250 658430 134490 658670
rect 134580 658430 134820 658670
rect 134910 658430 135150 658670
rect 135260 658430 135500 658670
rect 135590 658430 135830 658670
rect 135920 658430 136160 658670
rect 136250 658430 136490 658670
rect 136600 658430 136840 658670
rect 136930 658430 137170 658670
rect 137260 658430 137500 658670
rect 137590 658430 137830 658670
rect 137940 658430 138180 658670
rect 138270 658430 138510 658670
rect 138600 658430 138840 658670
rect 138930 658430 139170 658670
rect 139280 658430 139520 658670
rect 139610 658430 139850 658670
rect 139940 658430 140180 658670
rect 140270 658430 140510 658670
rect 140620 658430 140860 658670
rect 140950 658430 141190 658670
rect 141280 658430 141520 658670
rect 141610 658430 141850 658670
rect 141960 658430 142200 658670
rect 142290 658430 142530 658670
rect 142620 658430 142860 658670
rect 142950 658430 143190 658670
rect 143300 658430 143540 658670
rect 143630 658430 143870 658670
rect 143960 658430 144200 658670
rect 144290 658430 144530 658670
rect 133570 658100 133810 658340
rect 133920 658100 134160 658340
rect 134250 658100 134490 658340
rect 134580 658100 134820 658340
rect 134910 658100 135150 658340
rect 135260 658100 135500 658340
rect 135590 658100 135830 658340
rect 135920 658100 136160 658340
rect 136250 658100 136490 658340
rect 136600 658100 136840 658340
rect 136930 658100 137170 658340
rect 137260 658100 137500 658340
rect 137590 658100 137830 658340
rect 137940 658100 138180 658340
rect 138270 658100 138510 658340
rect 138600 658100 138840 658340
rect 138930 658100 139170 658340
rect 139280 658100 139520 658340
rect 139610 658100 139850 658340
rect 139940 658100 140180 658340
rect 140270 658100 140510 658340
rect 140620 658100 140860 658340
rect 140950 658100 141190 658340
rect 141280 658100 141520 658340
rect 141610 658100 141850 658340
rect 141960 658100 142200 658340
rect 142290 658100 142530 658340
rect 142620 658100 142860 658340
rect 142950 658100 143190 658340
rect 143300 658100 143540 658340
rect 143630 658100 143870 658340
rect 143960 658100 144200 658340
rect 144290 658100 144530 658340
rect 133570 657770 133810 658010
rect 133920 657770 134160 658010
rect 134250 657770 134490 658010
rect 134580 657770 134820 658010
rect 134910 657770 135150 658010
rect 135260 657770 135500 658010
rect 135590 657770 135830 658010
rect 135920 657770 136160 658010
rect 136250 657770 136490 658010
rect 136600 657770 136840 658010
rect 136930 657770 137170 658010
rect 137260 657770 137500 658010
rect 137590 657770 137830 658010
rect 137940 657770 138180 658010
rect 138270 657770 138510 658010
rect 138600 657770 138840 658010
rect 138930 657770 139170 658010
rect 139280 657770 139520 658010
rect 139610 657770 139850 658010
rect 139940 657770 140180 658010
rect 140270 657770 140510 658010
rect 140620 657770 140860 658010
rect 140950 657770 141190 658010
rect 141280 657770 141520 658010
rect 141610 657770 141850 658010
rect 141960 657770 142200 658010
rect 142290 657770 142530 658010
rect 142620 657770 142860 658010
rect 142950 657770 143190 658010
rect 143300 657770 143540 658010
rect 143630 657770 143870 658010
rect 143960 657770 144200 658010
rect 144290 657770 144530 658010
rect 133570 657420 133810 657660
rect 133920 657420 134160 657660
rect 134250 657420 134490 657660
rect 134580 657420 134820 657660
rect 134910 657420 135150 657660
rect 135260 657420 135500 657660
rect 135590 657420 135830 657660
rect 135920 657420 136160 657660
rect 136250 657420 136490 657660
rect 136600 657420 136840 657660
rect 136930 657420 137170 657660
rect 137260 657420 137500 657660
rect 137590 657420 137830 657660
rect 137940 657420 138180 657660
rect 138270 657420 138510 657660
rect 138600 657420 138840 657660
rect 138930 657420 139170 657660
rect 139280 657420 139520 657660
rect 139610 657420 139850 657660
rect 139940 657420 140180 657660
rect 140270 657420 140510 657660
rect 140620 657420 140860 657660
rect 140950 657420 141190 657660
rect 141280 657420 141520 657660
rect 141610 657420 141850 657660
rect 141960 657420 142200 657660
rect 142290 657420 142530 657660
rect 142620 657420 142860 657660
rect 142950 657420 143190 657660
rect 143300 657420 143540 657660
rect 143630 657420 143870 657660
rect 143960 657420 144200 657660
rect 144290 657420 144530 657660
rect 133570 657090 133810 657330
rect 133920 657090 134160 657330
rect 134250 657090 134490 657330
rect 134580 657090 134820 657330
rect 134910 657090 135150 657330
rect 135260 657090 135500 657330
rect 135590 657090 135830 657330
rect 135920 657090 136160 657330
rect 136250 657090 136490 657330
rect 136600 657090 136840 657330
rect 136930 657090 137170 657330
rect 137260 657090 137500 657330
rect 137590 657090 137830 657330
rect 137940 657090 138180 657330
rect 138270 657090 138510 657330
rect 138600 657090 138840 657330
rect 138930 657090 139170 657330
rect 139280 657090 139520 657330
rect 139610 657090 139850 657330
rect 139940 657090 140180 657330
rect 140270 657090 140510 657330
rect 140620 657090 140860 657330
rect 140950 657090 141190 657330
rect 141280 657090 141520 657330
rect 141610 657090 141850 657330
rect 141960 657090 142200 657330
rect 142290 657090 142530 657330
rect 142620 657090 142860 657330
rect 142950 657090 143190 657330
rect 143300 657090 143540 657330
rect 143630 657090 143870 657330
rect 143960 657090 144200 657330
rect 144290 657090 144530 657330
rect 133570 656760 133810 657000
rect 133920 656760 134160 657000
rect 134250 656760 134490 657000
rect 134580 656760 134820 657000
rect 134910 656760 135150 657000
rect 135260 656760 135500 657000
rect 135590 656760 135830 657000
rect 135920 656760 136160 657000
rect 136250 656760 136490 657000
rect 136600 656760 136840 657000
rect 136930 656760 137170 657000
rect 137260 656760 137500 657000
rect 137590 656760 137830 657000
rect 137940 656760 138180 657000
rect 138270 656760 138510 657000
rect 138600 656760 138840 657000
rect 138930 656760 139170 657000
rect 139280 656760 139520 657000
rect 139610 656760 139850 657000
rect 139940 656760 140180 657000
rect 140270 656760 140510 657000
rect 140620 656760 140860 657000
rect 140950 656760 141190 657000
rect 141280 656760 141520 657000
rect 141610 656760 141850 657000
rect 141960 656760 142200 657000
rect 142290 656760 142530 657000
rect 142620 656760 142860 657000
rect 142950 656760 143190 657000
rect 143300 656760 143540 657000
rect 143630 656760 143870 657000
rect 143960 656760 144200 657000
rect 144290 656760 144530 657000
rect 133570 656430 133810 656670
rect 133920 656430 134160 656670
rect 134250 656430 134490 656670
rect 134580 656430 134820 656670
rect 134910 656430 135150 656670
rect 135260 656430 135500 656670
rect 135590 656430 135830 656670
rect 135920 656430 136160 656670
rect 136250 656430 136490 656670
rect 136600 656430 136840 656670
rect 136930 656430 137170 656670
rect 137260 656430 137500 656670
rect 137590 656430 137830 656670
rect 137940 656430 138180 656670
rect 138270 656430 138510 656670
rect 138600 656430 138840 656670
rect 138930 656430 139170 656670
rect 139280 656430 139520 656670
rect 139610 656430 139850 656670
rect 139940 656430 140180 656670
rect 140270 656430 140510 656670
rect 140620 656430 140860 656670
rect 140950 656430 141190 656670
rect 141280 656430 141520 656670
rect 141610 656430 141850 656670
rect 141960 656430 142200 656670
rect 142290 656430 142530 656670
rect 142620 656430 142860 656670
rect 142950 656430 143190 656670
rect 143300 656430 143540 656670
rect 143630 656430 143870 656670
rect 143960 656430 144200 656670
rect 144290 656430 144530 656670
rect 133570 656080 133810 656320
rect 133920 656080 134160 656320
rect 134250 656080 134490 656320
rect 134580 656080 134820 656320
rect 134910 656080 135150 656320
rect 135260 656080 135500 656320
rect 135590 656080 135830 656320
rect 135920 656080 136160 656320
rect 136250 656080 136490 656320
rect 136600 656080 136840 656320
rect 136930 656080 137170 656320
rect 137260 656080 137500 656320
rect 137590 656080 137830 656320
rect 137940 656080 138180 656320
rect 138270 656080 138510 656320
rect 138600 656080 138840 656320
rect 138930 656080 139170 656320
rect 139280 656080 139520 656320
rect 139610 656080 139850 656320
rect 139940 656080 140180 656320
rect 140270 656080 140510 656320
rect 140620 656080 140860 656320
rect 140950 656080 141190 656320
rect 141280 656080 141520 656320
rect 141610 656080 141850 656320
rect 141960 656080 142200 656320
rect 142290 656080 142530 656320
rect 142620 656080 142860 656320
rect 142950 656080 143190 656320
rect 143300 656080 143540 656320
rect 143630 656080 143870 656320
rect 143960 656080 144200 656320
rect 144290 656080 144530 656320
rect 133570 655750 133810 655990
rect 133920 655750 134160 655990
rect 134250 655750 134490 655990
rect 134580 655750 134820 655990
rect 134910 655750 135150 655990
rect 135260 655750 135500 655990
rect 135590 655750 135830 655990
rect 135920 655750 136160 655990
rect 136250 655750 136490 655990
rect 136600 655750 136840 655990
rect 136930 655750 137170 655990
rect 137260 655750 137500 655990
rect 137590 655750 137830 655990
rect 137940 655750 138180 655990
rect 138270 655750 138510 655990
rect 138600 655750 138840 655990
rect 138930 655750 139170 655990
rect 139280 655750 139520 655990
rect 139610 655750 139850 655990
rect 139940 655750 140180 655990
rect 140270 655750 140510 655990
rect 140620 655750 140860 655990
rect 140950 655750 141190 655990
rect 141280 655750 141520 655990
rect 141610 655750 141850 655990
rect 141960 655750 142200 655990
rect 142290 655750 142530 655990
rect 142620 655750 142860 655990
rect 142950 655750 143190 655990
rect 143300 655750 143540 655990
rect 143630 655750 143870 655990
rect 143960 655750 144200 655990
rect 144290 655750 144530 655990
rect 133570 655420 133810 655660
rect 133920 655420 134160 655660
rect 134250 655420 134490 655660
rect 134580 655420 134820 655660
rect 134910 655420 135150 655660
rect 135260 655420 135500 655660
rect 135590 655420 135830 655660
rect 135920 655420 136160 655660
rect 136250 655420 136490 655660
rect 136600 655420 136840 655660
rect 136930 655420 137170 655660
rect 137260 655420 137500 655660
rect 137590 655420 137830 655660
rect 137940 655420 138180 655660
rect 138270 655420 138510 655660
rect 138600 655420 138840 655660
rect 138930 655420 139170 655660
rect 139280 655420 139520 655660
rect 139610 655420 139850 655660
rect 139940 655420 140180 655660
rect 140270 655420 140510 655660
rect 140620 655420 140860 655660
rect 140950 655420 141190 655660
rect 141280 655420 141520 655660
rect 141610 655420 141850 655660
rect 141960 655420 142200 655660
rect 142290 655420 142530 655660
rect 142620 655420 142860 655660
rect 142950 655420 143190 655660
rect 143300 655420 143540 655660
rect 143630 655420 143870 655660
rect 143960 655420 144200 655660
rect 144290 655420 144530 655660
rect 133570 655090 133810 655330
rect 133920 655090 134160 655330
rect 134250 655090 134490 655330
rect 134580 655090 134820 655330
rect 134910 655090 135150 655330
rect 135260 655090 135500 655330
rect 135590 655090 135830 655330
rect 135920 655090 136160 655330
rect 136250 655090 136490 655330
rect 136600 655090 136840 655330
rect 136930 655090 137170 655330
rect 137260 655090 137500 655330
rect 137590 655090 137830 655330
rect 137940 655090 138180 655330
rect 138270 655090 138510 655330
rect 138600 655090 138840 655330
rect 138930 655090 139170 655330
rect 139280 655090 139520 655330
rect 139610 655090 139850 655330
rect 139940 655090 140180 655330
rect 140270 655090 140510 655330
rect 140620 655090 140860 655330
rect 140950 655090 141190 655330
rect 141280 655090 141520 655330
rect 141610 655090 141850 655330
rect 141960 655090 142200 655330
rect 142290 655090 142530 655330
rect 142620 655090 142860 655330
rect 142950 655090 143190 655330
rect 143300 655090 143540 655330
rect 143630 655090 143870 655330
rect 143960 655090 144200 655330
rect 144290 655090 144530 655330
rect 133570 654740 133810 654980
rect 133920 654740 134160 654980
rect 134250 654740 134490 654980
rect 134580 654740 134820 654980
rect 134910 654740 135150 654980
rect 135260 654740 135500 654980
rect 135590 654740 135830 654980
rect 135920 654740 136160 654980
rect 136250 654740 136490 654980
rect 136600 654740 136840 654980
rect 136930 654740 137170 654980
rect 137260 654740 137500 654980
rect 137590 654740 137830 654980
rect 137940 654740 138180 654980
rect 138270 654740 138510 654980
rect 138600 654740 138840 654980
rect 138930 654740 139170 654980
rect 139280 654740 139520 654980
rect 139610 654740 139850 654980
rect 139940 654740 140180 654980
rect 140270 654740 140510 654980
rect 140620 654740 140860 654980
rect 140950 654740 141190 654980
rect 141280 654740 141520 654980
rect 141610 654740 141850 654980
rect 141960 654740 142200 654980
rect 142290 654740 142530 654980
rect 142620 654740 142860 654980
rect 142950 654740 143190 654980
rect 143300 654740 143540 654980
rect 143630 654740 143870 654980
rect 143960 654740 144200 654980
rect 144290 654740 144530 654980
rect 133570 654410 133810 654650
rect 133920 654410 134160 654650
rect 134250 654410 134490 654650
rect 134580 654410 134820 654650
rect 134910 654410 135150 654650
rect 135260 654410 135500 654650
rect 135590 654410 135830 654650
rect 135920 654410 136160 654650
rect 136250 654410 136490 654650
rect 136600 654410 136840 654650
rect 136930 654410 137170 654650
rect 137260 654410 137500 654650
rect 137590 654410 137830 654650
rect 137940 654410 138180 654650
rect 138270 654410 138510 654650
rect 138600 654410 138840 654650
rect 138930 654410 139170 654650
rect 139280 654410 139520 654650
rect 139610 654410 139850 654650
rect 139940 654410 140180 654650
rect 140270 654410 140510 654650
rect 140620 654410 140860 654650
rect 140950 654410 141190 654650
rect 141280 654410 141520 654650
rect 141610 654410 141850 654650
rect 141960 654410 142200 654650
rect 142290 654410 142530 654650
rect 142620 654410 142860 654650
rect 142950 654410 143190 654650
rect 143300 654410 143540 654650
rect 143630 654410 143870 654650
rect 143960 654410 144200 654650
rect 144290 654410 144530 654650
rect 133570 654080 133810 654320
rect 133920 654080 134160 654320
rect 134250 654080 134490 654320
rect 134580 654080 134820 654320
rect 134910 654080 135150 654320
rect 135260 654080 135500 654320
rect 135590 654080 135830 654320
rect 135920 654080 136160 654320
rect 136250 654080 136490 654320
rect 136600 654080 136840 654320
rect 136930 654080 137170 654320
rect 137260 654080 137500 654320
rect 137590 654080 137830 654320
rect 137940 654080 138180 654320
rect 138270 654080 138510 654320
rect 138600 654080 138840 654320
rect 138930 654080 139170 654320
rect 139280 654080 139520 654320
rect 139610 654080 139850 654320
rect 139940 654080 140180 654320
rect 140270 654080 140510 654320
rect 140620 654080 140860 654320
rect 140950 654080 141190 654320
rect 141280 654080 141520 654320
rect 141610 654080 141850 654320
rect 141960 654080 142200 654320
rect 142290 654080 142530 654320
rect 142620 654080 142860 654320
rect 142950 654080 143190 654320
rect 143300 654080 143540 654320
rect 143630 654080 143870 654320
rect 143960 654080 144200 654320
rect 144290 654080 144530 654320
rect 133570 653750 133810 653990
rect 133920 653750 134160 653990
rect 134250 653750 134490 653990
rect 134580 653750 134820 653990
rect 134910 653750 135150 653990
rect 135260 653750 135500 653990
rect 135590 653750 135830 653990
rect 135920 653750 136160 653990
rect 136250 653750 136490 653990
rect 136600 653750 136840 653990
rect 136930 653750 137170 653990
rect 137260 653750 137500 653990
rect 137590 653750 137830 653990
rect 137940 653750 138180 653990
rect 138270 653750 138510 653990
rect 138600 653750 138840 653990
rect 138930 653750 139170 653990
rect 139280 653750 139520 653990
rect 139610 653750 139850 653990
rect 139940 653750 140180 653990
rect 140270 653750 140510 653990
rect 140620 653750 140860 653990
rect 140950 653750 141190 653990
rect 141280 653750 141520 653990
rect 141610 653750 141850 653990
rect 141960 653750 142200 653990
rect 142290 653750 142530 653990
rect 142620 653750 142860 653990
rect 142950 653750 143190 653990
rect 143300 653750 143540 653990
rect 143630 653750 143870 653990
rect 143960 653750 144200 653990
rect 144290 653750 144530 653990
rect 133570 653400 133810 653640
rect 133920 653400 134160 653640
rect 134250 653400 134490 653640
rect 134580 653400 134820 653640
rect 134910 653400 135150 653640
rect 135260 653400 135500 653640
rect 135590 653400 135830 653640
rect 135920 653400 136160 653640
rect 136250 653400 136490 653640
rect 136600 653400 136840 653640
rect 136930 653400 137170 653640
rect 137260 653400 137500 653640
rect 137590 653400 137830 653640
rect 137940 653400 138180 653640
rect 138270 653400 138510 653640
rect 138600 653400 138840 653640
rect 138930 653400 139170 653640
rect 139280 653400 139520 653640
rect 139610 653400 139850 653640
rect 139940 653400 140180 653640
rect 140270 653400 140510 653640
rect 140620 653400 140860 653640
rect 140950 653400 141190 653640
rect 141280 653400 141520 653640
rect 141610 653400 141850 653640
rect 141960 653400 142200 653640
rect 142290 653400 142530 653640
rect 142620 653400 142860 653640
rect 142950 653400 143190 653640
rect 143300 653400 143540 653640
rect 143630 653400 143870 653640
rect 143960 653400 144200 653640
rect 144290 653400 144530 653640
rect 133570 653070 133810 653310
rect 133920 653070 134160 653310
rect 134250 653070 134490 653310
rect 134580 653070 134820 653310
rect 134910 653070 135150 653310
rect 135260 653070 135500 653310
rect 135590 653070 135830 653310
rect 135920 653070 136160 653310
rect 136250 653070 136490 653310
rect 136600 653070 136840 653310
rect 136930 653070 137170 653310
rect 137260 653070 137500 653310
rect 137590 653070 137830 653310
rect 137940 653070 138180 653310
rect 138270 653070 138510 653310
rect 138600 653070 138840 653310
rect 138930 653070 139170 653310
rect 139280 653070 139520 653310
rect 139610 653070 139850 653310
rect 139940 653070 140180 653310
rect 140270 653070 140510 653310
rect 140620 653070 140860 653310
rect 140950 653070 141190 653310
rect 141280 653070 141520 653310
rect 141610 653070 141850 653310
rect 141960 653070 142200 653310
rect 142290 653070 142530 653310
rect 142620 653070 142860 653310
rect 142950 653070 143190 653310
rect 143300 653070 143540 653310
rect 143630 653070 143870 653310
rect 143960 653070 144200 653310
rect 144290 653070 144530 653310
rect 133570 652740 133810 652980
rect 133920 652740 134160 652980
rect 134250 652740 134490 652980
rect 134580 652740 134820 652980
rect 134910 652740 135150 652980
rect 135260 652740 135500 652980
rect 135590 652740 135830 652980
rect 135920 652740 136160 652980
rect 136250 652740 136490 652980
rect 136600 652740 136840 652980
rect 136930 652740 137170 652980
rect 137260 652740 137500 652980
rect 137590 652740 137830 652980
rect 137940 652740 138180 652980
rect 138270 652740 138510 652980
rect 138600 652740 138840 652980
rect 138930 652740 139170 652980
rect 139280 652740 139520 652980
rect 139610 652740 139850 652980
rect 139940 652740 140180 652980
rect 140270 652740 140510 652980
rect 140620 652740 140860 652980
rect 140950 652740 141190 652980
rect 141280 652740 141520 652980
rect 141610 652740 141850 652980
rect 141960 652740 142200 652980
rect 142290 652740 142530 652980
rect 142620 652740 142860 652980
rect 142950 652740 143190 652980
rect 143300 652740 143540 652980
rect 143630 652740 143870 652980
rect 143960 652740 144200 652980
rect 144290 652740 144530 652980
rect 133570 652410 133810 652650
rect 133920 652410 134160 652650
rect 134250 652410 134490 652650
rect 134580 652410 134820 652650
rect 134910 652410 135150 652650
rect 135260 652410 135500 652650
rect 135590 652410 135830 652650
rect 135920 652410 136160 652650
rect 136250 652410 136490 652650
rect 136600 652410 136840 652650
rect 136930 652410 137170 652650
rect 137260 652410 137500 652650
rect 137590 652410 137830 652650
rect 137940 652410 138180 652650
rect 138270 652410 138510 652650
rect 138600 652410 138840 652650
rect 138930 652410 139170 652650
rect 139280 652410 139520 652650
rect 139610 652410 139850 652650
rect 139940 652410 140180 652650
rect 140270 652410 140510 652650
rect 140620 652410 140860 652650
rect 140950 652410 141190 652650
rect 141280 652410 141520 652650
rect 141610 652410 141850 652650
rect 141960 652410 142200 652650
rect 142290 652410 142530 652650
rect 142620 652410 142860 652650
rect 142950 652410 143190 652650
rect 143300 652410 143540 652650
rect 143630 652410 143870 652650
rect 143960 652410 144200 652650
rect 144290 652410 144530 652650
rect 133570 652060 133810 652300
rect 133920 652060 134160 652300
rect 134250 652060 134490 652300
rect 134580 652060 134820 652300
rect 134910 652060 135150 652300
rect 135260 652060 135500 652300
rect 135590 652060 135830 652300
rect 135920 652060 136160 652300
rect 136250 652060 136490 652300
rect 136600 652060 136840 652300
rect 136930 652060 137170 652300
rect 137260 652060 137500 652300
rect 137590 652060 137830 652300
rect 137940 652060 138180 652300
rect 138270 652060 138510 652300
rect 138600 652060 138840 652300
rect 138930 652060 139170 652300
rect 139280 652060 139520 652300
rect 139610 652060 139850 652300
rect 139940 652060 140180 652300
rect 140270 652060 140510 652300
rect 140620 652060 140860 652300
rect 140950 652060 141190 652300
rect 141280 652060 141520 652300
rect 141610 652060 141850 652300
rect 141960 652060 142200 652300
rect 142290 652060 142530 652300
rect 142620 652060 142860 652300
rect 142950 652060 143190 652300
rect 143300 652060 143540 652300
rect 143630 652060 143870 652300
rect 143960 652060 144200 652300
rect 144290 652060 144530 652300
rect 133570 651730 133810 651970
rect 133920 651730 134160 651970
rect 134250 651730 134490 651970
rect 134580 651730 134820 651970
rect 134910 651730 135150 651970
rect 135260 651730 135500 651970
rect 135590 651730 135830 651970
rect 135920 651730 136160 651970
rect 136250 651730 136490 651970
rect 136600 651730 136840 651970
rect 136930 651730 137170 651970
rect 137260 651730 137500 651970
rect 137590 651730 137830 651970
rect 137940 651730 138180 651970
rect 138270 651730 138510 651970
rect 138600 651730 138840 651970
rect 138930 651730 139170 651970
rect 139280 651730 139520 651970
rect 139610 651730 139850 651970
rect 139940 651730 140180 651970
rect 140270 651730 140510 651970
rect 140620 651730 140860 651970
rect 140950 651730 141190 651970
rect 141280 651730 141520 651970
rect 141610 651730 141850 651970
rect 141960 651730 142200 651970
rect 142290 651730 142530 651970
rect 142620 651730 142860 651970
rect 142950 651730 143190 651970
rect 143300 651730 143540 651970
rect 143630 651730 143870 651970
rect 143960 651730 144200 651970
rect 144290 651730 144530 651970
rect 133570 651400 133810 651640
rect 133920 651400 134160 651640
rect 134250 651400 134490 651640
rect 134580 651400 134820 651640
rect 134910 651400 135150 651640
rect 135260 651400 135500 651640
rect 135590 651400 135830 651640
rect 135920 651400 136160 651640
rect 136250 651400 136490 651640
rect 136600 651400 136840 651640
rect 136930 651400 137170 651640
rect 137260 651400 137500 651640
rect 137590 651400 137830 651640
rect 137940 651400 138180 651640
rect 138270 651400 138510 651640
rect 138600 651400 138840 651640
rect 138930 651400 139170 651640
rect 139280 651400 139520 651640
rect 139610 651400 139850 651640
rect 139940 651400 140180 651640
rect 140270 651400 140510 651640
rect 140620 651400 140860 651640
rect 140950 651400 141190 651640
rect 141280 651400 141520 651640
rect 141610 651400 141850 651640
rect 141960 651400 142200 651640
rect 142290 651400 142530 651640
rect 142620 651400 142860 651640
rect 142950 651400 143190 651640
rect 143300 651400 143540 651640
rect 143630 651400 143870 651640
rect 143960 651400 144200 651640
rect 144290 651400 144530 651640
rect 133570 651070 133810 651310
rect 133920 651070 134160 651310
rect 134250 651070 134490 651310
rect 134580 651070 134820 651310
rect 134910 651070 135150 651310
rect 135260 651070 135500 651310
rect 135590 651070 135830 651310
rect 135920 651070 136160 651310
rect 136250 651070 136490 651310
rect 136600 651070 136840 651310
rect 136930 651070 137170 651310
rect 137260 651070 137500 651310
rect 137590 651070 137830 651310
rect 137940 651070 138180 651310
rect 138270 651070 138510 651310
rect 138600 651070 138840 651310
rect 138930 651070 139170 651310
rect 139280 651070 139520 651310
rect 139610 651070 139850 651310
rect 139940 651070 140180 651310
rect 140270 651070 140510 651310
rect 140620 651070 140860 651310
rect 140950 651070 141190 651310
rect 141280 651070 141520 651310
rect 141610 651070 141850 651310
rect 141960 651070 142200 651310
rect 142290 651070 142530 651310
rect 142620 651070 142860 651310
rect 142950 651070 143190 651310
rect 143300 651070 143540 651310
rect 143630 651070 143870 651310
rect 143960 651070 144200 651310
rect 144290 651070 144530 651310
rect 133570 650720 133810 650960
rect 133920 650720 134160 650960
rect 134250 650720 134490 650960
rect 134580 650720 134820 650960
rect 134910 650720 135150 650960
rect 135260 650720 135500 650960
rect 135590 650720 135830 650960
rect 135920 650720 136160 650960
rect 136250 650720 136490 650960
rect 136600 650720 136840 650960
rect 136930 650720 137170 650960
rect 137260 650720 137500 650960
rect 137590 650720 137830 650960
rect 137940 650720 138180 650960
rect 138270 650720 138510 650960
rect 138600 650720 138840 650960
rect 138930 650720 139170 650960
rect 139280 650720 139520 650960
rect 139610 650720 139850 650960
rect 139940 650720 140180 650960
rect 140270 650720 140510 650960
rect 140620 650720 140860 650960
rect 140950 650720 141190 650960
rect 141280 650720 141520 650960
rect 141610 650720 141850 650960
rect 141960 650720 142200 650960
rect 142290 650720 142530 650960
rect 142620 650720 142860 650960
rect 142950 650720 143190 650960
rect 143300 650720 143540 650960
rect 143630 650720 143870 650960
rect 143960 650720 144200 650960
rect 144290 650720 144530 650960
rect 133570 650390 133810 650630
rect 133920 650390 134160 650630
rect 134250 650390 134490 650630
rect 134580 650390 134820 650630
rect 134910 650390 135150 650630
rect 135260 650390 135500 650630
rect 135590 650390 135830 650630
rect 135920 650390 136160 650630
rect 136250 650390 136490 650630
rect 136600 650390 136840 650630
rect 136930 650390 137170 650630
rect 137260 650390 137500 650630
rect 137590 650390 137830 650630
rect 137940 650390 138180 650630
rect 138270 650390 138510 650630
rect 138600 650390 138840 650630
rect 138930 650390 139170 650630
rect 139280 650390 139520 650630
rect 139610 650390 139850 650630
rect 139940 650390 140180 650630
rect 140270 650390 140510 650630
rect 140620 650390 140860 650630
rect 140950 650390 141190 650630
rect 141280 650390 141520 650630
rect 141610 650390 141850 650630
rect 141960 650390 142200 650630
rect 142290 650390 142530 650630
rect 142620 650390 142860 650630
rect 142950 650390 143190 650630
rect 143300 650390 143540 650630
rect 143630 650390 143870 650630
rect 143960 650390 144200 650630
rect 144290 650390 144530 650630
rect 133570 650060 133810 650300
rect 133920 650060 134160 650300
rect 134250 650060 134490 650300
rect 134580 650060 134820 650300
rect 134910 650060 135150 650300
rect 135260 650060 135500 650300
rect 135590 650060 135830 650300
rect 135920 650060 136160 650300
rect 136250 650060 136490 650300
rect 136600 650060 136840 650300
rect 136930 650060 137170 650300
rect 137260 650060 137500 650300
rect 137590 650060 137830 650300
rect 137940 650060 138180 650300
rect 138270 650060 138510 650300
rect 138600 650060 138840 650300
rect 138930 650060 139170 650300
rect 139280 650060 139520 650300
rect 139610 650060 139850 650300
rect 139940 650060 140180 650300
rect 140270 650060 140510 650300
rect 140620 650060 140860 650300
rect 140950 650060 141190 650300
rect 141280 650060 141520 650300
rect 141610 650060 141850 650300
rect 141960 650060 142200 650300
rect 142290 650060 142530 650300
rect 142620 650060 142860 650300
rect 142950 650060 143190 650300
rect 143300 650060 143540 650300
rect 143630 650060 143870 650300
rect 143960 650060 144200 650300
rect 144290 650060 144530 650300
rect 133570 649730 133810 649970
rect 133920 649730 134160 649970
rect 134250 649730 134490 649970
rect 134580 649730 134820 649970
rect 134910 649730 135150 649970
rect 135260 649730 135500 649970
rect 135590 649730 135830 649970
rect 135920 649730 136160 649970
rect 136250 649730 136490 649970
rect 136600 649730 136840 649970
rect 136930 649730 137170 649970
rect 137260 649730 137500 649970
rect 137590 649730 137830 649970
rect 137940 649730 138180 649970
rect 138270 649730 138510 649970
rect 138600 649730 138840 649970
rect 138930 649730 139170 649970
rect 139280 649730 139520 649970
rect 139610 649730 139850 649970
rect 139940 649730 140180 649970
rect 140270 649730 140510 649970
rect 140620 649730 140860 649970
rect 140950 649730 141190 649970
rect 141280 649730 141520 649970
rect 141610 649730 141850 649970
rect 141960 649730 142200 649970
rect 142290 649730 142530 649970
rect 142620 649730 142860 649970
rect 142950 649730 143190 649970
rect 143300 649730 143540 649970
rect 143630 649730 143870 649970
rect 143960 649730 144200 649970
rect 144290 649730 144530 649970
rect 133570 649380 133810 649620
rect 133920 649380 134160 649620
rect 134250 649380 134490 649620
rect 134580 649380 134820 649620
rect 134910 649380 135150 649620
rect 135260 649380 135500 649620
rect 135590 649380 135830 649620
rect 135920 649380 136160 649620
rect 136250 649380 136490 649620
rect 136600 649380 136840 649620
rect 136930 649380 137170 649620
rect 137260 649380 137500 649620
rect 137590 649380 137830 649620
rect 137940 649380 138180 649620
rect 138270 649380 138510 649620
rect 138600 649380 138840 649620
rect 138930 649380 139170 649620
rect 139280 649380 139520 649620
rect 139610 649380 139850 649620
rect 139940 649380 140180 649620
rect 140270 649380 140510 649620
rect 140620 649380 140860 649620
rect 140950 649380 141190 649620
rect 141280 649380 141520 649620
rect 141610 649380 141850 649620
rect 141960 649380 142200 649620
rect 142290 649380 142530 649620
rect 142620 649380 142860 649620
rect 142950 649380 143190 649620
rect 143300 649380 143540 649620
rect 143630 649380 143870 649620
rect 143960 649380 144200 649620
rect 144290 649380 144530 649620
rect 144950 660100 145190 660340
rect 145300 660100 145540 660340
rect 145630 660100 145870 660340
rect 145960 660100 146200 660340
rect 146290 660100 146530 660340
rect 146640 660100 146880 660340
rect 146970 660100 147210 660340
rect 147300 660100 147540 660340
rect 147630 660100 147870 660340
rect 147980 660100 148220 660340
rect 148310 660100 148550 660340
rect 148640 660100 148880 660340
rect 148970 660100 149210 660340
rect 149320 660100 149560 660340
rect 149650 660100 149890 660340
rect 149980 660100 150220 660340
rect 150310 660100 150550 660340
rect 150660 660100 150900 660340
rect 150990 660100 151230 660340
rect 151320 660100 151560 660340
rect 151650 660100 151890 660340
rect 152000 660100 152240 660340
rect 152330 660100 152570 660340
rect 152660 660100 152900 660340
rect 152990 660100 153230 660340
rect 153340 660100 153580 660340
rect 153670 660100 153910 660340
rect 154000 660100 154240 660340
rect 154330 660100 154570 660340
rect 154680 660100 154920 660340
rect 155010 660100 155250 660340
rect 155340 660100 155580 660340
rect 155670 660100 155910 660340
rect 144950 659770 145190 660010
rect 145300 659770 145540 660010
rect 145630 659770 145870 660010
rect 145960 659770 146200 660010
rect 146290 659770 146530 660010
rect 146640 659770 146880 660010
rect 146970 659770 147210 660010
rect 147300 659770 147540 660010
rect 147630 659770 147870 660010
rect 147980 659770 148220 660010
rect 148310 659770 148550 660010
rect 148640 659770 148880 660010
rect 148970 659770 149210 660010
rect 149320 659770 149560 660010
rect 149650 659770 149890 660010
rect 149980 659770 150220 660010
rect 150310 659770 150550 660010
rect 150660 659770 150900 660010
rect 150990 659770 151230 660010
rect 151320 659770 151560 660010
rect 151650 659770 151890 660010
rect 152000 659770 152240 660010
rect 152330 659770 152570 660010
rect 152660 659770 152900 660010
rect 152990 659770 153230 660010
rect 153340 659770 153580 660010
rect 153670 659770 153910 660010
rect 154000 659770 154240 660010
rect 154330 659770 154570 660010
rect 154680 659770 154920 660010
rect 155010 659770 155250 660010
rect 155340 659770 155580 660010
rect 155670 659770 155910 660010
rect 144950 659440 145190 659680
rect 145300 659440 145540 659680
rect 145630 659440 145870 659680
rect 145960 659440 146200 659680
rect 146290 659440 146530 659680
rect 146640 659440 146880 659680
rect 146970 659440 147210 659680
rect 147300 659440 147540 659680
rect 147630 659440 147870 659680
rect 147980 659440 148220 659680
rect 148310 659440 148550 659680
rect 148640 659440 148880 659680
rect 148970 659440 149210 659680
rect 149320 659440 149560 659680
rect 149650 659440 149890 659680
rect 149980 659440 150220 659680
rect 150310 659440 150550 659680
rect 150660 659440 150900 659680
rect 150990 659440 151230 659680
rect 151320 659440 151560 659680
rect 151650 659440 151890 659680
rect 152000 659440 152240 659680
rect 152330 659440 152570 659680
rect 152660 659440 152900 659680
rect 152990 659440 153230 659680
rect 153340 659440 153580 659680
rect 153670 659440 153910 659680
rect 154000 659440 154240 659680
rect 154330 659440 154570 659680
rect 154680 659440 154920 659680
rect 155010 659440 155250 659680
rect 155340 659440 155580 659680
rect 155670 659440 155910 659680
rect 144950 659110 145190 659350
rect 145300 659110 145540 659350
rect 145630 659110 145870 659350
rect 145960 659110 146200 659350
rect 146290 659110 146530 659350
rect 146640 659110 146880 659350
rect 146970 659110 147210 659350
rect 147300 659110 147540 659350
rect 147630 659110 147870 659350
rect 147980 659110 148220 659350
rect 148310 659110 148550 659350
rect 148640 659110 148880 659350
rect 148970 659110 149210 659350
rect 149320 659110 149560 659350
rect 149650 659110 149890 659350
rect 149980 659110 150220 659350
rect 150310 659110 150550 659350
rect 150660 659110 150900 659350
rect 150990 659110 151230 659350
rect 151320 659110 151560 659350
rect 151650 659110 151890 659350
rect 152000 659110 152240 659350
rect 152330 659110 152570 659350
rect 152660 659110 152900 659350
rect 152990 659110 153230 659350
rect 153340 659110 153580 659350
rect 153670 659110 153910 659350
rect 154000 659110 154240 659350
rect 154330 659110 154570 659350
rect 154680 659110 154920 659350
rect 155010 659110 155250 659350
rect 155340 659110 155580 659350
rect 155670 659110 155910 659350
rect 144950 658760 145190 659000
rect 145300 658760 145540 659000
rect 145630 658760 145870 659000
rect 145960 658760 146200 659000
rect 146290 658760 146530 659000
rect 146640 658760 146880 659000
rect 146970 658760 147210 659000
rect 147300 658760 147540 659000
rect 147630 658760 147870 659000
rect 147980 658760 148220 659000
rect 148310 658760 148550 659000
rect 148640 658760 148880 659000
rect 148970 658760 149210 659000
rect 149320 658760 149560 659000
rect 149650 658760 149890 659000
rect 149980 658760 150220 659000
rect 150310 658760 150550 659000
rect 150660 658760 150900 659000
rect 150990 658760 151230 659000
rect 151320 658760 151560 659000
rect 151650 658760 151890 659000
rect 152000 658760 152240 659000
rect 152330 658760 152570 659000
rect 152660 658760 152900 659000
rect 152990 658760 153230 659000
rect 153340 658760 153580 659000
rect 153670 658760 153910 659000
rect 154000 658760 154240 659000
rect 154330 658760 154570 659000
rect 154680 658760 154920 659000
rect 155010 658760 155250 659000
rect 155340 658760 155580 659000
rect 155670 658760 155910 659000
rect 144950 658430 145190 658670
rect 145300 658430 145540 658670
rect 145630 658430 145870 658670
rect 145960 658430 146200 658670
rect 146290 658430 146530 658670
rect 146640 658430 146880 658670
rect 146970 658430 147210 658670
rect 147300 658430 147540 658670
rect 147630 658430 147870 658670
rect 147980 658430 148220 658670
rect 148310 658430 148550 658670
rect 148640 658430 148880 658670
rect 148970 658430 149210 658670
rect 149320 658430 149560 658670
rect 149650 658430 149890 658670
rect 149980 658430 150220 658670
rect 150310 658430 150550 658670
rect 150660 658430 150900 658670
rect 150990 658430 151230 658670
rect 151320 658430 151560 658670
rect 151650 658430 151890 658670
rect 152000 658430 152240 658670
rect 152330 658430 152570 658670
rect 152660 658430 152900 658670
rect 152990 658430 153230 658670
rect 153340 658430 153580 658670
rect 153670 658430 153910 658670
rect 154000 658430 154240 658670
rect 154330 658430 154570 658670
rect 154680 658430 154920 658670
rect 155010 658430 155250 658670
rect 155340 658430 155580 658670
rect 155670 658430 155910 658670
rect 144950 658100 145190 658340
rect 145300 658100 145540 658340
rect 145630 658100 145870 658340
rect 145960 658100 146200 658340
rect 146290 658100 146530 658340
rect 146640 658100 146880 658340
rect 146970 658100 147210 658340
rect 147300 658100 147540 658340
rect 147630 658100 147870 658340
rect 147980 658100 148220 658340
rect 148310 658100 148550 658340
rect 148640 658100 148880 658340
rect 148970 658100 149210 658340
rect 149320 658100 149560 658340
rect 149650 658100 149890 658340
rect 149980 658100 150220 658340
rect 150310 658100 150550 658340
rect 150660 658100 150900 658340
rect 150990 658100 151230 658340
rect 151320 658100 151560 658340
rect 151650 658100 151890 658340
rect 152000 658100 152240 658340
rect 152330 658100 152570 658340
rect 152660 658100 152900 658340
rect 152990 658100 153230 658340
rect 153340 658100 153580 658340
rect 153670 658100 153910 658340
rect 154000 658100 154240 658340
rect 154330 658100 154570 658340
rect 154680 658100 154920 658340
rect 155010 658100 155250 658340
rect 155340 658100 155580 658340
rect 155670 658100 155910 658340
rect 144950 657770 145190 658010
rect 145300 657770 145540 658010
rect 145630 657770 145870 658010
rect 145960 657770 146200 658010
rect 146290 657770 146530 658010
rect 146640 657770 146880 658010
rect 146970 657770 147210 658010
rect 147300 657770 147540 658010
rect 147630 657770 147870 658010
rect 147980 657770 148220 658010
rect 148310 657770 148550 658010
rect 148640 657770 148880 658010
rect 148970 657770 149210 658010
rect 149320 657770 149560 658010
rect 149650 657770 149890 658010
rect 149980 657770 150220 658010
rect 150310 657770 150550 658010
rect 150660 657770 150900 658010
rect 150990 657770 151230 658010
rect 151320 657770 151560 658010
rect 151650 657770 151890 658010
rect 152000 657770 152240 658010
rect 152330 657770 152570 658010
rect 152660 657770 152900 658010
rect 152990 657770 153230 658010
rect 153340 657770 153580 658010
rect 153670 657770 153910 658010
rect 154000 657770 154240 658010
rect 154330 657770 154570 658010
rect 154680 657770 154920 658010
rect 155010 657770 155250 658010
rect 155340 657770 155580 658010
rect 155670 657770 155910 658010
rect 144950 657420 145190 657660
rect 145300 657420 145540 657660
rect 145630 657420 145870 657660
rect 145960 657420 146200 657660
rect 146290 657420 146530 657660
rect 146640 657420 146880 657660
rect 146970 657420 147210 657660
rect 147300 657420 147540 657660
rect 147630 657420 147870 657660
rect 147980 657420 148220 657660
rect 148310 657420 148550 657660
rect 148640 657420 148880 657660
rect 148970 657420 149210 657660
rect 149320 657420 149560 657660
rect 149650 657420 149890 657660
rect 149980 657420 150220 657660
rect 150310 657420 150550 657660
rect 150660 657420 150900 657660
rect 150990 657420 151230 657660
rect 151320 657420 151560 657660
rect 151650 657420 151890 657660
rect 152000 657420 152240 657660
rect 152330 657420 152570 657660
rect 152660 657420 152900 657660
rect 152990 657420 153230 657660
rect 153340 657420 153580 657660
rect 153670 657420 153910 657660
rect 154000 657420 154240 657660
rect 154330 657420 154570 657660
rect 154680 657420 154920 657660
rect 155010 657420 155250 657660
rect 155340 657420 155580 657660
rect 155670 657420 155910 657660
rect 144950 657090 145190 657330
rect 145300 657090 145540 657330
rect 145630 657090 145870 657330
rect 145960 657090 146200 657330
rect 146290 657090 146530 657330
rect 146640 657090 146880 657330
rect 146970 657090 147210 657330
rect 147300 657090 147540 657330
rect 147630 657090 147870 657330
rect 147980 657090 148220 657330
rect 148310 657090 148550 657330
rect 148640 657090 148880 657330
rect 148970 657090 149210 657330
rect 149320 657090 149560 657330
rect 149650 657090 149890 657330
rect 149980 657090 150220 657330
rect 150310 657090 150550 657330
rect 150660 657090 150900 657330
rect 150990 657090 151230 657330
rect 151320 657090 151560 657330
rect 151650 657090 151890 657330
rect 152000 657090 152240 657330
rect 152330 657090 152570 657330
rect 152660 657090 152900 657330
rect 152990 657090 153230 657330
rect 153340 657090 153580 657330
rect 153670 657090 153910 657330
rect 154000 657090 154240 657330
rect 154330 657090 154570 657330
rect 154680 657090 154920 657330
rect 155010 657090 155250 657330
rect 155340 657090 155580 657330
rect 155670 657090 155910 657330
rect 144950 656760 145190 657000
rect 145300 656760 145540 657000
rect 145630 656760 145870 657000
rect 145960 656760 146200 657000
rect 146290 656760 146530 657000
rect 146640 656760 146880 657000
rect 146970 656760 147210 657000
rect 147300 656760 147540 657000
rect 147630 656760 147870 657000
rect 147980 656760 148220 657000
rect 148310 656760 148550 657000
rect 148640 656760 148880 657000
rect 148970 656760 149210 657000
rect 149320 656760 149560 657000
rect 149650 656760 149890 657000
rect 149980 656760 150220 657000
rect 150310 656760 150550 657000
rect 150660 656760 150900 657000
rect 150990 656760 151230 657000
rect 151320 656760 151560 657000
rect 151650 656760 151890 657000
rect 152000 656760 152240 657000
rect 152330 656760 152570 657000
rect 152660 656760 152900 657000
rect 152990 656760 153230 657000
rect 153340 656760 153580 657000
rect 153670 656760 153910 657000
rect 154000 656760 154240 657000
rect 154330 656760 154570 657000
rect 154680 656760 154920 657000
rect 155010 656760 155250 657000
rect 155340 656760 155580 657000
rect 155670 656760 155910 657000
rect 144950 656430 145190 656670
rect 145300 656430 145540 656670
rect 145630 656430 145870 656670
rect 145960 656430 146200 656670
rect 146290 656430 146530 656670
rect 146640 656430 146880 656670
rect 146970 656430 147210 656670
rect 147300 656430 147540 656670
rect 147630 656430 147870 656670
rect 147980 656430 148220 656670
rect 148310 656430 148550 656670
rect 148640 656430 148880 656670
rect 148970 656430 149210 656670
rect 149320 656430 149560 656670
rect 149650 656430 149890 656670
rect 149980 656430 150220 656670
rect 150310 656430 150550 656670
rect 150660 656430 150900 656670
rect 150990 656430 151230 656670
rect 151320 656430 151560 656670
rect 151650 656430 151890 656670
rect 152000 656430 152240 656670
rect 152330 656430 152570 656670
rect 152660 656430 152900 656670
rect 152990 656430 153230 656670
rect 153340 656430 153580 656670
rect 153670 656430 153910 656670
rect 154000 656430 154240 656670
rect 154330 656430 154570 656670
rect 154680 656430 154920 656670
rect 155010 656430 155250 656670
rect 155340 656430 155580 656670
rect 155670 656430 155910 656670
rect 144950 656080 145190 656320
rect 145300 656080 145540 656320
rect 145630 656080 145870 656320
rect 145960 656080 146200 656320
rect 146290 656080 146530 656320
rect 146640 656080 146880 656320
rect 146970 656080 147210 656320
rect 147300 656080 147540 656320
rect 147630 656080 147870 656320
rect 147980 656080 148220 656320
rect 148310 656080 148550 656320
rect 148640 656080 148880 656320
rect 148970 656080 149210 656320
rect 149320 656080 149560 656320
rect 149650 656080 149890 656320
rect 149980 656080 150220 656320
rect 150310 656080 150550 656320
rect 150660 656080 150900 656320
rect 150990 656080 151230 656320
rect 151320 656080 151560 656320
rect 151650 656080 151890 656320
rect 152000 656080 152240 656320
rect 152330 656080 152570 656320
rect 152660 656080 152900 656320
rect 152990 656080 153230 656320
rect 153340 656080 153580 656320
rect 153670 656080 153910 656320
rect 154000 656080 154240 656320
rect 154330 656080 154570 656320
rect 154680 656080 154920 656320
rect 155010 656080 155250 656320
rect 155340 656080 155580 656320
rect 155670 656080 155910 656320
rect 144950 655750 145190 655990
rect 145300 655750 145540 655990
rect 145630 655750 145870 655990
rect 145960 655750 146200 655990
rect 146290 655750 146530 655990
rect 146640 655750 146880 655990
rect 146970 655750 147210 655990
rect 147300 655750 147540 655990
rect 147630 655750 147870 655990
rect 147980 655750 148220 655990
rect 148310 655750 148550 655990
rect 148640 655750 148880 655990
rect 148970 655750 149210 655990
rect 149320 655750 149560 655990
rect 149650 655750 149890 655990
rect 149980 655750 150220 655990
rect 150310 655750 150550 655990
rect 150660 655750 150900 655990
rect 150990 655750 151230 655990
rect 151320 655750 151560 655990
rect 151650 655750 151890 655990
rect 152000 655750 152240 655990
rect 152330 655750 152570 655990
rect 152660 655750 152900 655990
rect 152990 655750 153230 655990
rect 153340 655750 153580 655990
rect 153670 655750 153910 655990
rect 154000 655750 154240 655990
rect 154330 655750 154570 655990
rect 154680 655750 154920 655990
rect 155010 655750 155250 655990
rect 155340 655750 155580 655990
rect 155670 655750 155910 655990
rect 144950 655420 145190 655660
rect 145300 655420 145540 655660
rect 145630 655420 145870 655660
rect 145960 655420 146200 655660
rect 146290 655420 146530 655660
rect 146640 655420 146880 655660
rect 146970 655420 147210 655660
rect 147300 655420 147540 655660
rect 147630 655420 147870 655660
rect 147980 655420 148220 655660
rect 148310 655420 148550 655660
rect 148640 655420 148880 655660
rect 148970 655420 149210 655660
rect 149320 655420 149560 655660
rect 149650 655420 149890 655660
rect 149980 655420 150220 655660
rect 150310 655420 150550 655660
rect 150660 655420 150900 655660
rect 150990 655420 151230 655660
rect 151320 655420 151560 655660
rect 151650 655420 151890 655660
rect 152000 655420 152240 655660
rect 152330 655420 152570 655660
rect 152660 655420 152900 655660
rect 152990 655420 153230 655660
rect 153340 655420 153580 655660
rect 153670 655420 153910 655660
rect 154000 655420 154240 655660
rect 154330 655420 154570 655660
rect 154680 655420 154920 655660
rect 155010 655420 155250 655660
rect 155340 655420 155580 655660
rect 155670 655420 155910 655660
rect 144950 655090 145190 655330
rect 145300 655090 145540 655330
rect 145630 655090 145870 655330
rect 145960 655090 146200 655330
rect 146290 655090 146530 655330
rect 146640 655090 146880 655330
rect 146970 655090 147210 655330
rect 147300 655090 147540 655330
rect 147630 655090 147870 655330
rect 147980 655090 148220 655330
rect 148310 655090 148550 655330
rect 148640 655090 148880 655330
rect 148970 655090 149210 655330
rect 149320 655090 149560 655330
rect 149650 655090 149890 655330
rect 149980 655090 150220 655330
rect 150310 655090 150550 655330
rect 150660 655090 150900 655330
rect 150990 655090 151230 655330
rect 151320 655090 151560 655330
rect 151650 655090 151890 655330
rect 152000 655090 152240 655330
rect 152330 655090 152570 655330
rect 152660 655090 152900 655330
rect 152990 655090 153230 655330
rect 153340 655090 153580 655330
rect 153670 655090 153910 655330
rect 154000 655090 154240 655330
rect 154330 655090 154570 655330
rect 154680 655090 154920 655330
rect 155010 655090 155250 655330
rect 155340 655090 155580 655330
rect 155670 655090 155910 655330
rect 144950 654740 145190 654980
rect 145300 654740 145540 654980
rect 145630 654740 145870 654980
rect 145960 654740 146200 654980
rect 146290 654740 146530 654980
rect 146640 654740 146880 654980
rect 146970 654740 147210 654980
rect 147300 654740 147540 654980
rect 147630 654740 147870 654980
rect 147980 654740 148220 654980
rect 148310 654740 148550 654980
rect 148640 654740 148880 654980
rect 148970 654740 149210 654980
rect 149320 654740 149560 654980
rect 149650 654740 149890 654980
rect 149980 654740 150220 654980
rect 150310 654740 150550 654980
rect 150660 654740 150900 654980
rect 150990 654740 151230 654980
rect 151320 654740 151560 654980
rect 151650 654740 151890 654980
rect 152000 654740 152240 654980
rect 152330 654740 152570 654980
rect 152660 654740 152900 654980
rect 152990 654740 153230 654980
rect 153340 654740 153580 654980
rect 153670 654740 153910 654980
rect 154000 654740 154240 654980
rect 154330 654740 154570 654980
rect 154680 654740 154920 654980
rect 155010 654740 155250 654980
rect 155340 654740 155580 654980
rect 155670 654740 155910 654980
rect 144950 654410 145190 654650
rect 145300 654410 145540 654650
rect 145630 654410 145870 654650
rect 145960 654410 146200 654650
rect 146290 654410 146530 654650
rect 146640 654410 146880 654650
rect 146970 654410 147210 654650
rect 147300 654410 147540 654650
rect 147630 654410 147870 654650
rect 147980 654410 148220 654650
rect 148310 654410 148550 654650
rect 148640 654410 148880 654650
rect 148970 654410 149210 654650
rect 149320 654410 149560 654650
rect 149650 654410 149890 654650
rect 149980 654410 150220 654650
rect 150310 654410 150550 654650
rect 150660 654410 150900 654650
rect 150990 654410 151230 654650
rect 151320 654410 151560 654650
rect 151650 654410 151890 654650
rect 152000 654410 152240 654650
rect 152330 654410 152570 654650
rect 152660 654410 152900 654650
rect 152990 654410 153230 654650
rect 153340 654410 153580 654650
rect 153670 654410 153910 654650
rect 154000 654410 154240 654650
rect 154330 654410 154570 654650
rect 154680 654410 154920 654650
rect 155010 654410 155250 654650
rect 155340 654410 155580 654650
rect 155670 654410 155910 654650
rect 144950 654080 145190 654320
rect 145300 654080 145540 654320
rect 145630 654080 145870 654320
rect 145960 654080 146200 654320
rect 146290 654080 146530 654320
rect 146640 654080 146880 654320
rect 146970 654080 147210 654320
rect 147300 654080 147540 654320
rect 147630 654080 147870 654320
rect 147980 654080 148220 654320
rect 148310 654080 148550 654320
rect 148640 654080 148880 654320
rect 148970 654080 149210 654320
rect 149320 654080 149560 654320
rect 149650 654080 149890 654320
rect 149980 654080 150220 654320
rect 150310 654080 150550 654320
rect 150660 654080 150900 654320
rect 150990 654080 151230 654320
rect 151320 654080 151560 654320
rect 151650 654080 151890 654320
rect 152000 654080 152240 654320
rect 152330 654080 152570 654320
rect 152660 654080 152900 654320
rect 152990 654080 153230 654320
rect 153340 654080 153580 654320
rect 153670 654080 153910 654320
rect 154000 654080 154240 654320
rect 154330 654080 154570 654320
rect 154680 654080 154920 654320
rect 155010 654080 155250 654320
rect 155340 654080 155580 654320
rect 155670 654080 155910 654320
rect 144950 653750 145190 653990
rect 145300 653750 145540 653990
rect 145630 653750 145870 653990
rect 145960 653750 146200 653990
rect 146290 653750 146530 653990
rect 146640 653750 146880 653990
rect 146970 653750 147210 653990
rect 147300 653750 147540 653990
rect 147630 653750 147870 653990
rect 147980 653750 148220 653990
rect 148310 653750 148550 653990
rect 148640 653750 148880 653990
rect 148970 653750 149210 653990
rect 149320 653750 149560 653990
rect 149650 653750 149890 653990
rect 149980 653750 150220 653990
rect 150310 653750 150550 653990
rect 150660 653750 150900 653990
rect 150990 653750 151230 653990
rect 151320 653750 151560 653990
rect 151650 653750 151890 653990
rect 152000 653750 152240 653990
rect 152330 653750 152570 653990
rect 152660 653750 152900 653990
rect 152990 653750 153230 653990
rect 153340 653750 153580 653990
rect 153670 653750 153910 653990
rect 154000 653750 154240 653990
rect 154330 653750 154570 653990
rect 154680 653750 154920 653990
rect 155010 653750 155250 653990
rect 155340 653750 155580 653990
rect 155670 653750 155910 653990
rect 144950 653400 145190 653640
rect 145300 653400 145540 653640
rect 145630 653400 145870 653640
rect 145960 653400 146200 653640
rect 146290 653400 146530 653640
rect 146640 653400 146880 653640
rect 146970 653400 147210 653640
rect 147300 653400 147540 653640
rect 147630 653400 147870 653640
rect 147980 653400 148220 653640
rect 148310 653400 148550 653640
rect 148640 653400 148880 653640
rect 148970 653400 149210 653640
rect 149320 653400 149560 653640
rect 149650 653400 149890 653640
rect 149980 653400 150220 653640
rect 150310 653400 150550 653640
rect 150660 653400 150900 653640
rect 150990 653400 151230 653640
rect 151320 653400 151560 653640
rect 151650 653400 151890 653640
rect 152000 653400 152240 653640
rect 152330 653400 152570 653640
rect 152660 653400 152900 653640
rect 152990 653400 153230 653640
rect 153340 653400 153580 653640
rect 153670 653400 153910 653640
rect 154000 653400 154240 653640
rect 154330 653400 154570 653640
rect 154680 653400 154920 653640
rect 155010 653400 155250 653640
rect 155340 653400 155580 653640
rect 155670 653400 155910 653640
rect 144950 653070 145190 653310
rect 145300 653070 145540 653310
rect 145630 653070 145870 653310
rect 145960 653070 146200 653310
rect 146290 653070 146530 653310
rect 146640 653070 146880 653310
rect 146970 653070 147210 653310
rect 147300 653070 147540 653310
rect 147630 653070 147870 653310
rect 147980 653070 148220 653310
rect 148310 653070 148550 653310
rect 148640 653070 148880 653310
rect 148970 653070 149210 653310
rect 149320 653070 149560 653310
rect 149650 653070 149890 653310
rect 149980 653070 150220 653310
rect 150310 653070 150550 653310
rect 150660 653070 150900 653310
rect 150990 653070 151230 653310
rect 151320 653070 151560 653310
rect 151650 653070 151890 653310
rect 152000 653070 152240 653310
rect 152330 653070 152570 653310
rect 152660 653070 152900 653310
rect 152990 653070 153230 653310
rect 153340 653070 153580 653310
rect 153670 653070 153910 653310
rect 154000 653070 154240 653310
rect 154330 653070 154570 653310
rect 154680 653070 154920 653310
rect 155010 653070 155250 653310
rect 155340 653070 155580 653310
rect 155670 653070 155910 653310
rect 144950 652740 145190 652980
rect 145300 652740 145540 652980
rect 145630 652740 145870 652980
rect 145960 652740 146200 652980
rect 146290 652740 146530 652980
rect 146640 652740 146880 652980
rect 146970 652740 147210 652980
rect 147300 652740 147540 652980
rect 147630 652740 147870 652980
rect 147980 652740 148220 652980
rect 148310 652740 148550 652980
rect 148640 652740 148880 652980
rect 148970 652740 149210 652980
rect 149320 652740 149560 652980
rect 149650 652740 149890 652980
rect 149980 652740 150220 652980
rect 150310 652740 150550 652980
rect 150660 652740 150900 652980
rect 150990 652740 151230 652980
rect 151320 652740 151560 652980
rect 151650 652740 151890 652980
rect 152000 652740 152240 652980
rect 152330 652740 152570 652980
rect 152660 652740 152900 652980
rect 152990 652740 153230 652980
rect 153340 652740 153580 652980
rect 153670 652740 153910 652980
rect 154000 652740 154240 652980
rect 154330 652740 154570 652980
rect 154680 652740 154920 652980
rect 155010 652740 155250 652980
rect 155340 652740 155580 652980
rect 155670 652740 155910 652980
rect 144950 652410 145190 652650
rect 145300 652410 145540 652650
rect 145630 652410 145870 652650
rect 145960 652410 146200 652650
rect 146290 652410 146530 652650
rect 146640 652410 146880 652650
rect 146970 652410 147210 652650
rect 147300 652410 147540 652650
rect 147630 652410 147870 652650
rect 147980 652410 148220 652650
rect 148310 652410 148550 652650
rect 148640 652410 148880 652650
rect 148970 652410 149210 652650
rect 149320 652410 149560 652650
rect 149650 652410 149890 652650
rect 149980 652410 150220 652650
rect 150310 652410 150550 652650
rect 150660 652410 150900 652650
rect 150990 652410 151230 652650
rect 151320 652410 151560 652650
rect 151650 652410 151890 652650
rect 152000 652410 152240 652650
rect 152330 652410 152570 652650
rect 152660 652410 152900 652650
rect 152990 652410 153230 652650
rect 153340 652410 153580 652650
rect 153670 652410 153910 652650
rect 154000 652410 154240 652650
rect 154330 652410 154570 652650
rect 154680 652410 154920 652650
rect 155010 652410 155250 652650
rect 155340 652410 155580 652650
rect 155670 652410 155910 652650
rect 144950 652060 145190 652300
rect 145300 652060 145540 652300
rect 145630 652060 145870 652300
rect 145960 652060 146200 652300
rect 146290 652060 146530 652300
rect 146640 652060 146880 652300
rect 146970 652060 147210 652300
rect 147300 652060 147540 652300
rect 147630 652060 147870 652300
rect 147980 652060 148220 652300
rect 148310 652060 148550 652300
rect 148640 652060 148880 652300
rect 148970 652060 149210 652300
rect 149320 652060 149560 652300
rect 149650 652060 149890 652300
rect 149980 652060 150220 652300
rect 150310 652060 150550 652300
rect 150660 652060 150900 652300
rect 150990 652060 151230 652300
rect 151320 652060 151560 652300
rect 151650 652060 151890 652300
rect 152000 652060 152240 652300
rect 152330 652060 152570 652300
rect 152660 652060 152900 652300
rect 152990 652060 153230 652300
rect 153340 652060 153580 652300
rect 153670 652060 153910 652300
rect 154000 652060 154240 652300
rect 154330 652060 154570 652300
rect 154680 652060 154920 652300
rect 155010 652060 155250 652300
rect 155340 652060 155580 652300
rect 155670 652060 155910 652300
rect 144950 651730 145190 651970
rect 145300 651730 145540 651970
rect 145630 651730 145870 651970
rect 145960 651730 146200 651970
rect 146290 651730 146530 651970
rect 146640 651730 146880 651970
rect 146970 651730 147210 651970
rect 147300 651730 147540 651970
rect 147630 651730 147870 651970
rect 147980 651730 148220 651970
rect 148310 651730 148550 651970
rect 148640 651730 148880 651970
rect 148970 651730 149210 651970
rect 149320 651730 149560 651970
rect 149650 651730 149890 651970
rect 149980 651730 150220 651970
rect 150310 651730 150550 651970
rect 150660 651730 150900 651970
rect 150990 651730 151230 651970
rect 151320 651730 151560 651970
rect 151650 651730 151890 651970
rect 152000 651730 152240 651970
rect 152330 651730 152570 651970
rect 152660 651730 152900 651970
rect 152990 651730 153230 651970
rect 153340 651730 153580 651970
rect 153670 651730 153910 651970
rect 154000 651730 154240 651970
rect 154330 651730 154570 651970
rect 154680 651730 154920 651970
rect 155010 651730 155250 651970
rect 155340 651730 155580 651970
rect 155670 651730 155910 651970
rect 144950 651400 145190 651640
rect 145300 651400 145540 651640
rect 145630 651400 145870 651640
rect 145960 651400 146200 651640
rect 146290 651400 146530 651640
rect 146640 651400 146880 651640
rect 146970 651400 147210 651640
rect 147300 651400 147540 651640
rect 147630 651400 147870 651640
rect 147980 651400 148220 651640
rect 148310 651400 148550 651640
rect 148640 651400 148880 651640
rect 148970 651400 149210 651640
rect 149320 651400 149560 651640
rect 149650 651400 149890 651640
rect 149980 651400 150220 651640
rect 150310 651400 150550 651640
rect 150660 651400 150900 651640
rect 150990 651400 151230 651640
rect 151320 651400 151560 651640
rect 151650 651400 151890 651640
rect 152000 651400 152240 651640
rect 152330 651400 152570 651640
rect 152660 651400 152900 651640
rect 152990 651400 153230 651640
rect 153340 651400 153580 651640
rect 153670 651400 153910 651640
rect 154000 651400 154240 651640
rect 154330 651400 154570 651640
rect 154680 651400 154920 651640
rect 155010 651400 155250 651640
rect 155340 651400 155580 651640
rect 155670 651400 155910 651640
rect 144950 651070 145190 651310
rect 145300 651070 145540 651310
rect 145630 651070 145870 651310
rect 145960 651070 146200 651310
rect 146290 651070 146530 651310
rect 146640 651070 146880 651310
rect 146970 651070 147210 651310
rect 147300 651070 147540 651310
rect 147630 651070 147870 651310
rect 147980 651070 148220 651310
rect 148310 651070 148550 651310
rect 148640 651070 148880 651310
rect 148970 651070 149210 651310
rect 149320 651070 149560 651310
rect 149650 651070 149890 651310
rect 149980 651070 150220 651310
rect 150310 651070 150550 651310
rect 150660 651070 150900 651310
rect 150990 651070 151230 651310
rect 151320 651070 151560 651310
rect 151650 651070 151890 651310
rect 152000 651070 152240 651310
rect 152330 651070 152570 651310
rect 152660 651070 152900 651310
rect 152990 651070 153230 651310
rect 153340 651070 153580 651310
rect 153670 651070 153910 651310
rect 154000 651070 154240 651310
rect 154330 651070 154570 651310
rect 154680 651070 154920 651310
rect 155010 651070 155250 651310
rect 155340 651070 155580 651310
rect 155670 651070 155910 651310
rect 144950 650720 145190 650960
rect 145300 650720 145540 650960
rect 145630 650720 145870 650960
rect 145960 650720 146200 650960
rect 146290 650720 146530 650960
rect 146640 650720 146880 650960
rect 146970 650720 147210 650960
rect 147300 650720 147540 650960
rect 147630 650720 147870 650960
rect 147980 650720 148220 650960
rect 148310 650720 148550 650960
rect 148640 650720 148880 650960
rect 148970 650720 149210 650960
rect 149320 650720 149560 650960
rect 149650 650720 149890 650960
rect 149980 650720 150220 650960
rect 150310 650720 150550 650960
rect 150660 650720 150900 650960
rect 150990 650720 151230 650960
rect 151320 650720 151560 650960
rect 151650 650720 151890 650960
rect 152000 650720 152240 650960
rect 152330 650720 152570 650960
rect 152660 650720 152900 650960
rect 152990 650720 153230 650960
rect 153340 650720 153580 650960
rect 153670 650720 153910 650960
rect 154000 650720 154240 650960
rect 154330 650720 154570 650960
rect 154680 650720 154920 650960
rect 155010 650720 155250 650960
rect 155340 650720 155580 650960
rect 155670 650720 155910 650960
rect 144950 650390 145190 650630
rect 145300 650390 145540 650630
rect 145630 650390 145870 650630
rect 145960 650390 146200 650630
rect 146290 650390 146530 650630
rect 146640 650390 146880 650630
rect 146970 650390 147210 650630
rect 147300 650390 147540 650630
rect 147630 650390 147870 650630
rect 147980 650390 148220 650630
rect 148310 650390 148550 650630
rect 148640 650390 148880 650630
rect 148970 650390 149210 650630
rect 149320 650390 149560 650630
rect 149650 650390 149890 650630
rect 149980 650390 150220 650630
rect 150310 650390 150550 650630
rect 150660 650390 150900 650630
rect 150990 650390 151230 650630
rect 151320 650390 151560 650630
rect 151650 650390 151890 650630
rect 152000 650390 152240 650630
rect 152330 650390 152570 650630
rect 152660 650390 152900 650630
rect 152990 650390 153230 650630
rect 153340 650390 153580 650630
rect 153670 650390 153910 650630
rect 154000 650390 154240 650630
rect 154330 650390 154570 650630
rect 154680 650390 154920 650630
rect 155010 650390 155250 650630
rect 155340 650390 155580 650630
rect 155670 650390 155910 650630
rect 144950 650060 145190 650300
rect 145300 650060 145540 650300
rect 145630 650060 145870 650300
rect 145960 650060 146200 650300
rect 146290 650060 146530 650300
rect 146640 650060 146880 650300
rect 146970 650060 147210 650300
rect 147300 650060 147540 650300
rect 147630 650060 147870 650300
rect 147980 650060 148220 650300
rect 148310 650060 148550 650300
rect 148640 650060 148880 650300
rect 148970 650060 149210 650300
rect 149320 650060 149560 650300
rect 149650 650060 149890 650300
rect 149980 650060 150220 650300
rect 150310 650060 150550 650300
rect 150660 650060 150900 650300
rect 150990 650060 151230 650300
rect 151320 650060 151560 650300
rect 151650 650060 151890 650300
rect 152000 650060 152240 650300
rect 152330 650060 152570 650300
rect 152660 650060 152900 650300
rect 152990 650060 153230 650300
rect 153340 650060 153580 650300
rect 153670 650060 153910 650300
rect 154000 650060 154240 650300
rect 154330 650060 154570 650300
rect 154680 650060 154920 650300
rect 155010 650060 155250 650300
rect 155340 650060 155580 650300
rect 155670 650060 155910 650300
rect 144950 649730 145190 649970
rect 145300 649730 145540 649970
rect 145630 649730 145870 649970
rect 145960 649730 146200 649970
rect 146290 649730 146530 649970
rect 146640 649730 146880 649970
rect 146970 649730 147210 649970
rect 147300 649730 147540 649970
rect 147630 649730 147870 649970
rect 147980 649730 148220 649970
rect 148310 649730 148550 649970
rect 148640 649730 148880 649970
rect 148970 649730 149210 649970
rect 149320 649730 149560 649970
rect 149650 649730 149890 649970
rect 149980 649730 150220 649970
rect 150310 649730 150550 649970
rect 150660 649730 150900 649970
rect 150990 649730 151230 649970
rect 151320 649730 151560 649970
rect 151650 649730 151890 649970
rect 152000 649730 152240 649970
rect 152330 649730 152570 649970
rect 152660 649730 152900 649970
rect 152990 649730 153230 649970
rect 153340 649730 153580 649970
rect 153670 649730 153910 649970
rect 154000 649730 154240 649970
rect 154330 649730 154570 649970
rect 154680 649730 154920 649970
rect 155010 649730 155250 649970
rect 155340 649730 155580 649970
rect 155670 649730 155910 649970
rect 144950 649380 145190 649620
rect 145300 649380 145540 649620
rect 145630 649380 145870 649620
rect 145960 649380 146200 649620
rect 146290 649380 146530 649620
rect 146640 649380 146880 649620
rect 146970 649380 147210 649620
rect 147300 649380 147540 649620
rect 147630 649380 147870 649620
rect 147980 649380 148220 649620
rect 148310 649380 148550 649620
rect 148640 649380 148880 649620
rect 148970 649380 149210 649620
rect 149320 649380 149560 649620
rect 149650 649380 149890 649620
rect 149980 649380 150220 649620
rect 150310 649380 150550 649620
rect 150660 649380 150900 649620
rect 150990 649380 151230 649620
rect 151320 649380 151560 649620
rect 151650 649380 151890 649620
rect 152000 649380 152240 649620
rect 152330 649380 152570 649620
rect 152660 649380 152900 649620
rect 152990 649380 153230 649620
rect 153340 649380 153580 649620
rect 153670 649380 153910 649620
rect 154000 649380 154240 649620
rect 154330 649380 154570 649620
rect 154680 649380 154920 649620
rect 155010 649380 155250 649620
rect 155340 649380 155580 649620
rect 155670 649380 155910 649620
<< metal5 >>
rect 16194 703800 21194 704000
rect 16194 703500 16352 703800
rect 16652 703500 16852 703800
rect 17152 703500 17352 703800
rect 17652 703500 17852 703800
rect 18152 703500 18352 703800
rect 18652 703500 18852 703800
rect 19152 703500 19352 703800
rect 19652 703500 19852 703800
rect 20152 703500 20352 703800
rect 20652 703500 20852 703800
rect 21152 703500 21194 703800
rect 16194 703300 21194 703500
rect 16194 703000 16352 703300
rect 16652 703000 16852 703300
rect 17152 703000 17352 703300
rect 17652 703000 17852 703300
rect 18152 703000 18352 703300
rect 18652 703000 18852 703300
rect 19152 703000 19352 703300
rect 19652 703000 19852 703300
rect 20152 703000 20352 703300
rect 20652 703000 20852 703300
rect 21152 703000 21194 703300
rect 16194 702800 21194 703000
rect 16194 702500 16352 702800
rect 16652 702500 16852 702800
rect 17152 702500 17352 702800
rect 17652 702500 17852 702800
rect 18152 702500 18352 702800
rect 18652 702500 18852 702800
rect 19152 702500 19352 702800
rect 19652 702500 19852 702800
rect 20152 702500 20352 702800
rect 20652 702500 20852 702800
rect 21152 702500 21194 702800
rect 16194 697044 21194 702500
rect 165594 702300 170594 704800
rect 0 685237 2500 685242
rect 0 685200 7495 685237
rect 0 684900 200 685200
rect 500 684900 700 685200
rect 1000 684900 1200 685200
rect 1500 684900 7495 685200
rect 0 684700 7495 684900
rect 0 684400 200 684700
rect 500 684400 700 684700
rect 1000 684400 1200 684700
rect 1500 684400 7495 684700
rect 0 684200 7495 684400
rect 0 683900 200 684200
rect 500 683900 700 684200
rect 1000 683900 1200 684200
rect 1500 683900 7495 684200
rect 0 683700 7495 683900
rect 0 683400 200 683700
rect 500 683400 700 683700
rect 1000 683400 1200 683700
rect 1500 683400 7495 683700
rect 0 683200 7495 683400
rect 0 682900 200 683200
rect 500 682900 700 683200
rect 1000 682900 1200 683200
rect 1500 682900 7495 683200
rect 0 682700 7495 682900
rect 0 682400 200 682700
rect 500 682400 700 682700
rect 1000 682400 1200 682700
rect 1500 682400 7495 682700
rect 0 682200 7495 682400
rect 0 681900 200 682200
rect 500 681900 700 682200
rect 1000 681900 1200 682200
rect 1500 681900 7495 682200
rect 0 681700 7495 681900
rect 0 681400 200 681700
rect 500 681400 700 681700
rect 1000 681400 1200 681700
rect 1500 681400 7495 681700
rect 0 681200 7495 681400
rect 0 680900 200 681200
rect 500 680900 700 681200
rect 1000 680900 1200 681200
rect 1500 680900 7495 681200
rect 0 680700 7495 680900
rect 0 680400 200 680700
rect 500 680400 700 680700
rect 1000 680400 1200 680700
rect 1500 680400 7495 680700
rect 0 680242 7495 680400
rect 2500 665500 7495 680242
rect 16197 679147 21192 697044
rect 110760 694840 155960 694890
rect 110760 694600 110810 694840
rect 111050 694600 111140 694840
rect 111380 694600 111470 694840
rect 111710 694600 111800 694840
rect 112040 694600 112150 694840
rect 112390 694600 112480 694840
rect 112720 694600 112810 694840
rect 113050 694600 113140 694840
rect 113380 694600 113490 694840
rect 113730 694600 113820 694840
rect 114060 694600 114150 694840
rect 114390 694600 114480 694840
rect 114720 694600 114830 694840
rect 115070 694600 115160 694840
rect 115400 694600 115490 694840
rect 115730 694600 115820 694840
rect 116060 694600 116170 694840
rect 116410 694600 116500 694840
rect 116740 694600 116830 694840
rect 117070 694600 117160 694840
rect 117400 694600 117510 694840
rect 117750 694600 117840 694840
rect 118080 694600 118170 694840
rect 118410 694600 118500 694840
rect 118740 694600 118850 694840
rect 119090 694600 119180 694840
rect 119420 694600 119510 694840
rect 119750 694600 119840 694840
rect 120080 694600 120190 694840
rect 120430 694600 120520 694840
rect 120760 694600 120850 694840
rect 121090 694600 121180 694840
rect 121420 694600 121530 694840
rect 121770 694600 122190 694840
rect 122430 694600 122520 694840
rect 122760 694600 122850 694840
rect 123090 694600 123180 694840
rect 123420 694600 123530 694840
rect 123770 694600 123860 694840
rect 124100 694600 124190 694840
rect 124430 694600 124520 694840
rect 124760 694600 124870 694840
rect 125110 694600 125200 694840
rect 125440 694600 125530 694840
rect 125770 694600 125860 694840
rect 126100 694600 126210 694840
rect 126450 694600 126540 694840
rect 126780 694600 126870 694840
rect 127110 694600 127200 694840
rect 127440 694600 127550 694840
rect 127790 694600 127880 694840
rect 128120 694600 128210 694840
rect 128450 694600 128540 694840
rect 128780 694600 128890 694840
rect 129130 694600 129220 694840
rect 129460 694600 129550 694840
rect 129790 694600 129880 694840
rect 130120 694600 130230 694840
rect 130470 694600 130560 694840
rect 130800 694600 130890 694840
rect 131130 694600 131220 694840
rect 131460 694600 131570 694840
rect 131810 694600 131900 694840
rect 132140 694600 132230 694840
rect 132470 694600 132560 694840
rect 132800 694600 132910 694840
rect 133150 694600 133570 694840
rect 133810 694600 133900 694840
rect 134140 694600 134230 694840
rect 134470 694600 134560 694840
rect 134800 694600 134910 694840
rect 135150 694600 135240 694840
rect 135480 694600 135570 694840
rect 135810 694600 135900 694840
rect 136140 694600 136250 694840
rect 136490 694600 136580 694840
rect 136820 694600 136910 694840
rect 137150 694600 137240 694840
rect 137480 694600 137590 694840
rect 137830 694600 137920 694840
rect 138160 694600 138250 694840
rect 138490 694600 138580 694840
rect 138820 694600 138930 694840
rect 139170 694600 139260 694840
rect 139500 694600 139590 694840
rect 139830 694600 139920 694840
rect 140160 694600 140270 694840
rect 140510 694600 140600 694840
rect 140840 694600 140930 694840
rect 141170 694600 141260 694840
rect 141500 694600 141610 694840
rect 141850 694600 141940 694840
rect 142180 694600 142270 694840
rect 142510 694600 142600 694840
rect 142840 694600 142950 694840
rect 143190 694600 143280 694840
rect 143520 694600 143610 694840
rect 143850 694600 143940 694840
rect 144180 694600 144290 694840
rect 144530 694600 144950 694840
rect 145190 694600 145280 694840
rect 145520 694600 145610 694840
rect 145850 694600 145940 694840
rect 146180 694600 146290 694840
rect 146530 694600 146620 694840
rect 146860 694600 146950 694840
rect 147190 694600 147280 694840
rect 147520 694600 147630 694840
rect 147870 694600 147960 694840
rect 148200 694600 148290 694840
rect 148530 694600 148620 694840
rect 148860 694600 148970 694840
rect 149210 694600 149300 694840
rect 149540 694600 149630 694840
rect 149870 694600 149960 694840
rect 150200 694600 150310 694840
rect 150550 694600 150640 694840
rect 150880 694600 150970 694840
rect 151210 694600 151300 694840
rect 151540 694600 151650 694840
rect 151890 694600 151980 694840
rect 152220 694600 152310 694840
rect 152550 694600 152640 694840
rect 152880 694600 152990 694840
rect 153230 694600 153320 694840
rect 153560 694600 153650 694840
rect 153890 694600 153980 694840
rect 154220 694600 154330 694840
rect 154570 694600 154660 694840
rect 154900 694600 154990 694840
rect 155230 694600 155320 694840
rect 155560 694600 155670 694840
rect 155910 694600 155960 694840
rect 110760 694490 155960 694600
rect 110760 694250 110810 694490
rect 111050 694250 111140 694490
rect 111380 694250 111470 694490
rect 111710 694250 111800 694490
rect 112040 694250 112150 694490
rect 112390 694250 112480 694490
rect 112720 694250 112810 694490
rect 113050 694250 113140 694490
rect 113380 694250 113490 694490
rect 113730 694250 113820 694490
rect 114060 694250 114150 694490
rect 114390 694250 114480 694490
rect 114720 694250 114830 694490
rect 115070 694250 115160 694490
rect 115400 694250 115490 694490
rect 115730 694250 115820 694490
rect 116060 694250 116170 694490
rect 116410 694250 116500 694490
rect 116740 694250 116830 694490
rect 117070 694250 117160 694490
rect 117400 694250 117510 694490
rect 117750 694250 117840 694490
rect 118080 694250 118170 694490
rect 118410 694250 118500 694490
rect 118740 694250 118850 694490
rect 119090 694250 119180 694490
rect 119420 694250 119510 694490
rect 119750 694250 119840 694490
rect 120080 694250 120190 694490
rect 120430 694250 120520 694490
rect 120760 694250 120850 694490
rect 121090 694250 121180 694490
rect 121420 694250 121530 694490
rect 121770 694250 122190 694490
rect 122430 694250 122520 694490
rect 122760 694250 122850 694490
rect 123090 694250 123180 694490
rect 123420 694250 123530 694490
rect 123770 694250 123860 694490
rect 124100 694250 124190 694490
rect 124430 694250 124520 694490
rect 124760 694250 124870 694490
rect 125110 694250 125200 694490
rect 125440 694250 125530 694490
rect 125770 694250 125860 694490
rect 126100 694250 126210 694490
rect 126450 694250 126540 694490
rect 126780 694250 126870 694490
rect 127110 694250 127200 694490
rect 127440 694250 127550 694490
rect 127790 694250 127880 694490
rect 128120 694250 128210 694490
rect 128450 694250 128540 694490
rect 128780 694250 128890 694490
rect 129130 694250 129220 694490
rect 129460 694250 129550 694490
rect 129790 694250 129880 694490
rect 130120 694250 130230 694490
rect 130470 694250 130560 694490
rect 130800 694250 130890 694490
rect 131130 694250 131220 694490
rect 131460 694250 131570 694490
rect 131810 694250 131900 694490
rect 132140 694250 132230 694490
rect 132470 694250 132560 694490
rect 132800 694250 132910 694490
rect 133150 694250 133570 694490
rect 133810 694250 133900 694490
rect 134140 694250 134230 694490
rect 134470 694250 134560 694490
rect 134800 694250 134910 694490
rect 135150 694250 135240 694490
rect 135480 694250 135570 694490
rect 135810 694250 135900 694490
rect 136140 694250 136250 694490
rect 136490 694250 136580 694490
rect 136820 694250 136910 694490
rect 137150 694250 137240 694490
rect 137480 694250 137590 694490
rect 137830 694250 137920 694490
rect 138160 694250 138250 694490
rect 138490 694250 138580 694490
rect 138820 694250 138930 694490
rect 139170 694250 139260 694490
rect 139500 694250 139590 694490
rect 139830 694250 139920 694490
rect 140160 694250 140270 694490
rect 140510 694250 140600 694490
rect 140840 694250 140930 694490
rect 141170 694250 141260 694490
rect 141500 694250 141610 694490
rect 141850 694250 141940 694490
rect 142180 694250 142270 694490
rect 142510 694250 142600 694490
rect 142840 694250 142950 694490
rect 143190 694250 143280 694490
rect 143520 694250 143610 694490
rect 143850 694250 143940 694490
rect 144180 694250 144290 694490
rect 144530 694250 144950 694490
rect 145190 694250 145280 694490
rect 145520 694250 145610 694490
rect 145850 694250 145940 694490
rect 146180 694250 146290 694490
rect 146530 694250 146620 694490
rect 146860 694250 146950 694490
rect 147190 694250 147280 694490
rect 147520 694250 147630 694490
rect 147870 694250 147960 694490
rect 148200 694250 148290 694490
rect 148530 694250 148620 694490
rect 148860 694250 148970 694490
rect 149210 694250 149300 694490
rect 149540 694250 149630 694490
rect 149870 694250 149960 694490
rect 150200 694250 150310 694490
rect 150550 694250 150640 694490
rect 150880 694250 150970 694490
rect 151210 694250 151300 694490
rect 151540 694250 151650 694490
rect 151890 694250 151980 694490
rect 152220 694250 152310 694490
rect 152550 694250 152640 694490
rect 152880 694250 152990 694490
rect 153230 694250 153320 694490
rect 153560 694250 153650 694490
rect 153890 694250 153980 694490
rect 154220 694250 154330 694490
rect 154570 694250 154660 694490
rect 154900 694250 154990 694490
rect 155230 694250 155320 694490
rect 155560 694250 155670 694490
rect 155910 694250 155960 694490
rect 110760 694160 155960 694250
rect 110760 693920 110810 694160
rect 111050 693920 111140 694160
rect 111380 693920 111470 694160
rect 111710 693920 111800 694160
rect 112040 693920 112150 694160
rect 112390 693920 112480 694160
rect 112720 693920 112810 694160
rect 113050 693920 113140 694160
rect 113380 693920 113490 694160
rect 113730 693920 113820 694160
rect 114060 693920 114150 694160
rect 114390 693920 114480 694160
rect 114720 693920 114830 694160
rect 115070 693920 115160 694160
rect 115400 693920 115490 694160
rect 115730 693920 115820 694160
rect 116060 693920 116170 694160
rect 116410 693920 116500 694160
rect 116740 693920 116830 694160
rect 117070 693920 117160 694160
rect 117400 693920 117510 694160
rect 117750 693920 117840 694160
rect 118080 693920 118170 694160
rect 118410 693920 118500 694160
rect 118740 693920 118850 694160
rect 119090 693920 119180 694160
rect 119420 693920 119510 694160
rect 119750 693920 119840 694160
rect 120080 693920 120190 694160
rect 120430 693920 120520 694160
rect 120760 693920 120850 694160
rect 121090 693920 121180 694160
rect 121420 693920 121530 694160
rect 121770 693920 122190 694160
rect 122430 693920 122520 694160
rect 122760 693920 122850 694160
rect 123090 693920 123180 694160
rect 123420 693920 123530 694160
rect 123770 693920 123860 694160
rect 124100 693920 124190 694160
rect 124430 693920 124520 694160
rect 124760 693920 124870 694160
rect 125110 693920 125200 694160
rect 125440 693920 125530 694160
rect 125770 693920 125860 694160
rect 126100 693920 126210 694160
rect 126450 693920 126540 694160
rect 126780 693920 126870 694160
rect 127110 693920 127200 694160
rect 127440 693920 127550 694160
rect 127790 693920 127880 694160
rect 128120 693920 128210 694160
rect 128450 693920 128540 694160
rect 128780 693920 128890 694160
rect 129130 693920 129220 694160
rect 129460 693920 129550 694160
rect 129790 693920 129880 694160
rect 130120 693920 130230 694160
rect 130470 693920 130560 694160
rect 130800 693920 130890 694160
rect 131130 693920 131220 694160
rect 131460 693920 131570 694160
rect 131810 693920 131900 694160
rect 132140 693920 132230 694160
rect 132470 693920 132560 694160
rect 132800 693920 132910 694160
rect 133150 693920 133570 694160
rect 133810 693920 133900 694160
rect 134140 693920 134230 694160
rect 134470 693920 134560 694160
rect 134800 693920 134910 694160
rect 135150 693920 135240 694160
rect 135480 693920 135570 694160
rect 135810 693920 135900 694160
rect 136140 693920 136250 694160
rect 136490 693920 136580 694160
rect 136820 693920 136910 694160
rect 137150 693920 137240 694160
rect 137480 693920 137590 694160
rect 137830 693920 137920 694160
rect 138160 693920 138250 694160
rect 138490 693920 138580 694160
rect 138820 693920 138930 694160
rect 139170 693920 139260 694160
rect 139500 693920 139590 694160
rect 139830 693920 139920 694160
rect 140160 693920 140270 694160
rect 140510 693920 140600 694160
rect 140840 693920 140930 694160
rect 141170 693920 141260 694160
rect 141500 693920 141610 694160
rect 141850 693920 141940 694160
rect 142180 693920 142270 694160
rect 142510 693920 142600 694160
rect 142840 693920 142950 694160
rect 143190 693920 143280 694160
rect 143520 693920 143610 694160
rect 143850 693920 143940 694160
rect 144180 693920 144290 694160
rect 144530 693920 144950 694160
rect 145190 693920 145280 694160
rect 145520 693920 145610 694160
rect 145850 693920 145940 694160
rect 146180 693920 146290 694160
rect 146530 693920 146620 694160
rect 146860 693920 146950 694160
rect 147190 693920 147280 694160
rect 147520 693920 147630 694160
rect 147870 693920 147960 694160
rect 148200 693920 148290 694160
rect 148530 693920 148620 694160
rect 148860 693920 148970 694160
rect 149210 693920 149300 694160
rect 149540 693920 149630 694160
rect 149870 693920 149960 694160
rect 150200 693920 150310 694160
rect 150550 693920 150640 694160
rect 150880 693920 150970 694160
rect 151210 693920 151300 694160
rect 151540 693920 151650 694160
rect 151890 693920 151980 694160
rect 152220 693920 152310 694160
rect 152550 693920 152640 694160
rect 152880 693920 152990 694160
rect 153230 693920 153320 694160
rect 153560 693920 153650 694160
rect 153890 693920 153980 694160
rect 154220 693920 154330 694160
rect 154570 693920 154660 694160
rect 154900 693920 154990 694160
rect 155230 693920 155320 694160
rect 155560 693920 155670 694160
rect 155910 693920 155960 694160
rect 110760 693830 155960 693920
rect 110760 693590 110810 693830
rect 111050 693590 111140 693830
rect 111380 693590 111470 693830
rect 111710 693590 111800 693830
rect 112040 693590 112150 693830
rect 112390 693590 112480 693830
rect 112720 693590 112810 693830
rect 113050 693590 113140 693830
rect 113380 693590 113490 693830
rect 113730 693590 113820 693830
rect 114060 693590 114150 693830
rect 114390 693590 114480 693830
rect 114720 693590 114830 693830
rect 115070 693590 115160 693830
rect 115400 693590 115490 693830
rect 115730 693590 115820 693830
rect 116060 693590 116170 693830
rect 116410 693590 116500 693830
rect 116740 693590 116830 693830
rect 117070 693590 117160 693830
rect 117400 693590 117510 693830
rect 117750 693590 117840 693830
rect 118080 693590 118170 693830
rect 118410 693590 118500 693830
rect 118740 693590 118850 693830
rect 119090 693590 119180 693830
rect 119420 693590 119510 693830
rect 119750 693590 119840 693830
rect 120080 693590 120190 693830
rect 120430 693590 120520 693830
rect 120760 693590 120850 693830
rect 121090 693590 121180 693830
rect 121420 693590 121530 693830
rect 121770 693590 122190 693830
rect 122430 693590 122520 693830
rect 122760 693590 122850 693830
rect 123090 693590 123180 693830
rect 123420 693590 123530 693830
rect 123770 693590 123860 693830
rect 124100 693590 124190 693830
rect 124430 693590 124520 693830
rect 124760 693590 124870 693830
rect 125110 693590 125200 693830
rect 125440 693590 125530 693830
rect 125770 693590 125860 693830
rect 126100 693590 126210 693830
rect 126450 693590 126540 693830
rect 126780 693590 126870 693830
rect 127110 693590 127200 693830
rect 127440 693590 127550 693830
rect 127790 693590 127880 693830
rect 128120 693590 128210 693830
rect 128450 693590 128540 693830
rect 128780 693590 128890 693830
rect 129130 693590 129220 693830
rect 129460 693590 129550 693830
rect 129790 693590 129880 693830
rect 130120 693590 130230 693830
rect 130470 693590 130560 693830
rect 130800 693590 130890 693830
rect 131130 693590 131220 693830
rect 131460 693590 131570 693830
rect 131810 693590 131900 693830
rect 132140 693590 132230 693830
rect 132470 693590 132560 693830
rect 132800 693590 132910 693830
rect 133150 693590 133570 693830
rect 133810 693590 133900 693830
rect 134140 693590 134230 693830
rect 134470 693590 134560 693830
rect 134800 693590 134910 693830
rect 135150 693590 135240 693830
rect 135480 693590 135570 693830
rect 135810 693590 135900 693830
rect 136140 693590 136250 693830
rect 136490 693590 136580 693830
rect 136820 693590 136910 693830
rect 137150 693590 137240 693830
rect 137480 693590 137590 693830
rect 137830 693590 137920 693830
rect 138160 693590 138250 693830
rect 138490 693590 138580 693830
rect 138820 693590 138930 693830
rect 139170 693590 139260 693830
rect 139500 693590 139590 693830
rect 139830 693590 139920 693830
rect 140160 693590 140270 693830
rect 140510 693590 140600 693830
rect 140840 693590 140930 693830
rect 141170 693590 141260 693830
rect 141500 693590 141610 693830
rect 141850 693590 141940 693830
rect 142180 693590 142270 693830
rect 142510 693590 142600 693830
rect 142840 693590 142950 693830
rect 143190 693590 143280 693830
rect 143520 693590 143610 693830
rect 143850 693590 143940 693830
rect 144180 693590 144290 693830
rect 144530 693590 144950 693830
rect 145190 693590 145280 693830
rect 145520 693590 145610 693830
rect 145850 693590 145940 693830
rect 146180 693590 146290 693830
rect 146530 693590 146620 693830
rect 146860 693590 146950 693830
rect 147190 693590 147280 693830
rect 147520 693590 147630 693830
rect 147870 693590 147960 693830
rect 148200 693590 148290 693830
rect 148530 693590 148620 693830
rect 148860 693590 148970 693830
rect 149210 693590 149300 693830
rect 149540 693590 149630 693830
rect 149870 693590 149960 693830
rect 150200 693590 150310 693830
rect 150550 693590 150640 693830
rect 150880 693590 150970 693830
rect 151210 693590 151300 693830
rect 151540 693590 151650 693830
rect 151890 693590 151980 693830
rect 152220 693590 152310 693830
rect 152550 693590 152640 693830
rect 152880 693590 152990 693830
rect 153230 693590 153320 693830
rect 153560 693590 153650 693830
rect 153890 693590 153980 693830
rect 154220 693590 154330 693830
rect 154570 693590 154660 693830
rect 154900 693590 154990 693830
rect 155230 693590 155320 693830
rect 155560 693590 155670 693830
rect 155910 693590 155960 693830
rect 110760 693500 155960 693590
rect 110760 693260 110810 693500
rect 111050 693260 111140 693500
rect 111380 693260 111470 693500
rect 111710 693260 111800 693500
rect 112040 693260 112150 693500
rect 112390 693260 112480 693500
rect 112720 693260 112810 693500
rect 113050 693260 113140 693500
rect 113380 693260 113490 693500
rect 113730 693260 113820 693500
rect 114060 693260 114150 693500
rect 114390 693260 114480 693500
rect 114720 693260 114830 693500
rect 115070 693260 115160 693500
rect 115400 693260 115490 693500
rect 115730 693260 115820 693500
rect 116060 693260 116170 693500
rect 116410 693260 116500 693500
rect 116740 693260 116830 693500
rect 117070 693260 117160 693500
rect 117400 693260 117510 693500
rect 117750 693260 117840 693500
rect 118080 693260 118170 693500
rect 118410 693260 118500 693500
rect 118740 693260 118850 693500
rect 119090 693260 119180 693500
rect 119420 693260 119510 693500
rect 119750 693260 119840 693500
rect 120080 693260 120190 693500
rect 120430 693260 120520 693500
rect 120760 693260 120850 693500
rect 121090 693260 121180 693500
rect 121420 693260 121530 693500
rect 121770 693260 122190 693500
rect 122430 693260 122520 693500
rect 122760 693260 122850 693500
rect 123090 693260 123180 693500
rect 123420 693260 123530 693500
rect 123770 693260 123860 693500
rect 124100 693260 124190 693500
rect 124430 693260 124520 693500
rect 124760 693260 124870 693500
rect 125110 693260 125200 693500
rect 125440 693260 125530 693500
rect 125770 693260 125860 693500
rect 126100 693260 126210 693500
rect 126450 693260 126540 693500
rect 126780 693260 126870 693500
rect 127110 693260 127200 693500
rect 127440 693260 127550 693500
rect 127790 693260 127880 693500
rect 128120 693260 128210 693500
rect 128450 693260 128540 693500
rect 128780 693260 128890 693500
rect 129130 693260 129220 693500
rect 129460 693260 129550 693500
rect 129790 693260 129880 693500
rect 130120 693260 130230 693500
rect 130470 693260 130560 693500
rect 130800 693260 130890 693500
rect 131130 693260 131220 693500
rect 131460 693260 131570 693500
rect 131810 693260 131900 693500
rect 132140 693260 132230 693500
rect 132470 693260 132560 693500
rect 132800 693260 132910 693500
rect 133150 693260 133570 693500
rect 133810 693260 133900 693500
rect 134140 693260 134230 693500
rect 134470 693260 134560 693500
rect 134800 693260 134910 693500
rect 135150 693260 135240 693500
rect 135480 693260 135570 693500
rect 135810 693260 135900 693500
rect 136140 693260 136250 693500
rect 136490 693260 136580 693500
rect 136820 693260 136910 693500
rect 137150 693260 137240 693500
rect 137480 693260 137590 693500
rect 137830 693260 137920 693500
rect 138160 693260 138250 693500
rect 138490 693260 138580 693500
rect 138820 693260 138930 693500
rect 139170 693260 139260 693500
rect 139500 693260 139590 693500
rect 139830 693260 139920 693500
rect 140160 693260 140270 693500
rect 140510 693260 140600 693500
rect 140840 693260 140930 693500
rect 141170 693260 141260 693500
rect 141500 693260 141610 693500
rect 141850 693260 141940 693500
rect 142180 693260 142270 693500
rect 142510 693260 142600 693500
rect 142840 693260 142950 693500
rect 143190 693260 143280 693500
rect 143520 693260 143610 693500
rect 143850 693260 143940 693500
rect 144180 693260 144290 693500
rect 144530 693260 144950 693500
rect 145190 693260 145280 693500
rect 145520 693260 145610 693500
rect 145850 693260 145940 693500
rect 146180 693260 146290 693500
rect 146530 693260 146620 693500
rect 146860 693260 146950 693500
rect 147190 693260 147280 693500
rect 147520 693260 147630 693500
rect 147870 693260 147960 693500
rect 148200 693260 148290 693500
rect 148530 693260 148620 693500
rect 148860 693260 148970 693500
rect 149210 693260 149300 693500
rect 149540 693260 149630 693500
rect 149870 693260 149960 693500
rect 150200 693260 150310 693500
rect 150550 693260 150640 693500
rect 150880 693260 150970 693500
rect 151210 693260 151300 693500
rect 151540 693260 151650 693500
rect 151890 693260 151980 693500
rect 152220 693260 152310 693500
rect 152550 693260 152640 693500
rect 152880 693260 152990 693500
rect 153230 693260 153320 693500
rect 153560 693260 153650 693500
rect 153890 693260 153980 693500
rect 154220 693260 154330 693500
rect 154570 693260 154660 693500
rect 154900 693260 154990 693500
rect 155230 693260 155320 693500
rect 155560 693260 155670 693500
rect 155910 693260 155960 693500
rect 110760 693150 155960 693260
rect 110760 692910 110810 693150
rect 111050 692910 111140 693150
rect 111380 692910 111470 693150
rect 111710 692910 111800 693150
rect 112040 692910 112150 693150
rect 112390 692910 112480 693150
rect 112720 692910 112810 693150
rect 113050 692910 113140 693150
rect 113380 692910 113490 693150
rect 113730 692910 113820 693150
rect 114060 692910 114150 693150
rect 114390 692910 114480 693150
rect 114720 692910 114830 693150
rect 115070 692910 115160 693150
rect 115400 692910 115490 693150
rect 115730 692910 115820 693150
rect 116060 692910 116170 693150
rect 116410 692910 116500 693150
rect 116740 692910 116830 693150
rect 117070 692910 117160 693150
rect 117400 692910 117510 693150
rect 117750 692910 117840 693150
rect 118080 692910 118170 693150
rect 118410 692910 118500 693150
rect 118740 692910 118850 693150
rect 119090 692910 119180 693150
rect 119420 692910 119510 693150
rect 119750 692910 119840 693150
rect 120080 692910 120190 693150
rect 120430 692910 120520 693150
rect 120760 692910 120850 693150
rect 121090 692910 121180 693150
rect 121420 692910 121530 693150
rect 121770 692910 122190 693150
rect 122430 692910 122520 693150
rect 122760 692910 122850 693150
rect 123090 692910 123180 693150
rect 123420 692910 123530 693150
rect 123770 692910 123860 693150
rect 124100 692910 124190 693150
rect 124430 692910 124520 693150
rect 124760 692910 124870 693150
rect 125110 692910 125200 693150
rect 125440 692910 125530 693150
rect 125770 692910 125860 693150
rect 126100 692910 126210 693150
rect 126450 692910 126540 693150
rect 126780 692910 126870 693150
rect 127110 692910 127200 693150
rect 127440 692910 127550 693150
rect 127790 692910 127880 693150
rect 128120 692910 128210 693150
rect 128450 692910 128540 693150
rect 128780 692910 128890 693150
rect 129130 692910 129220 693150
rect 129460 692910 129550 693150
rect 129790 692910 129880 693150
rect 130120 692910 130230 693150
rect 130470 692910 130560 693150
rect 130800 692910 130890 693150
rect 131130 692910 131220 693150
rect 131460 692910 131570 693150
rect 131810 692910 131900 693150
rect 132140 692910 132230 693150
rect 132470 692910 132560 693150
rect 132800 692910 132910 693150
rect 133150 692910 133570 693150
rect 133810 692910 133900 693150
rect 134140 692910 134230 693150
rect 134470 692910 134560 693150
rect 134800 692910 134910 693150
rect 135150 692910 135240 693150
rect 135480 692910 135570 693150
rect 135810 692910 135900 693150
rect 136140 692910 136250 693150
rect 136490 692910 136580 693150
rect 136820 692910 136910 693150
rect 137150 692910 137240 693150
rect 137480 692910 137590 693150
rect 137830 692910 137920 693150
rect 138160 692910 138250 693150
rect 138490 692910 138580 693150
rect 138820 692910 138930 693150
rect 139170 692910 139260 693150
rect 139500 692910 139590 693150
rect 139830 692910 139920 693150
rect 140160 692910 140270 693150
rect 140510 692910 140600 693150
rect 140840 692910 140930 693150
rect 141170 692910 141260 693150
rect 141500 692910 141610 693150
rect 141850 692910 141940 693150
rect 142180 692910 142270 693150
rect 142510 692910 142600 693150
rect 142840 692910 142950 693150
rect 143190 692910 143280 693150
rect 143520 692910 143610 693150
rect 143850 692910 143940 693150
rect 144180 692910 144290 693150
rect 144530 692910 144950 693150
rect 145190 692910 145280 693150
rect 145520 692910 145610 693150
rect 145850 692910 145940 693150
rect 146180 692910 146290 693150
rect 146530 692910 146620 693150
rect 146860 692910 146950 693150
rect 147190 692910 147280 693150
rect 147520 692910 147630 693150
rect 147870 692910 147960 693150
rect 148200 692910 148290 693150
rect 148530 692910 148620 693150
rect 148860 692910 148970 693150
rect 149210 692910 149300 693150
rect 149540 692910 149630 693150
rect 149870 692910 149960 693150
rect 150200 692910 150310 693150
rect 150550 692910 150640 693150
rect 150880 692910 150970 693150
rect 151210 692910 151300 693150
rect 151540 692910 151650 693150
rect 151890 692910 151980 693150
rect 152220 692910 152310 693150
rect 152550 692910 152640 693150
rect 152880 692910 152990 693150
rect 153230 692910 153320 693150
rect 153560 692910 153650 693150
rect 153890 692910 153980 693150
rect 154220 692910 154330 693150
rect 154570 692910 154660 693150
rect 154900 692910 154990 693150
rect 155230 692910 155320 693150
rect 155560 692910 155670 693150
rect 155910 692910 155960 693150
rect 110760 692820 155960 692910
rect 110760 692580 110810 692820
rect 111050 692580 111140 692820
rect 111380 692580 111470 692820
rect 111710 692580 111800 692820
rect 112040 692580 112150 692820
rect 112390 692580 112480 692820
rect 112720 692580 112810 692820
rect 113050 692580 113140 692820
rect 113380 692580 113490 692820
rect 113730 692580 113820 692820
rect 114060 692580 114150 692820
rect 114390 692580 114480 692820
rect 114720 692580 114830 692820
rect 115070 692580 115160 692820
rect 115400 692580 115490 692820
rect 115730 692580 115820 692820
rect 116060 692580 116170 692820
rect 116410 692580 116500 692820
rect 116740 692580 116830 692820
rect 117070 692580 117160 692820
rect 117400 692580 117510 692820
rect 117750 692580 117840 692820
rect 118080 692580 118170 692820
rect 118410 692580 118500 692820
rect 118740 692580 118850 692820
rect 119090 692580 119180 692820
rect 119420 692580 119510 692820
rect 119750 692580 119840 692820
rect 120080 692580 120190 692820
rect 120430 692580 120520 692820
rect 120760 692580 120850 692820
rect 121090 692580 121180 692820
rect 121420 692580 121530 692820
rect 121770 692580 122190 692820
rect 122430 692580 122520 692820
rect 122760 692580 122850 692820
rect 123090 692580 123180 692820
rect 123420 692580 123530 692820
rect 123770 692580 123860 692820
rect 124100 692580 124190 692820
rect 124430 692580 124520 692820
rect 124760 692580 124870 692820
rect 125110 692580 125200 692820
rect 125440 692580 125530 692820
rect 125770 692580 125860 692820
rect 126100 692580 126210 692820
rect 126450 692580 126540 692820
rect 126780 692580 126870 692820
rect 127110 692580 127200 692820
rect 127440 692580 127550 692820
rect 127790 692580 127880 692820
rect 128120 692580 128210 692820
rect 128450 692580 128540 692820
rect 128780 692580 128890 692820
rect 129130 692580 129220 692820
rect 129460 692580 129550 692820
rect 129790 692580 129880 692820
rect 130120 692580 130230 692820
rect 130470 692580 130560 692820
rect 130800 692580 130890 692820
rect 131130 692580 131220 692820
rect 131460 692580 131570 692820
rect 131810 692580 131900 692820
rect 132140 692580 132230 692820
rect 132470 692580 132560 692820
rect 132800 692580 132910 692820
rect 133150 692580 133570 692820
rect 133810 692580 133900 692820
rect 134140 692580 134230 692820
rect 134470 692580 134560 692820
rect 134800 692580 134910 692820
rect 135150 692580 135240 692820
rect 135480 692580 135570 692820
rect 135810 692580 135900 692820
rect 136140 692580 136250 692820
rect 136490 692580 136580 692820
rect 136820 692580 136910 692820
rect 137150 692580 137240 692820
rect 137480 692580 137590 692820
rect 137830 692580 137920 692820
rect 138160 692580 138250 692820
rect 138490 692580 138580 692820
rect 138820 692580 138930 692820
rect 139170 692580 139260 692820
rect 139500 692580 139590 692820
rect 139830 692580 139920 692820
rect 140160 692580 140270 692820
rect 140510 692580 140600 692820
rect 140840 692580 140930 692820
rect 141170 692580 141260 692820
rect 141500 692580 141610 692820
rect 141850 692580 141940 692820
rect 142180 692580 142270 692820
rect 142510 692580 142600 692820
rect 142840 692580 142950 692820
rect 143190 692580 143280 692820
rect 143520 692580 143610 692820
rect 143850 692580 143940 692820
rect 144180 692580 144290 692820
rect 144530 692580 144950 692820
rect 145190 692580 145280 692820
rect 145520 692580 145610 692820
rect 145850 692580 145940 692820
rect 146180 692580 146290 692820
rect 146530 692580 146620 692820
rect 146860 692580 146950 692820
rect 147190 692580 147280 692820
rect 147520 692580 147630 692820
rect 147870 692580 147960 692820
rect 148200 692580 148290 692820
rect 148530 692580 148620 692820
rect 148860 692580 148970 692820
rect 149210 692580 149300 692820
rect 149540 692580 149630 692820
rect 149870 692580 149960 692820
rect 150200 692580 150310 692820
rect 150550 692580 150640 692820
rect 150880 692580 150970 692820
rect 151210 692580 151300 692820
rect 151540 692580 151650 692820
rect 151890 692580 151980 692820
rect 152220 692580 152310 692820
rect 152550 692580 152640 692820
rect 152880 692580 152990 692820
rect 153230 692580 153320 692820
rect 153560 692580 153650 692820
rect 153890 692580 153980 692820
rect 154220 692580 154330 692820
rect 154570 692580 154660 692820
rect 154900 692580 154990 692820
rect 155230 692580 155320 692820
rect 155560 692580 155670 692820
rect 155910 692580 155960 692820
rect 110760 692490 155960 692580
rect 110760 692250 110810 692490
rect 111050 692250 111140 692490
rect 111380 692250 111470 692490
rect 111710 692250 111800 692490
rect 112040 692250 112150 692490
rect 112390 692250 112480 692490
rect 112720 692250 112810 692490
rect 113050 692250 113140 692490
rect 113380 692250 113490 692490
rect 113730 692250 113820 692490
rect 114060 692250 114150 692490
rect 114390 692250 114480 692490
rect 114720 692250 114830 692490
rect 115070 692250 115160 692490
rect 115400 692250 115490 692490
rect 115730 692250 115820 692490
rect 116060 692250 116170 692490
rect 116410 692250 116500 692490
rect 116740 692250 116830 692490
rect 117070 692250 117160 692490
rect 117400 692250 117510 692490
rect 117750 692250 117840 692490
rect 118080 692250 118170 692490
rect 118410 692250 118500 692490
rect 118740 692250 118850 692490
rect 119090 692250 119180 692490
rect 119420 692250 119510 692490
rect 119750 692250 119840 692490
rect 120080 692250 120190 692490
rect 120430 692250 120520 692490
rect 120760 692250 120850 692490
rect 121090 692250 121180 692490
rect 121420 692250 121530 692490
rect 121770 692250 122190 692490
rect 122430 692250 122520 692490
rect 122760 692250 122850 692490
rect 123090 692250 123180 692490
rect 123420 692250 123530 692490
rect 123770 692250 123860 692490
rect 124100 692250 124190 692490
rect 124430 692250 124520 692490
rect 124760 692250 124870 692490
rect 125110 692250 125200 692490
rect 125440 692250 125530 692490
rect 125770 692250 125860 692490
rect 126100 692250 126210 692490
rect 126450 692250 126540 692490
rect 126780 692250 126870 692490
rect 127110 692250 127200 692490
rect 127440 692250 127550 692490
rect 127790 692250 127880 692490
rect 128120 692250 128210 692490
rect 128450 692250 128540 692490
rect 128780 692250 128890 692490
rect 129130 692250 129220 692490
rect 129460 692250 129550 692490
rect 129790 692250 129880 692490
rect 130120 692250 130230 692490
rect 130470 692250 130560 692490
rect 130800 692250 130890 692490
rect 131130 692250 131220 692490
rect 131460 692250 131570 692490
rect 131810 692250 131900 692490
rect 132140 692250 132230 692490
rect 132470 692250 132560 692490
rect 132800 692250 132910 692490
rect 133150 692250 133570 692490
rect 133810 692250 133900 692490
rect 134140 692250 134230 692490
rect 134470 692250 134560 692490
rect 134800 692250 134910 692490
rect 135150 692250 135240 692490
rect 135480 692250 135570 692490
rect 135810 692250 135900 692490
rect 136140 692250 136250 692490
rect 136490 692250 136580 692490
rect 136820 692250 136910 692490
rect 137150 692250 137240 692490
rect 137480 692250 137590 692490
rect 137830 692250 137920 692490
rect 138160 692250 138250 692490
rect 138490 692250 138580 692490
rect 138820 692250 138930 692490
rect 139170 692250 139260 692490
rect 139500 692250 139590 692490
rect 139830 692250 139920 692490
rect 140160 692250 140270 692490
rect 140510 692250 140600 692490
rect 140840 692250 140930 692490
rect 141170 692250 141260 692490
rect 141500 692250 141610 692490
rect 141850 692250 141940 692490
rect 142180 692250 142270 692490
rect 142510 692250 142600 692490
rect 142840 692250 142950 692490
rect 143190 692250 143280 692490
rect 143520 692250 143610 692490
rect 143850 692250 143940 692490
rect 144180 692250 144290 692490
rect 144530 692250 144950 692490
rect 145190 692250 145280 692490
rect 145520 692250 145610 692490
rect 145850 692250 145940 692490
rect 146180 692250 146290 692490
rect 146530 692250 146620 692490
rect 146860 692250 146950 692490
rect 147190 692250 147280 692490
rect 147520 692250 147630 692490
rect 147870 692250 147960 692490
rect 148200 692250 148290 692490
rect 148530 692250 148620 692490
rect 148860 692250 148970 692490
rect 149210 692250 149300 692490
rect 149540 692250 149630 692490
rect 149870 692250 149960 692490
rect 150200 692250 150310 692490
rect 150550 692250 150640 692490
rect 150880 692250 150970 692490
rect 151210 692250 151300 692490
rect 151540 692250 151650 692490
rect 151890 692250 151980 692490
rect 152220 692250 152310 692490
rect 152550 692250 152640 692490
rect 152880 692250 152990 692490
rect 153230 692250 153320 692490
rect 153560 692250 153650 692490
rect 153890 692250 153980 692490
rect 154220 692250 154330 692490
rect 154570 692250 154660 692490
rect 154900 692250 154990 692490
rect 155230 692250 155320 692490
rect 155560 692250 155670 692490
rect 155910 692250 155960 692490
rect 110760 692160 155960 692250
rect 110760 691920 110810 692160
rect 111050 691920 111140 692160
rect 111380 691920 111470 692160
rect 111710 691920 111800 692160
rect 112040 691920 112150 692160
rect 112390 691920 112480 692160
rect 112720 691920 112810 692160
rect 113050 691920 113140 692160
rect 113380 691920 113490 692160
rect 113730 691920 113820 692160
rect 114060 691920 114150 692160
rect 114390 691920 114480 692160
rect 114720 691920 114830 692160
rect 115070 691920 115160 692160
rect 115400 691920 115490 692160
rect 115730 691920 115820 692160
rect 116060 691920 116170 692160
rect 116410 691920 116500 692160
rect 116740 691920 116830 692160
rect 117070 691920 117160 692160
rect 117400 691920 117510 692160
rect 117750 691920 117840 692160
rect 118080 691920 118170 692160
rect 118410 691920 118500 692160
rect 118740 691920 118850 692160
rect 119090 691920 119180 692160
rect 119420 691920 119510 692160
rect 119750 691920 119840 692160
rect 120080 691920 120190 692160
rect 120430 691920 120520 692160
rect 120760 691920 120850 692160
rect 121090 691920 121180 692160
rect 121420 691920 121530 692160
rect 121770 691920 122190 692160
rect 122430 691920 122520 692160
rect 122760 691920 122850 692160
rect 123090 691920 123180 692160
rect 123420 691920 123530 692160
rect 123770 691920 123860 692160
rect 124100 691920 124190 692160
rect 124430 691920 124520 692160
rect 124760 691920 124870 692160
rect 125110 691920 125200 692160
rect 125440 691920 125530 692160
rect 125770 691920 125860 692160
rect 126100 691920 126210 692160
rect 126450 691920 126540 692160
rect 126780 691920 126870 692160
rect 127110 691920 127200 692160
rect 127440 691920 127550 692160
rect 127790 691920 127880 692160
rect 128120 691920 128210 692160
rect 128450 691920 128540 692160
rect 128780 691920 128890 692160
rect 129130 691920 129220 692160
rect 129460 691920 129550 692160
rect 129790 691920 129880 692160
rect 130120 691920 130230 692160
rect 130470 691920 130560 692160
rect 130800 691920 130890 692160
rect 131130 691920 131220 692160
rect 131460 691920 131570 692160
rect 131810 691920 131900 692160
rect 132140 691920 132230 692160
rect 132470 691920 132560 692160
rect 132800 691920 132910 692160
rect 133150 691920 133570 692160
rect 133810 691920 133900 692160
rect 134140 691920 134230 692160
rect 134470 691920 134560 692160
rect 134800 691920 134910 692160
rect 135150 691920 135240 692160
rect 135480 691920 135570 692160
rect 135810 691920 135900 692160
rect 136140 691920 136250 692160
rect 136490 691920 136580 692160
rect 136820 691920 136910 692160
rect 137150 691920 137240 692160
rect 137480 691920 137590 692160
rect 137830 691920 137920 692160
rect 138160 691920 138250 692160
rect 138490 691920 138580 692160
rect 138820 691920 138930 692160
rect 139170 691920 139260 692160
rect 139500 691920 139590 692160
rect 139830 691920 139920 692160
rect 140160 691920 140270 692160
rect 140510 691920 140600 692160
rect 140840 691920 140930 692160
rect 141170 691920 141260 692160
rect 141500 691920 141610 692160
rect 141850 691920 141940 692160
rect 142180 691920 142270 692160
rect 142510 691920 142600 692160
rect 142840 691920 142950 692160
rect 143190 691920 143280 692160
rect 143520 691920 143610 692160
rect 143850 691920 143940 692160
rect 144180 691920 144290 692160
rect 144530 691920 144950 692160
rect 145190 691920 145280 692160
rect 145520 691920 145610 692160
rect 145850 691920 145940 692160
rect 146180 691920 146290 692160
rect 146530 691920 146620 692160
rect 146860 691920 146950 692160
rect 147190 691920 147280 692160
rect 147520 691920 147630 692160
rect 147870 691920 147960 692160
rect 148200 691920 148290 692160
rect 148530 691920 148620 692160
rect 148860 691920 148970 692160
rect 149210 691920 149300 692160
rect 149540 691920 149630 692160
rect 149870 691920 149960 692160
rect 150200 691920 150310 692160
rect 150550 691920 150640 692160
rect 150880 691920 150970 692160
rect 151210 691920 151300 692160
rect 151540 691920 151650 692160
rect 151890 691920 151980 692160
rect 152220 691920 152310 692160
rect 152550 691920 152640 692160
rect 152880 691920 152990 692160
rect 153230 691920 153320 692160
rect 153560 691920 153650 692160
rect 153890 691920 153980 692160
rect 154220 691920 154330 692160
rect 154570 691920 154660 692160
rect 154900 691920 154990 692160
rect 155230 691920 155320 692160
rect 155560 691920 155670 692160
rect 155910 691920 155960 692160
rect 110760 691810 155960 691920
rect 110760 691570 110810 691810
rect 111050 691570 111140 691810
rect 111380 691570 111470 691810
rect 111710 691570 111800 691810
rect 112040 691570 112150 691810
rect 112390 691570 112480 691810
rect 112720 691570 112810 691810
rect 113050 691570 113140 691810
rect 113380 691570 113490 691810
rect 113730 691570 113820 691810
rect 114060 691570 114150 691810
rect 114390 691570 114480 691810
rect 114720 691570 114830 691810
rect 115070 691570 115160 691810
rect 115400 691570 115490 691810
rect 115730 691570 115820 691810
rect 116060 691570 116170 691810
rect 116410 691570 116500 691810
rect 116740 691570 116830 691810
rect 117070 691570 117160 691810
rect 117400 691570 117510 691810
rect 117750 691570 117840 691810
rect 118080 691570 118170 691810
rect 118410 691570 118500 691810
rect 118740 691570 118850 691810
rect 119090 691570 119180 691810
rect 119420 691570 119510 691810
rect 119750 691570 119840 691810
rect 120080 691570 120190 691810
rect 120430 691570 120520 691810
rect 120760 691570 120850 691810
rect 121090 691570 121180 691810
rect 121420 691570 121530 691810
rect 121770 691570 122190 691810
rect 122430 691570 122520 691810
rect 122760 691570 122850 691810
rect 123090 691570 123180 691810
rect 123420 691570 123530 691810
rect 123770 691570 123860 691810
rect 124100 691570 124190 691810
rect 124430 691570 124520 691810
rect 124760 691570 124870 691810
rect 125110 691570 125200 691810
rect 125440 691570 125530 691810
rect 125770 691570 125860 691810
rect 126100 691570 126210 691810
rect 126450 691570 126540 691810
rect 126780 691570 126870 691810
rect 127110 691570 127200 691810
rect 127440 691570 127550 691810
rect 127790 691570 127880 691810
rect 128120 691570 128210 691810
rect 128450 691570 128540 691810
rect 128780 691570 128890 691810
rect 129130 691570 129220 691810
rect 129460 691570 129550 691810
rect 129790 691570 129880 691810
rect 130120 691570 130230 691810
rect 130470 691570 130560 691810
rect 130800 691570 130890 691810
rect 131130 691570 131220 691810
rect 131460 691570 131570 691810
rect 131810 691570 131900 691810
rect 132140 691570 132230 691810
rect 132470 691570 132560 691810
rect 132800 691570 132910 691810
rect 133150 691570 133570 691810
rect 133810 691570 133900 691810
rect 134140 691570 134230 691810
rect 134470 691570 134560 691810
rect 134800 691570 134910 691810
rect 135150 691570 135240 691810
rect 135480 691570 135570 691810
rect 135810 691570 135900 691810
rect 136140 691570 136250 691810
rect 136490 691570 136580 691810
rect 136820 691570 136910 691810
rect 137150 691570 137240 691810
rect 137480 691570 137590 691810
rect 137830 691570 137920 691810
rect 138160 691570 138250 691810
rect 138490 691570 138580 691810
rect 138820 691570 138930 691810
rect 139170 691570 139260 691810
rect 139500 691570 139590 691810
rect 139830 691570 139920 691810
rect 140160 691570 140270 691810
rect 140510 691570 140600 691810
rect 140840 691570 140930 691810
rect 141170 691570 141260 691810
rect 141500 691570 141610 691810
rect 141850 691570 141940 691810
rect 142180 691570 142270 691810
rect 142510 691570 142600 691810
rect 142840 691570 142950 691810
rect 143190 691570 143280 691810
rect 143520 691570 143610 691810
rect 143850 691570 143940 691810
rect 144180 691570 144290 691810
rect 144530 691570 144950 691810
rect 145190 691570 145280 691810
rect 145520 691570 145610 691810
rect 145850 691570 145940 691810
rect 146180 691570 146290 691810
rect 146530 691570 146620 691810
rect 146860 691570 146950 691810
rect 147190 691570 147280 691810
rect 147520 691570 147630 691810
rect 147870 691570 147960 691810
rect 148200 691570 148290 691810
rect 148530 691570 148620 691810
rect 148860 691570 148970 691810
rect 149210 691570 149300 691810
rect 149540 691570 149630 691810
rect 149870 691570 149960 691810
rect 150200 691570 150310 691810
rect 150550 691570 150640 691810
rect 150880 691570 150970 691810
rect 151210 691570 151300 691810
rect 151540 691570 151650 691810
rect 151890 691570 151980 691810
rect 152220 691570 152310 691810
rect 152550 691570 152640 691810
rect 152880 691570 152990 691810
rect 153230 691570 153320 691810
rect 153560 691570 153650 691810
rect 153890 691570 153980 691810
rect 154220 691570 154330 691810
rect 154570 691570 154660 691810
rect 154900 691570 154990 691810
rect 155230 691570 155320 691810
rect 155560 691570 155670 691810
rect 155910 691570 155960 691810
rect 110760 691480 155960 691570
rect 110760 691240 110810 691480
rect 111050 691240 111140 691480
rect 111380 691240 111470 691480
rect 111710 691240 111800 691480
rect 112040 691240 112150 691480
rect 112390 691240 112480 691480
rect 112720 691240 112810 691480
rect 113050 691240 113140 691480
rect 113380 691240 113490 691480
rect 113730 691240 113820 691480
rect 114060 691240 114150 691480
rect 114390 691240 114480 691480
rect 114720 691240 114830 691480
rect 115070 691240 115160 691480
rect 115400 691240 115490 691480
rect 115730 691240 115820 691480
rect 116060 691240 116170 691480
rect 116410 691240 116500 691480
rect 116740 691240 116830 691480
rect 117070 691240 117160 691480
rect 117400 691240 117510 691480
rect 117750 691240 117840 691480
rect 118080 691240 118170 691480
rect 118410 691240 118500 691480
rect 118740 691240 118850 691480
rect 119090 691240 119180 691480
rect 119420 691240 119510 691480
rect 119750 691240 119840 691480
rect 120080 691240 120190 691480
rect 120430 691240 120520 691480
rect 120760 691240 120850 691480
rect 121090 691240 121180 691480
rect 121420 691240 121530 691480
rect 121770 691240 122190 691480
rect 122430 691240 122520 691480
rect 122760 691240 122850 691480
rect 123090 691240 123180 691480
rect 123420 691240 123530 691480
rect 123770 691240 123860 691480
rect 124100 691240 124190 691480
rect 124430 691240 124520 691480
rect 124760 691240 124870 691480
rect 125110 691240 125200 691480
rect 125440 691240 125530 691480
rect 125770 691240 125860 691480
rect 126100 691240 126210 691480
rect 126450 691240 126540 691480
rect 126780 691240 126870 691480
rect 127110 691240 127200 691480
rect 127440 691240 127550 691480
rect 127790 691240 127880 691480
rect 128120 691240 128210 691480
rect 128450 691240 128540 691480
rect 128780 691240 128890 691480
rect 129130 691240 129220 691480
rect 129460 691240 129550 691480
rect 129790 691240 129880 691480
rect 130120 691240 130230 691480
rect 130470 691240 130560 691480
rect 130800 691240 130890 691480
rect 131130 691240 131220 691480
rect 131460 691240 131570 691480
rect 131810 691240 131900 691480
rect 132140 691240 132230 691480
rect 132470 691240 132560 691480
rect 132800 691240 132910 691480
rect 133150 691240 133570 691480
rect 133810 691240 133900 691480
rect 134140 691240 134230 691480
rect 134470 691240 134560 691480
rect 134800 691240 134910 691480
rect 135150 691240 135240 691480
rect 135480 691240 135570 691480
rect 135810 691240 135900 691480
rect 136140 691240 136250 691480
rect 136490 691240 136580 691480
rect 136820 691240 136910 691480
rect 137150 691240 137240 691480
rect 137480 691240 137590 691480
rect 137830 691240 137920 691480
rect 138160 691240 138250 691480
rect 138490 691240 138580 691480
rect 138820 691240 138930 691480
rect 139170 691240 139260 691480
rect 139500 691240 139590 691480
rect 139830 691240 139920 691480
rect 140160 691240 140270 691480
rect 140510 691240 140600 691480
rect 140840 691240 140930 691480
rect 141170 691240 141260 691480
rect 141500 691240 141610 691480
rect 141850 691240 141940 691480
rect 142180 691240 142270 691480
rect 142510 691240 142600 691480
rect 142840 691240 142950 691480
rect 143190 691240 143280 691480
rect 143520 691240 143610 691480
rect 143850 691240 143940 691480
rect 144180 691240 144290 691480
rect 144530 691240 144950 691480
rect 145190 691240 145280 691480
rect 145520 691240 145610 691480
rect 145850 691240 145940 691480
rect 146180 691240 146290 691480
rect 146530 691240 146620 691480
rect 146860 691240 146950 691480
rect 147190 691240 147280 691480
rect 147520 691240 147630 691480
rect 147870 691240 147960 691480
rect 148200 691240 148290 691480
rect 148530 691240 148620 691480
rect 148860 691240 148970 691480
rect 149210 691240 149300 691480
rect 149540 691240 149630 691480
rect 149870 691240 149960 691480
rect 150200 691240 150310 691480
rect 150550 691240 150640 691480
rect 150880 691240 150970 691480
rect 151210 691240 151300 691480
rect 151540 691240 151650 691480
rect 151890 691240 151980 691480
rect 152220 691240 152310 691480
rect 152550 691240 152640 691480
rect 152880 691240 152990 691480
rect 153230 691240 153320 691480
rect 153560 691240 153650 691480
rect 153890 691240 153980 691480
rect 154220 691240 154330 691480
rect 154570 691240 154660 691480
rect 154900 691240 154990 691480
rect 155230 691240 155320 691480
rect 155560 691240 155670 691480
rect 155910 691240 155960 691480
rect 110760 691150 155960 691240
rect 110760 690910 110810 691150
rect 111050 690910 111140 691150
rect 111380 690910 111470 691150
rect 111710 690910 111800 691150
rect 112040 690910 112150 691150
rect 112390 690910 112480 691150
rect 112720 690910 112810 691150
rect 113050 690910 113140 691150
rect 113380 690910 113490 691150
rect 113730 690910 113820 691150
rect 114060 690910 114150 691150
rect 114390 690910 114480 691150
rect 114720 690910 114830 691150
rect 115070 690910 115160 691150
rect 115400 690910 115490 691150
rect 115730 690910 115820 691150
rect 116060 690910 116170 691150
rect 116410 690910 116500 691150
rect 116740 690910 116830 691150
rect 117070 690910 117160 691150
rect 117400 690910 117510 691150
rect 117750 690910 117840 691150
rect 118080 690910 118170 691150
rect 118410 690910 118500 691150
rect 118740 690910 118850 691150
rect 119090 690910 119180 691150
rect 119420 690910 119510 691150
rect 119750 690910 119840 691150
rect 120080 690910 120190 691150
rect 120430 690910 120520 691150
rect 120760 690910 120850 691150
rect 121090 690910 121180 691150
rect 121420 690910 121530 691150
rect 121770 690910 122190 691150
rect 122430 690910 122520 691150
rect 122760 690910 122850 691150
rect 123090 690910 123180 691150
rect 123420 690910 123530 691150
rect 123770 690910 123860 691150
rect 124100 690910 124190 691150
rect 124430 690910 124520 691150
rect 124760 690910 124870 691150
rect 125110 690910 125200 691150
rect 125440 690910 125530 691150
rect 125770 690910 125860 691150
rect 126100 690910 126210 691150
rect 126450 690910 126540 691150
rect 126780 690910 126870 691150
rect 127110 690910 127200 691150
rect 127440 690910 127550 691150
rect 127790 690910 127880 691150
rect 128120 690910 128210 691150
rect 128450 690910 128540 691150
rect 128780 690910 128890 691150
rect 129130 690910 129220 691150
rect 129460 690910 129550 691150
rect 129790 690910 129880 691150
rect 130120 690910 130230 691150
rect 130470 690910 130560 691150
rect 130800 690910 130890 691150
rect 131130 690910 131220 691150
rect 131460 690910 131570 691150
rect 131810 690910 131900 691150
rect 132140 690910 132230 691150
rect 132470 690910 132560 691150
rect 132800 690910 132910 691150
rect 133150 690910 133570 691150
rect 133810 690910 133900 691150
rect 134140 690910 134230 691150
rect 134470 690910 134560 691150
rect 134800 690910 134910 691150
rect 135150 690910 135240 691150
rect 135480 690910 135570 691150
rect 135810 690910 135900 691150
rect 136140 690910 136250 691150
rect 136490 690910 136580 691150
rect 136820 690910 136910 691150
rect 137150 690910 137240 691150
rect 137480 690910 137590 691150
rect 137830 690910 137920 691150
rect 138160 690910 138250 691150
rect 138490 690910 138580 691150
rect 138820 690910 138930 691150
rect 139170 690910 139260 691150
rect 139500 690910 139590 691150
rect 139830 690910 139920 691150
rect 140160 690910 140270 691150
rect 140510 690910 140600 691150
rect 140840 690910 140930 691150
rect 141170 690910 141260 691150
rect 141500 690910 141610 691150
rect 141850 690910 141940 691150
rect 142180 690910 142270 691150
rect 142510 690910 142600 691150
rect 142840 690910 142950 691150
rect 143190 690910 143280 691150
rect 143520 690910 143610 691150
rect 143850 690910 143940 691150
rect 144180 690910 144290 691150
rect 144530 690910 144950 691150
rect 145190 690910 145280 691150
rect 145520 690910 145610 691150
rect 145850 690910 145940 691150
rect 146180 690910 146290 691150
rect 146530 690910 146620 691150
rect 146860 690910 146950 691150
rect 147190 690910 147280 691150
rect 147520 690910 147630 691150
rect 147870 690910 147960 691150
rect 148200 690910 148290 691150
rect 148530 690910 148620 691150
rect 148860 690910 148970 691150
rect 149210 690910 149300 691150
rect 149540 690910 149630 691150
rect 149870 690910 149960 691150
rect 150200 690910 150310 691150
rect 150550 690910 150640 691150
rect 150880 690910 150970 691150
rect 151210 690910 151300 691150
rect 151540 690910 151650 691150
rect 151890 690910 151980 691150
rect 152220 690910 152310 691150
rect 152550 690910 152640 691150
rect 152880 690910 152990 691150
rect 153230 690910 153320 691150
rect 153560 690910 153650 691150
rect 153890 690910 153980 691150
rect 154220 690910 154330 691150
rect 154570 690910 154660 691150
rect 154900 690910 154990 691150
rect 155230 690910 155320 691150
rect 155560 690910 155670 691150
rect 155910 690910 155960 691150
rect 110760 690820 155960 690910
rect 110760 690580 110810 690820
rect 111050 690580 111140 690820
rect 111380 690580 111470 690820
rect 111710 690580 111800 690820
rect 112040 690580 112150 690820
rect 112390 690580 112480 690820
rect 112720 690580 112810 690820
rect 113050 690580 113140 690820
rect 113380 690580 113490 690820
rect 113730 690580 113820 690820
rect 114060 690580 114150 690820
rect 114390 690580 114480 690820
rect 114720 690580 114830 690820
rect 115070 690580 115160 690820
rect 115400 690580 115490 690820
rect 115730 690580 115820 690820
rect 116060 690580 116170 690820
rect 116410 690580 116500 690820
rect 116740 690580 116830 690820
rect 117070 690580 117160 690820
rect 117400 690580 117510 690820
rect 117750 690580 117840 690820
rect 118080 690580 118170 690820
rect 118410 690580 118500 690820
rect 118740 690580 118850 690820
rect 119090 690580 119180 690820
rect 119420 690580 119510 690820
rect 119750 690580 119840 690820
rect 120080 690580 120190 690820
rect 120430 690580 120520 690820
rect 120760 690580 120850 690820
rect 121090 690580 121180 690820
rect 121420 690580 121530 690820
rect 121770 690580 122190 690820
rect 122430 690580 122520 690820
rect 122760 690580 122850 690820
rect 123090 690580 123180 690820
rect 123420 690580 123530 690820
rect 123770 690580 123860 690820
rect 124100 690580 124190 690820
rect 124430 690580 124520 690820
rect 124760 690580 124870 690820
rect 125110 690580 125200 690820
rect 125440 690580 125530 690820
rect 125770 690580 125860 690820
rect 126100 690580 126210 690820
rect 126450 690580 126540 690820
rect 126780 690580 126870 690820
rect 127110 690580 127200 690820
rect 127440 690580 127550 690820
rect 127790 690580 127880 690820
rect 128120 690580 128210 690820
rect 128450 690580 128540 690820
rect 128780 690580 128890 690820
rect 129130 690580 129220 690820
rect 129460 690580 129550 690820
rect 129790 690580 129880 690820
rect 130120 690580 130230 690820
rect 130470 690580 130560 690820
rect 130800 690580 130890 690820
rect 131130 690580 131220 690820
rect 131460 690580 131570 690820
rect 131810 690580 131900 690820
rect 132140 690580 132230 690820
rect 132470 690580 132560 690820
rect 132800 690580 132910 690820
rect 133150 690580 133570 690820
rect 133810 690580 133900 690820
rect 134140 690580 134230 690820
rect 134470 690580 134560 690820
rect 134800 690580 134910 690820
rect 135150 690580 135240 690820
rect 135480 690580 135570 690820
rect 135810 690580 135900 690820
rect 136140 690580 136250 690820
rect 136490 690580 136580 690820
rect 136820 690580 136910 690820
rect 137150 690580 137240 690820
rect 137480 690580 137590 690820
rect 137830 690580 137920 690820
rect 138160 690580 138250 690820
rect 138490 690580 138580 690820
rect 138820 690580 138930 690820
rect 139170 690580 139260 690820
rect 139500 690580 139590 690820
rect 139830 690580 139920 690820
rect 140160 690580 140270 690820
rect 140510 690580 140600 690820
rect 140840 690580 140930 690820
rect 141170 690580 141260 690820
rect 141500 690580 141610 690820
rect 141850 690580 141940 690820
rect 142180 690580 142270 690820
rect 142510 690580 142600 690820
rect 142840 690580 142950 690820
rect 143190 690580 143280 690820
rect 143520 690580 143610 690820
rect 143850 690580 143940 690820
rect 144180 690580 144290 690820
rect 144530 690580 144950 690820
rect 145190 690580 145280 690820
rect 145520 690580 145610 690820
rect 145850 690580 145940 690820
rect 146180 690580 146290 690820
rect 146530 690580 146620 690820
rect 146860 690580 146950 690820
rect 147190 690580 147280 690820
rect 147520 690580 147630 690820
rect 147870 690580 147960 690820
rect 148200 690580 148290 690820
rect 148530 690580 148620 690820
rect 148860 690580 148970 690820
rect 149210 690580 149300 690820
rect 149540 690580 149630 690820
rect 149870 690580 149960 690820
rect 150200 690580 150310 690820
rect 150550 690580 150640 690820
rect 150880 690580 150970 690820
rect 151210 690580 151300 690820
rect 151540 690580 151650 690820
rect 151890 690580 151980 690820
rect 152220 690580 152310 690820
rect 152550 690580 152640 690820
rect 152880 690580 152990 690820
rect 153230 690580 153320 690820
rect 153560 690580 153650 690820
rect 153890 690580 153980 690820
rect 154220 690580 154330 690820
rect 154570 690580 154660 690820
rect 154900 690580 154990 690820
rect 155230 690580 155320 690820
rect 155560 690580 155670 690820
rect 155910 690580 155960 690820
rect 110760 690470 155960 690580
rect 110760 690230 110810 690470
rect 111050 690230 111140 690470
rect 111380 690230 111470 690470
rect 111710 690230 111800 690470
rect 112040 690230 112150 690470
rect 112390 690230 112480 690470
rect 112720 690230 112810 690470
rect 113050 690230 113140 690470
rect 113380 690230 113490 690470
rect 113730 690230 113820 690470
rect 114060 690230 114150 690470
rect 114390 690230 114480 690470
rect 114720 690230 114830 690470
rect 115070 690230 115160 690470
rect 115400 690230 115490 690470
rect 115730 690230 115820 690470
rect 116060 690230 116170 690470
rect 116410 690230 116500 690470
rect 116740 690230 116830 690470
rect 117070 690230 117160 690470
rect 117400 690230 117510 690470
rect 117750 690230 117840 690470
rect 118080 690230 118170 690470
rect 118410 690230 118500 690470
rect 118740 690230 118850 690470
rect 119090 690230 119180 690470
rect 119420 690230 119510 690470
rect 119750 690230 119840 690470
rect 120080 690230 120190 690470
rect 120430 690230 120520 690470
rect 120760 690230 120850 690470
rect 121090 690230 121180 690470
rect 121420 690230 121530 690470
rect 121770 690230 122190 690470
rect 122430 690230 122520 690470
rect 122760 690230 122850 690470
rect 123090 690230 123180 690470
rect 123420 690230 123530 690470
rect 123770 690230 123860 690470
rect 124100 690230 124190 690470
rect 124430 690230 124520 690470
rect 124760 690230 124870 690470
rect 125110 690230 125200 690470
rect 125440 690230 125530 690470
rect 125770 690230 125860 690470
rect 126100 690230 126210 690470
rect 126450 690230 126540 690470
rect 126780 690230 126870 690470
rect 127110 690230 127200 690470
rect 127440 690230 127550 690470
rect 127790 690230 127880 690470
rect 128120 690230 128210 690470
rect 128450 690230 128540 690470
rect 128780 690230 128890 690470
rect 129130 690230 129220 690470
rect 129460 690230 129550 690470
rect 129790 690230 129880 690470
rect 130120 690230 130230 690470
rect 130470 690230 130560 690470
rect 130800 690230 130890 690470
rect 131130 690230 131220 690470
rect 131460 690230 131570 690470
rect 131810 690230 131900 690470
rect 132140 690230 132230 690470
rect 132470 690230 132560 690470
rect 132800 690230 132910 690470
rect 133150 690230 133570 690470
rect 133810 690230 133900 690470
rect 134140 690230 134230 690470
rect 134470 690230 134560 690470
rect 134800 690230 134910 690470
rect 135150 690230 135240 690470
rect 135480 690230 135570 690470
rect 135810 690230 135900 690470
rect 136140 690230 136250 690470
rect 136490 690230 136580 690470
rect 136820 690230 136910 690470
rect 137150 690230 137240 690470
rect 137480 690230 137590 690470
rect 137830 690230 137920 690470
rect 138160 690230 138250 690470
rect 138490 690230 138580 690470
rect 138820 690230 138930 690470
rect 139170 690230 139260 690470
rect 139500 690230 139590 690470
rect 139830 690230 139920 690470
rect 140160 690230 140270 690470
rect 140510 690230 140600 690470
rect 140840 690230 140930 690470
rect 141170 690230 141260 690470
rect 141500 690230 141610 690470
rect 141850 690230 141940 690470
rect 142180 690230 142270 690470
rect 142510 690230 142600 690470
rect 142840 690230 142950 690470
rect 143190 690230 143280 690470
rect 143520 690230 143610 690470
rect 143850 690230 143940 690470
rect 144180 690230 144290 690470
rect 144530 690230 144950 690470
rect 145190 690230 145280 690470
rect 145520 690230 145610 690470
rect 145850 690230 145940 690470
rect 146180 690230 146290 690470
rect 146530 690230 146620 690470
rect 146860 690230 146950 690470
rect 147190 690230 147280 690470
rect 147520 690230 147630 690470
rect 147870 690230 147960 690470
rect 148200 690230 148290 690470
rect 148530 690230 148620 690470
rect 148860 690230 148970 690470
rect 149210 690230 149300 690470
rect 149540 690230 149630 690470
rect 149870 690230 149960 690470
rect 150200 690230 150310 690470
rect 150550 690230 150640 690470
rect 150880 690230 150970 690470
rect 151210 690230 151300 690470
rect 151540 690230 151650 690470
rect 151890 690230 151980 690470
rect 152220 690230 152310 690470
rect 152550 690230 152640 690470
rect 152880 690230 152990 690470
rect 153230 690230 153320 690470
rect 153560 690230 153650 690470
rect 153890 690230 153980 690470
rect 154220 690230 154330 690470
rect 154570 690230 154660 690470
rect 154900 690230 154990 690470
rect 155230 690230 155320 690470
rect 155560 690230 155670 690470
rect 155910 690230 155960 690470
rect 110760 690140 155960 690230
rect 110760 689900 110810 690140
rect 111050 689900 111140 690140
rect 111380 689900 111470 690140
rect 111710 689900 111800 690140
rect 112040 689900 112150 690140
rect 112390 689900 112480 690140
rect 112720 689900 112810 690140
rect 113050 689900 113140 690140
rect 113380 689900 113490 690140
rect 113730 689900 113820 690140
rect 114060 689900 114150 690140
rect 114390 689900 114480 690140
rect 114720 689900 114830 690140
rect 115070 689900 115160 690140
rect 115400 689900 115490 690140
rect 115730 689900 115820 690140
rect 116060 689900 116170 690140
rect 116410 689900 116500 690140
rect 116740 689900 116830 690140
rect 117070 689900 117160 690140
rect 117400 689900 117510 690140
rect 117750 689900 117840 690140
rect 118080 689900 118170 690140
rect 118410 689900 118500 690140
rect 118740 689900 118850 690140
rect 119090 689900 119180 690140
rect 119420 689900 119510 690140
rect 119750 689900 119840 690140
rect 120080 689900 120190 690140
rect 120430 689900 120520 690140
rect 120760 689900 120850 690140
rect 121090 689900 121180 690140
rect 121420 689900 121530 690140
rect 121770 689900 122190 690140
rect 122430 689900 122520 690140
rect 122760 689900 122850 690140
rect 123090 689900 123180 690140
rect 123420 689900 123530 690140
rect 123770 689900 123860 690140
rect 124100 689900 124190 690140
rect 124430 689900 124520 690140
rect 124760 689900 124870 690140
rect 125110 689900 125200 690140
rect 125440 689900 125530 690140
rect 125770 689900 125860 690140
rect 126100 689900 126210 690140
rect 126450 689900 126540 690140
rect 126780 689900 126870 690140
rect 127110 689900 127200 690140
rect 127440 689900 127550 690140
rect 127790 689900 127880 690140
rect 128120 689900 128210 690140
rect 128450 689900 128540 690140
rect 128780 689900 128890 690140
rect 129130 689900 129220 690140
rect 129460 689900 129550 690140
rect 129790 689900 129880 690140
rect 130120 689900 130230 690140
rect 130470 689900 130560 690140
rect 130800 689900 130890 690140
rect 131130 689900 131220 690140
rect 131460 689900 131570 690140
rect 131810 689900 131900 690140
rect 132140 689900 132230 690140
rect 132470 689900 132560 690140
rect 132800 689900 132910 690140
rect 133150 689900 133570 690140
rect 133810 689900 133900 690140
rect 134140 689900 134230 690140
rect 134470 689900 134560 690140
rect 134800 689900 134910 690140
rect 135150 689900 135240 690140
rect 135480 689900 135570 690140
rect 135810 689900 135900 690140
rect 136140 689900 136250 690140
rect 136490 689900 136580 690140
rect 136820 689900 136910 690140
rect 137150 689900 137240 690140
rect 137480 689900 137590 690140
rect 137830 689900 137920 690140
rect 138160 689900 138250 690140
rect 138490 689900 138580 690140
rect 138820 689900 138930 690140
rect 139170 689900 139260 690140
rect 139500 689900 139590 690140
rect 139830 689900 139920 690140
rect 140160 689900 140270 690140
rect 140510 689900 140600 690140
rect 140840 689900 140930 690140
rect 141170 689900 141260 690140
rect 141500 689900 141610 690140
rect 141850 689900 141940 690140
rect 142180 689900 142270 690140
rect 142510 689900 142600 690140
rect 142840 689900 142950 690140
rect 143190 689900 143280 690140
rect 143520 689900 143610 690140
rect 143850 689900 143940 690140
rect 144180 689900 144290 690140
rect 144530 689900 144950 690140
rect 145190 689900 145280 690140
rect 145520 689900 145610 690140
rect 145850 689900 145940 690140
rect 146180 689900 146290 690140
rect 146530 689900 146620 690140
rect 146860 689900 146950 690140
rect 147190 689900 147280 690140
rect 147520 689900 147630 690140
rect 147870 689900 147960 690140
rect 148200 689900 148290 690140
rect 148530 689900 148620 690140
rect 148860 689900 148970 690140
rect 149210 689900 149300 690140
rect 149540 689900 149630 690140
rect 149870 689900 149960 690140
rect 150200 689900 150310 690140
rect 150550 689900 150640 690140
rect 150880 689900 150970 690140
rect 151210 689900 151300 690140
rect 151540 689900 151650 690140
rect 151890 689900 151980 690140
rect 152220 689900 152310 690140
rect 152550 689900 152640 690140
rect 152880 689900 152990 690140
rect 153230 689900 153320 690140
rect 153560 689900 153650 690140
rect 153890 689900 153980 690140
rect 154220 689900 154330 690140
rect 154570 689900 154660 690140
rect 154900 689900 154990 690140
rect 155230 689900 155320 690140
rect 155560 689900 155670 690140
rect 155910 689900 155960 690140
rect 175894 693000 180894 704800
rect 217294 693000 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 175894 690100 186694 693000
rect 211494 690100 222294 693000
rect 110760 689810 155960 689900
rect 110760 689570 110810 689810
rect 111050 689570 111140 689810
rect 111380 689570 111470 689810
rect 111710 689570 111800 689810
rect 112040 689570 112150 689810
rect 112390 689570 112480 689810
rect 112720 689570 112810 689810
rect 113050 689570 113140 689810
rect 113380 689570 113490 689810
rect 113730 689570 113820 689810
rect 114060 689570 114150 689810
rect 114390 689570 114480 689810
rect 114720 689570 114830 689810
rect 115070 689570 115160 689810
rect 115400 689570 115490 689810
rect 115730 689570 115820 689810
rect 116060 689570 116170 689810
rect 116410 689570 116500 689810
rect 116740 689570 116830 689810
rect 117070 689570 117160 689810
rect 117400 689570 117510 689810
rect 117750 689570 117840 689810
rect 118080 689570 118170 689810
rect 118410 689570 118500 689810
rect 118740 689570 118850 689810
rect 119090 689570 119180 689810
rect 119420 689570 119510 689810
rect 119750 689570 119840 689810
rect 120080 689570 120190 689810
rect 120430 689570 120520 689810
rect 120760 689570 120850 689810
rect 121090 689570 121180 689810
rect 121420 689570 121530 689810
rect 121770 689570 122190 689810
rect 122430 689570 122520 689810
rect 122760 689570 122850 689810
rect 123090 689570 123180 689810
rect 123420 689570 123530 689810
rect 123770 689570 123860 689810
rect 124100 689570 124190 689810
rect 124430 689570 124520 689810
rect 124760 689570 124870 689810
rect 125110 689570 125200 689810
rect 125440 689570 125530 689810
rect 125770 689570 125860 689810
rect 126100 689570 126210 689810
rect 126450 689570 126540 689810
rect 126780 689570 126870 689810
rect 127110 689570 127200 689810
rect 127440 689570 127550 689810
rect 127790 689570 127880 689810
rect 128120 689570 128210 689810
rect 128450 689570 128540 689810
rect 128780 689570 128890 689810
rect 129130 689570 129220 689810
rect 129460 689570 129550 689810
rect 129790 689570 129880 689810
rect 130120 689570 130230 689810
rect 130470 689570 130560 689810
rect 130800 689570 130890 689810
rect 131130 689570 131220 689810
rect 131460 689570 131570 689810
rect 131810 689570 131900 689810
rect 132140 689570 132230 689810
rect 132470 689570 132560 689810
rect 132800 689570 132910 689810
rect 133150 689570 133570 689810
rect 133810 689570 133900 689810
rect 134140 689570 134230 689810
rect 134470 689570 134560 689810
rect 134800 689570 134910 689810
rect 135150 689570 135240 689810
rect 135480 689570 135570 689810
rect 135810 689570 135900 689810
rect 136140 689570 136250 689810
rect 136490 689570 136580 689810
rect 136820 689570 136910 689810
rect 137150 689570 137240 689810
rect 137480 689570 137590 689810
rect 137830 689570 137920 689810
rect 138160 689570 138250 689810
rect 138490 689570 138580 689810
rect 138820 689570 138930 689810
rect 139170 689570 139260 689810
rect 139500 689570 139590 689810
rect 139830 689570 139920 689810
rect 140160 689570 140270 689810
rect 140510 689570 140600 689810
rect 140840 689570 140930 689810
rect 141170 689570 141260 689810
rect 141500 689570 141610 689810
rect 141850 689570 141940 689810
rect 142180 689570 142270 689810
rect 142510 689570 142600 689810
rect 142840 689570 142950 689810
rect 143190 689570 143280 689810
rect 143520 689570 143610 689810
rect 143850 689570 143940 689810
rect 144180 689570 144290 689810
rect 144530 689570 144950 689810
rect 145190 689570 145280 689810
rect 145520 689570 145610 689810
rect 145850 689570 145940 689810
rect 146180 689570 146290 689810
rect 146530 689570 146620 689810
rect 146860 689570 146950 689810
rect 147190 689570 147280 689810
rect 147520 689570 147630 689810
rect 147870 689570 147960 689810
rect 148200 689570 148290 689810
rect 148530 689570 148620 689810
rect 148860 689570 148970 689810
rect 149210 689570 149300 689810
rect 149540 689570 149630 689810
rect 149870 689570 149960 689810
rect 150200 689570 150310 689810
rect 150550 689570 150640 689810
rect 150880 689570 150970 689810
rect 151210 689570 151300 689810
rect 151540 689570 151650 689810
rect 151890 689570 151980 689810
rect 152220 689570 152310 689810
rect 152550 689570 152640 689810
rect 152880 689570 152990 689810
rect 153230 689570 153320 689810
rect 153560 689570 153650 689810
rect 153890 689570 153980 689810
rect 154220 689570 154330 689810
rect 154570 689570 154660 689810
rect 154900 689570 154990 689810
rect 155230 689570 155320 689810
rect 155560 689570 155670 689810
rect 155910 689570 155960 689810
rect 110760 689480 155960 689570
rect 110760 689240 110810 689480
rect 111050 689240 111140 689480
rect 111380 689240 111470 689480
rect 111710 689240 111800 689480
rect 112040 689240 112150 689480
rect 112390 689240 112480 689480
rect 112720 689240 112810 689480
rect 113050 689240 113140 689480
rect 113380 689240 113490 689480
rect 113730 689240 113820 689480
rect 114060 689240 114150 689480
rect 114390 689240 114480 689480
rect 114720 689240 114830 689480
rect 115070 689240 115160 689480
rect 115400 689240 115490 689480
rect 115730 689240 115820 689480
rect 116060 689240 116170 689480
rect 116410 689240 116500 689480
rect 116740 689240 116830 689480
rect 117070 689240 117160 689480
rect 117400 689240 117510 689480
rect 117750 689240 117840 689480
rect 118080 689240 118170 689480
rect 118410 689240 118500 689480
rect 118740 689240 118850 689480
rect 119090 689240 119180 689480
rect 119420 689240 119510 689480
rect 119750 689240 119840 689480
rect 120080 689240 120190 689480
rect 120430 689240 120520 689480
rect 120760 689240 120850 689480
rect 121090 689240 121180 689480
rect 121420 689240 121530 689480
rect 121770 689240 122190 689480
rect 122430 689240 122520 689480
rect 122760 689240 122850 689480
rect 123090 689240 123180 689480
rect 123420 689240 123530 689480
rect 123770 689240 123860 689480
rect 124100 689240 124190 689480
rect 124430 689240 124520 689480
rect 124760 689240 124870 689480
rect 125110 689240 125200 689480
rect 125440 689240 125530 689480
rect 125770 689240 125860 689480
rect 126100 689240 126210 689480
rect 126450 689240 126540 689480
rect 126780 689240 126870 689480
rect 127110 689240 127200 689480
rect 127440 689240 127550 689480
rect 127790 689240 127880 689480
rect 128120 689240 128210 689480
rect 128450 689240 128540 689480
rect 128780 689240 128890 689480
rect 129130 689240 129220 689480
rect 129460 689240 129550 689480
rect 129790 689240 129880 689480
rect 130120 689240 130230 689480
rect 130470 689240 130560 689480
rect 130800 689240 130890 689480
rect 131130 689240 131220 689480
rect 131460 689240 131570 689480
rect 131810 689240 131900 689480
rect 132140 689240 132230 689480
rect 132470 689240 132560 689480
rect 132800 689240 132910 689480
rect 133150 689240 133570 689480
rect 133810 689240 133900 689480
rect 134140 689240 134230 689480
rect 134470 689240 134560 689480
rect 134800 689240 134910 689480
rect 135150 689240 135240 689480
rect 135480 689240 135570 689480
rect 135810 689240 135900 689480
rect 136140 689240 136250 689480
rect 136490 689240 136580 689480
rect 136820 689240 136910 689480
rect 137150 689240 137240 689480
rect 137480 689240 137590 689480
rect 137830 689240 137920 689480
rect 138160 689240 138250 689480
rect 138490 689240 138580 689480
rect 138820 689240 138930 689480
rect 139170 689240 139260 689480
rect 139500 689240 139590 689480
rect 139830 689240 139920 689480
rect 140160 689240 140270 689480
rect 140510 689240 140600 689480
rect 140840 689240 140930 689480
rect 141170 689240 141260 689480
rect 141500 689240 141610 689480
rect 141850 689240 141940 689480
rect 142180 689240 142270 689480
rect 142510 689240 142600 689480
rect 142840 689240 142950 689480
rect 143190 689240 143280 689480
rect 143520 689240 143610 689480
rect 143850 689240 143940 689480
rect 144180 689240 144290 689480
rect 144530 689240 144950 689480
rect 145190 689240 145280 689480
rect 145520 689240 145610 689480
rect 145850 689240 145940 689480
rect 146180 689240 146290 689480
rect 146530 689240 146620 689480
rect 146860 689240 146950 689480
rect 147190 689240 147280 689480
rect 147520 689240 147630 689480
rect 147870 689240 147960 689480
rect 148200 689240 148290 689480
rect 148530 689240 148620 689480
rect 148860 689240 148970 689480
rect 149210 689240 149300 689480
rect 149540 689240 149630 689480
rect 149870 689240 149960 689480
rect 150200 689240 150310 689480
rect 150550 689240 150640 689480
rect 150880 689240 150970 689480
rect 151210 689240 151300 689480
rect 151540 689240 151650 689480
rect 151890 689240 151980 689480
rect 152220 689240 152310 689480
rect 152550 689240 152640 689480
rect 152880 689240 152990 689480
rect 153230 689240 153320 689480
rect 153560 689240 153650 689480
rect 153890 689240 153980 689480
rect 154220 689240 154330 689480
rect 154570 689240 154660 689480
rect 154900 689240 154990 689480
rect 155230 689240 155320 689480
rect 155560 689240 155670 689480
rect 155910 689240 155960 689480
rect 110760 689130 155960 689240
rect 110760 688890 110810 689130
rect 111050 688890 111140 689130
rect 111380 688890 111470 689130
rect 111710 688890 111800 689130
rect 112040 688890 112150 689130
rect 112390 688890 112480 689130
rect 112720 688890 112810 689130
rect 113050 688890 113140 689130
rect 113380 688890 113490 689130
rect 113730 688890 113820 689130
rect 114060 688890 114150 689130
rect 114390 688890 114480 689130
rect 114720 688890 114830 689130
rect 115070 688890 115160 689130
rect 115400 688890 115490 689130
rect 115730 688890 115820 689130
rect 116060 688890 116170 689130
rect 116410 688890 116500 689130
rect 116740 688890 116830 689130
rect 117070 688890 117160 689130
rect 117400 688890 117510 689130
rect 117750 688890 117840 689130
rect 118080 688890 118170 689130
rect 118410 688890 118500 689130
rect 118740 688890 118850 689130
rect 119090 688890 119180 689130
rect 119420 688890 119510 689130
rect 119750 688890 119840 689130
rect 120080 688890 120190 689130
rect 120430 688890 120520 689130
rect 120760 688890 120850 689130
rect 121090 688890 121180 689130
rect 121420 688890 121530 689130
rect 121770 688890 122190 689130
rect 122430 688890 122520 689130
rect 122760 688890 122850 689130
rect 123090 688890 123180 689130
rect 123420 688890 123530 689130
rect 123770 688890 123860 689130
rect 124100 688890 124190 689130
rect 124430 688890 124520 689130
rect 124760 688890 124870 689130
rect 125110 688890 125200 689130
rect 125440 688890 125530 689130
rect 125770 688890 125860 689130
rect 126100 688890 126210 689130
rect 126450 688890 126540 689130
rect 126780 688890 126870 689130
rect 127110 688890 127200 689130
rect 127440 688890 127550 689130
rect 127790 688890 127880 689130
rect 128120 688890 128210 689130
rect 128450 688890 128540 689130
rect 128780 688890 128890 689130
rect 129130 688890 129220 689130
rect 129460 688890 129550 689130
rect 129790 688890 129880 689130
rect 130120 688890 130230 689130
rect 130470 688890 130560 689130
rect 130800 688890 130890 689130
rect 131130 688890 131220 689130
rect 131460 688890 131570 689130
rect 131810 688890 131900 689130
rect 132140 688890 132230 689130
rect 132470 688890 132560 689130
rect 132800 688890 132910 689130
rect 133150 688890 133570 689130
rect 133810 688890 133900 689130
rect 134140 688890 134230 689130
rect 134470 688890 134560 689130
rect 134800 688890 134910 689130
rect 135150 688890 135240 689130
rect 135480 688890 135570 689130
rect 135810 688890 135900 689130
rect 136140 688890 136250 689130
rect 136490 688890 136580 689130
rect 136820 688890 136910 689130
rect 137150 688890 137240 689130
rect 137480 688890 137590 689130
rect 137830 688890 137920 689130
rect 138160 688890 138250 689130
rect 138490 688890 138580 689130
rect 138820 688890 138930 689130
rect 139170 688890 139260 689130
rect 139500 688890 139590 689130
rect 139830 688890 139920 689130
rect 140160 688890 140270 689130
rect 140510 688890 140600 689130
rect 140840 688890 140930 689130
rect 141170 688890 141260 689130
rect 141500 688890 141610 689130
rect 141850 688890 141940 689130
rect 142180 688890 142270 689130
rect 142510 688890 142600 689130
rect 142840 688890 142950 689130
rect 143190 688890 143280 689130
rect 143520 688890 143610 689130
rect 143850 688890 143940 689130
rect 144180 688890 144290 689130
rect 144530 688890 144950 689130
rect 145190 688890 145280 689130
rect 145520 688890 145610 689130
rect 145850 688890 145940 689130
rect 146180 688890 146290 689130
rect 146530 688890 146620 689130
rect 146860 688890 146950 689130
rect 147190 688890 147280 689130
rect 147520 688890 147630 689130
rect 147870 688890 147960 689130
rect 148200 688890 148290 689130
rect 148530 688890 148620 689130
rect 148860 688890 148970 689130
rect 149210 688890 149300 689130
rect 149540 688890 149630 689130
rect 149870 688890 149960 689130
rect 150200 688890 150310 689130
rect 150550 688890 150640 689130
rect 150880 688890 150970 689130
rect 151210 688890 151300 689130
rect 151540 688890 151650 689130
rect 151890 688890 151980 689130
rect 152220 688890 152310 689130
rect 152550 688890 152640 689130
rect 152880 688890 152990 689130
rect 153230 688890 153320 689130
rect 153560 688890 153650 689130
rect 153890 688890 153980 689130
rect 154220 688890 154330 689130
rect 154570 688890 154660 689130
rect 154900 688890 154990 689130
rect 155230 688890 155320 689130
rect 155560 688890 155670 689130
rect 155910 688890 155960 689130
rect 110760 688800 155960 688890
rect 110760 688560 110810 688800
rect 111050 688560 111140 688800
rect 111380 688560 111470 688800
rect 111710 688560 111800 688800
rect 112040 688560 112150 688800
rect 112390 688560 112480 688800
rect 112720 688560 112810 688800
rect 113050 688560 113140 688800
rect 113380 688560 113490 688800
rect 113730 688560 113820 688800
rect 114060 688560 114150 688800
rect 114390 688560 114480 688800
rect 114720 688560 114830 688800
rect 115070 688560 115160 688800
rect 115400 688560 115490 688800
rect 115730 688560 115820 688800
rect 116060 688560 116170 688800
rect 116410 688560 116500 688800
rect 116740 688560 116830 688800
rect 117070 688560 117160 688800
rect 117400 688560 117510 688800
rect 117750 688560 117840 688800
rect 118080 688560 118170 688800
rect 118410 688560 118500 688800
rect 118740 688560 118850 688800
rect 119090 688560 119180 688800
rect 119420 688560 119510 688800
rect 119750 688560 119840 688800
rect 120080 688560 120190 688800
rect 120430 688560 120520 688800
rect 120760 688560 120850 688800
rect 121090 688560 121180 688800
rect 121420 688560 121530 688800
rect 121770 688560 122190 688800
rect 122430 688560 122520 688800
rect 122760 688560 122850 688800
rect 123090 688560 123180 688800
rect 123420 688560 123530 688800
rect 123770 688560 123860 688800
rect 124100 688560 124190 688800
rect 124430 688560 124520 688800
rect 124760 688560 124870 688800
rect 125110 688560 125200 688800
rect 125440 688560 125530 688800
rect 125770 688560 125860 688800
rect 126100 688560 126210 688800
rect 126450 688560 126540 688800
rect 126780 688560 126870 688800
rect 127110 688560 127200 688800
rect 127440 688560 127550 688800
rect 127790 688560 127880 688800
rect 128120 688560 128210 688800
rect 128450 688560 128540 688800
rect 128780 688560 128890 688800
rect 129130 688560 129220 688800
rect 129460 688560 129550 688800
rect 129790 688560 129880 688800
rect 130120 688560 130230 688800
rect 130470 688560 130560 688800
rect 130800 688560 130890 688800
rect 131130 688560 131220 688800
rect 131460 688560 131570 688800
rect 131810 688560 131900 688800
rect 132140 688560 132230 688800
rect 132470 688560 132560 688800
rect 132800 688560 132910 688800
rect 133150 688560 133570 688800
rect 133810 688560 133900 688800
rect 134140 688560 134230 688800
rect 134470 688560 134560 688800
rect 134800 688560 134910 688800
rect 135150 688560 135240 688800
rect 135480 688560 135570 688800
rect 135810 688560 135900 688800
rect 136140 688560 136250 688800
rect 136490 688560 136580 688800
rect 136820 688560 136910 688800
rect 137150 688560 137240 688800
rect 137480 688560 137590 688800
rect 137830 688560 137920 688800
rect 138160 688560 138250 688800
rect 138490 688560 138580 688800
rect 138820 688560 138930 688800
rect 139170 688560 139260 688800
rect 139500 688560 139590 688800
rect 139830 688560 139920 688800
rect 140160 688560 140270 688800
rect 140510 688560 140600 688800
rect 140840 688560 140930 688800
rect 141170 688560 141260 688800
rect 141500 688560 141610 688800
rect 141850 688560 141940 688800
rect 142180 688560 142270 688800
rect 142510 688560 142600 688800
rect 142840 688560 142950 688800
rect 143190 688560 143280 688800
rect 143520 688560 143610 688800
rect 143850 688560 143940 688800
rect 144180 688560 144290 688800
rect 144530 688560 144950 688800
rect 145190 688560 145280 688800
rect 145520 688560 145610 688800
rect 145850 688560 145940 688800
rect 146180 688560 146290 688800
rect 146530 688560 146620 688800
rect 146860 688560 146950 688800
rect 147190 688560 147280 688800
rect 147520 688560 147630 688800
rect 147870 688560 147960 688800
rect 148200 688560 148290 688800
rect 148530 688560 148620 688800
rect 148860 688560 148970 688800
rect 149210 688560 149300 688800
rect 149540 688560 149630 688800
rect 149870 688560 149960 688800
rect 150200 688560 150310 688800
rect 150550 688560 150640 688800
rect 150880 688560 150970 688800
rect 151210 688560 151300 688800
rect 151540 688560 151650 688800
rect 151890 688560 151980 688800
rect 152220 688560 152310 688800
rect 152550 688560 152640 688800
rect 152880 688560 152990 688800
rect 153230 688560 153320 688800
rect 153560 688560 153650 688800
rect 153890 688560 153980 688800
rect 154220 688560 154330 688800
rect 154570 688560 154660 688800
rect 154900 688560 154990 688800
rect 155230 688560 155320 688800
rect 155560 688560 155670 688800
rect 155910 688560 155960 688800
rect 110760 688470 155960 688560
rect 110760 688230 110810 688470
rect 111050 688230 111140 688470
rect 111380 688230 111470 688470
rect 111710 688230 111800 688470
rect 112040 688230 112150 688470
rect 112390 688230 112480 688470
rect 112720 688230 112810 688470
rect 113050 688230 113140 688470
rect 113380 688230 113490 688470
rect 113730 688230 113820 688470
rect 114060 688230 114150 688470
rect 114390 688230 114480 688470
rect 114720 688230 114830 688470
rect 115070 688230 115160 688470
rect 115400 688230 115490 688470
rect 115730 688230 115820 688470
rect 116060 688230 116170 688470
rect 116410 688230 116500 688470
rect 116740 688230 116830 688470
rect 117070 688230 117160 688470
rect 117400 688230 117510 688470
rect 117750 688230 117840 688470
rect 118080 688230 118170 688470
rect 118410 688230 118500 688470
rect 118740 688230 118850 688470
rect 119090 688230 119180 688470
rect 119420 688230 119510 688470
rect 119750 688230 119840 688470
rect 120080 688230 120190 688470
rect 120430 688230 120520 688470
rect 120760 688230 120850 688470
rect 121090 688230 121180 688470
rect 121420 688230 121530 688470
rect 121770 688230 122190 688470
rect 122430 688230 122520 688470
rect 122760 688230 122850 688470
rect 123090 688230 123180 688470
rect 123420 688230 123530 688470
rect 123770 688230 123860 688470
rect 124100 688230 124190 688470
rect 124430 688230 124520 688470
rect 124760 688230 124870 688470
rect 125110 688230 125200 688470
rect 125440 688230 125530 688470
rect 125770 688230 125860 688470
rect 126100 688230 126210 688470
rect 126450 688230 126540 688470
rect 126780 688230 126870 688470
rect 127110 688230 127200 688470
rect 127440 688230 127550 688470
rect 127790 688230 127880 688470
rect 128120 688230 128210 688470
rect 128450 688230 128540 688470
rect 128780 688230 128890 688470
rect 129130 688230 129220 688470
rect 129460 688230 129550 688470
rect 129790 688230 129880 688470
rect 130120 688230 130230 688470
rect 130470 688230 130560 688470
rect 130800 688230 130890 688470
rect 131130 688230 131220 688470
rect 131460 688230 131570 688470
rect 131810 688230 131900 688470
rect 132140 688230 132230 688470
rect 132470 688230 132560 688470
rect 132800 688230 132910 688470
rect 133150 688230 133570 688470
rect 133810 688230 133900 688470
rect 134140 688230 134230 688470
rect 134470 688230 134560 688470
rect 134800 688230 134910 688470
rect 135150 688230 135240 688470
rect 135480 688230 135570 688470
rect 135810 688230 135900 688470
rect 136140 688230 136250 688470
rect 136490 688230 136580 688470
rect 136820 688230 136910 688470
rect 137150 688230 137240 688470
rect 137480 688230 137590 688470
rect 137830 688230 137920 688470
rect 138160 688230 138250 688470
rect 138490 688230 138580 688470
rect 138820 688230 138930 688470
rect 139170 688230 139260 688470
rect 139500 688230 139590 688470
rect 139830 688230 139920 688470
rect 140160 688230 140270 688470
rect 140510 688230 140600 688470
rect 140840 688230 140930 688470
rect 141170 688230 141260 688470
rect 141500 688230 141610 688470
rect 141850 688230 141940 688470
rect 142180 688230 142270 688470
rect 142510 688230 142600 688470
rect 142840 688230 142950 688470
rect 143190 688230 143280 688470
rect 143520 688230 143610 688470
rect 143850 688230 143940 688470
rect 144180 688230 144290 688470
rect 144530 688230 144950 688470
rect 145190 688230 145280 688470
rect 145520 688230 145610 688470
rect 145850 688230 145940 688470
rect 146180 688230 146290 688470
rect 146530 688230 146620 688470
rect 146860 688230 146950 688470
rect 147190 688230 147280 688470
rect 147520 688230 147630 688470
rect 147870 688230 147960 688470
rect 148200 688230 148290 688470
rect 148530 688230 148620 688470
rect 148860 688230 148970 688470
rect 149210 688230 149300 688470
rect 149540 688230 149630 688470
rect 149870 688230 149960 688470
rect 150200 688230 150310 688470
rect 150550 688230 150640 688470
rect 150880 688230 150970 688470
rect 151210 688230 151300 688470
rect 151540 688230 151650 688470
rect 151890 688230 151980 688470
rect 152220 688230 152310 688470
rect 152550 688230 152640 688470
rect 152880 688230 152990 688470
rect 153230 688230 153320 688470
rect 153560 688230 153650 688470
rect 153890 688230 153980 688470
rect 154220 688230 154330 688470
rect 154570 688230 154660 688470
rect 154900 688230 154990 688470
rect 155230 688230 155320 688470
rect 155560 688230 155670 688470
rect 155910 688230 155960 688470
rect 110760 688140 155960 688230
rect 110760 687900 110810 688140
rect 111050 687900 111140 688140
rect 111380 687900 111470 688140
rect 111710 687900 111800 688140
rect 112040 687900 112150 688140
rect 112390 687900 112480 688140
rect 112720 687900 112810 688140
rect 113050 687900 113140 688140
rect 113380 687900 113490 688140
rect 113730 687900 113820 688140
rect 114060 687900 114150 688140
rect 114390 687900 114480 688140
rect 114720 687900 114830 688140
rect 115070 687900 115160 688140
rect 115400 687900 115490 688140
rect 115730 687900 115820 688140
rect 116060 687900 116170 688140
rect 116410 687900 116500 688140
rect 116740 687900 116830 688140
rect 117070 687900 117160 688140
rect 117400 687900 117510 688140
rect 117750 687900 117840 688140
rect 118080 687900 118170 688140
rect 118410 687900 118500 688140
rect 118740 687900 118850 688140
rect 119090 687900 119180 688140
rect 119420 687900 119510 688140
rect 119750 687900 119840 688140
rect 120080 687900 120190 688140
rect 120430 687900 120520 688140
rect 120760 687900 120850 688140
rect 121090 687900 121180 688140
rect 121420 687900 121530 688140
rect 121770 687900 122190 688140
rect 122430 687900 122520 688140
rect 122760 687900 122850 688140
rect 123090 687900 123180 688140
rect 123420 687900 123530 688140
rect 123770 687900 123860 688140
rect 124100 687900 124190 688140
rect 124430 687900 124520 688140
rect 124760 687900 124870 688140
rect 125110 687900 125200 688140
rect 125440 687900 125530 688140
rect 125770 687900 125860 688140
rect 126100 687900 126210 688140
rect 126450 687900 126540 688140
rect 126780 687900 126870 688140
rect 127110 687900 127200 688140
rect 127440 687900 127550 688140
rect 127790 687900 127880 688140
rect 128120 687900 128210 688140
rect 128450 687900 128540 688140
rect 128780 687900 128890 688140
rect 129130 687900 129220 688140
rect 129460 687900 129550 688140
rect 129790 687900 129880 688140
rect 130120 687900 130230 688140
rect 130470 687900 130560 688140
rect 130800 687900 130890 688140
rect 131130 687900 131220 688140
rect 131460 687900 131570 688140
rect 131810 687900 131900 688140
rect 132140 687900 132230 688140
rect 132470 687900 132560 688140
rect 132800 687900 132910 688140
rect 133150 687900 133570 688140
rect 133810 687900 133900 688140
rect 134140 687900 134230 688140
rect 134470 687900 134560 688140
rect 134800 687900 134910 688140
rect 135150 687900 135240 688140
rect 135480 687900 135570 688140
rect 135810 687900 135900 688140
rect 136140 687900 136250 688140
rect 136490 687900 136580 688140
rect 136820 687900 136910 688140
rect 137150 687900 137240 688140
rect 137480 687900 137590 688140
rect 137830 687900 137920 688140
rect 138160 687900 138250 688140
rect 138490 687900 138580 688140
rect 138820 687900 138930 688140
rect 139170 687900 139260 688140
rect 139500 687900 139590 688140
rect 139830 687900 139920 688140
rect 140160 687900 140270 688140
rect 140510 687900 140600 688140
rect 140840 687900 140930 688140
rect 141170 687900 141260 688140
rect 141500 687900 141610 688140
rect 141850 687900 141940 688140
rect 142180 687900 142270 688140
rect 142510 687900 142600 688140
rect 142840 687900 142950 688140
rect 143190 687900 143280 688140
rect 143520 687900 143610 688140
rect 143850 687900 143940 688140
rect 144180 687900 144290 688140
rect 144530 687900 144950 688140
rect 145190 687900 145280 688140
rect 145520 687900 145610 688140
rect 145850 687900 145940 688140
rect 146180 687900 146290 688140
rect 146530 687900 146620 688140
rect 146860 687900 146950 688140
rect 147190 687900 147280 688140
rect 147520 687900 147630 688140
rect 147870 687900 147960 688140
rect 148200 687900 148290 688140
rect 148530 687900 148620 688140
rect 148860 687900 148970 688140
rect 149210 687900 149300 688140
rect 149540 687900 149630 688140
rect 149870 687900 149960 688140
rect 150200 687900 150310 688140
rect 150550 687900 150640 688140
rect 150880 687900 150970 688140
rect 151210 687900 151300 688140
rect 151540 687900 151650 688140
rect 151890 687900 151980 688140
rect 152220 687900 152310 688140
rect 152550 687900 152640 688140
rect 152880 687900 152990 688140
rect 153230 687900 153320 688140
rect 153560 687900 153650 688140
rect 153890 687900 153980 688140
rect 154220 687900 154330 688140
rect 154570 687900 154660 688140
rect 154900 687900 154990 688140
rect 155230 687900 155320 688140
rect 155560 687900 155670 688140
rect 155910 687900 155960 688140
rect 110760 687790 155960 687900
rect 110760 687550 110810 687790
rect 111050 687550 111140 687790
rect 111380 687550 111470 687790
rect 111710 687550 111800 687790
rect 112040 687550 112150 687790
rect 112390 687550 112480 687790
rect 112720 687550 112810 687790
rect 113050 687550 113140 687790
rect 113380 687550 113490 687790
rect 113730 687550 113820 687790
rect 114060 687550 114150 687790
rect 114390 687550 114480 687790
rect 114720 687550 114830 687790
rect 115070 687550 115160 687790
rect 115400 687550 115490 687790
rect 115730 687550 115820 687790
rect 116060 687550 116170 687790
rect 116410 687550 116500 687790
rect 116740 687550 116830 687790
rect 117070 687550 117160 687790
rect 117400 687550 117510 687790
rect 117750 687550 117840 687790
rect 118080 687550 118170 687790
rect 118410 687550 118500 687790
rect 118740 687550 118850 687790
rect 119090 687550 119180 687790
rect 119420 687550 119510 687790
rect 119750 687550 119840 687790
rect 120080 687550 120190 687790
rect 120430 687550 120520 687790
rect 120760 687550 120850 687790
rect 121090 687550 121180 687790
rect 121420 687550 121530 687790
rect 121770 687550 122190 687790
rect 122430 687550 122520 687790
rect 122760 687550 122850 687790
rect 123090 687550 123180 687790
rect 123420 687550 123530 687790
rect 123770 687550 123860 687790
rect 124100 687550 124190 687790
rect 124430 687550 124520 687790
rect 124760 687550 124870 687790
rect 125110 687550 125200 687790
rect 125440 687550 125530 687790
rect 125770 687550 125860 687790
rect 126100 687550 126210 687790
rect 126450 687550 126540 687790
rect 126780 687550 126870 687790
rect 127110 687550 127200 687790
rect 127440 687550 127550 687790
rect 127790 687550 127880 687790
rect 128120 687550 128210 687790
rect 128450 687550 128540 687790
rect 128780 687550 128890 687790
rect 129130 687550 129220 687790
rect 129460 687550 129550 687790
rect 129790 687550 129880 687790
rect 130120 687550 130230 687790
rect 130470 687550 130560 687790
rect 130800 687550 130890 687790
rect 131130 687550 131220 687790
rect 131460 687550 131570 687790
rect 131810 687550 131900 687790
rect 132140 687550 132230 687790
rect 132470 687550 132560 687790
rect 132800 687550 132910 687790
rect 133150 687550 133570 687790
rect 133810 687550 133900 687790
rect 134140 687550 134230 687790
rect 134470 687550 134560 687790
rect 134800 687550 134910 687790
rect 135150 687550 135240 687790
rect 135480 687550 135570 687790
rect 135810 687550 135900 687790
rect 136140 687550 136250 687790
rect 136490 687550 136580 687790
rect 136820 687550 136910 687790
rect 137150 687550 137240 687790
rect 137480 687550 137590 687790
rect 137830 687550 137920 687790
rect 138160 687550 138250 687790
rect 138490 687550 138580 687790
rect 138820 687550 138930 687790
rect 139170 687550 139260 687790
rect 139500 687550 139590 687790
rect 139830 687550 139920 687790
rect 140160 687550 140270 687790
rect 140510 687550 140600 687790
rect 140840 687550 140930 687790
rect 141170 687550 141260 687790
rect 141500 687550 141610 687790
rect 141850 687550 141940 687790
rect 142180 687550 142270 687790
rect 142510 687550 142600 687790
rect 142840 687550 142950 687790
rect 143190 687550 143280 687790
rect 143520 687550 143610 687790
rect 143850 687550 143940 687790
rect 144180 687550 144290 687790
rect 144530 687550 144950 687790
rect 145190 687550 145280 687790
rect 145520 687550 145610 687790
rect 145850 687550 145940 687790
rect 146180 687550 146290 687790
rect 146530 687550 146620 687790
rect 146860 687550 146950 687790
rect 147190 687550 147280 687790
rect 147520 687550 147630 687790
rect 147870 687550 147960 687790
rect 148200 687550 148290 687790
rect 148530 687550 148620 687790
rect 148860 687550 148970 687790
rect 149210 687550 149300 687790
rect 149540 687550 149630 687790
rect 149870 687550 149960 687790
rect 150200 687550 150310 687790
rect 150550 687550 150640 687790
rect 150880 687550 150970 687790
rect 151210 687550 151300 687790
rect 151540 687550 151650 687790
rect 151890 687550 151980 687790
rect 152220 687550 152310 687790
rect 152550 687550 152640 687790
rect 152880 687550 152990 687790
rect 153230 687550 153320 687790
rect 153560 687550 153650 687790
rect 153890 687550 153980 687790
rect 154220 687550 154330 687790
rect 154570 687550 154660 687790
rect 154900 687550 154990 687790
rect 155230 687550 155320 687790
rect 155560 687550 155670 687790
rect 155910 687550 155960 687790
rect 110760 687460 155960 687550
rect 110760 687220 110810 687460
rect 111050 687220 111140 687460
rect 111380 687220 111470 687460
rect 111710 687220 111800 687460
rect 112040 687220 112150 687460
rect 112390 687220 112480 687460
rect 112720 687220 112810 687460
rect 113050 687220 113140 687460
rect 113380 687220 113490 687460
rect 113730 687220 113820 687460
rect 114060 687220 114150 687460
rect 114390 687220 114480 687460
rect 114720 687220 114830 687460
rect 115070 687220 115160 687460
rect 115400 687220 115490 687460
rect 115730 687220 115820 687460
rect 116060 687220 116170 687460
rect 116410 687220 116500 687460
rect 116740 687220 116830 687460
rect 117070 687220 117160 687460
rect 117400 687220 117510 687460
rect 117750 687220 117840 687460
rect 118080 687220 118170 687460
rect 118410 687220 118500 687460
rect 118740 687220 118850 687460
rect 119090 687220 119180 687460
rect 119420 687220 119510 687460
rect 119750 687220 119840 687460
rect 120080 687220 120190 687460
rect 120430 687220 120520 687460
rect 120760 687220 120850 687460
rect 121090 687220 121180 687460
rect 121420 687220 121530 687460
rect 121770 687220 122190 687460
rect 122430 687220 122520 687460
rect 122760 687220 122850 687460
rect 123090 687220 123180 687460
rect 123420 687220 123530 687460
rect 123770 687220 123860 687460
rect 124100 687220 124190 687460
rect 124430 687220 124520 687460
rect 124760 687220 124870 687460
rect 125110 687220 125200 687460
rect 125440 687220 125530 687460
rect 125770 687220 125860 687460
rect 126100 687220 126210 687460
rect 126450 687220 126540 687460
rect 126780 687220 126870 687460
rect 127110 687220 127200 687460
rect 127440 687220 127550 687460
rect 127790 687220 127880 687460
rect 128120 687220 128210 687460
rect 128450 687220 128540 687460
rect 128780 687220 128890 687460
rect 129130 687220 129220 687460
rect 129460 687220 129550 687460
rect 129790 687220 129880 687460
rect 130120 687220 130230 687460
rect 130470 687220 130560 687460
rect 130800 687220 130890 687460
rect 131130 687220 131220 687460
rect 131460 687220 131570 687460
rect 131810 687220 131900 687460
rect 132140 687220 132230 687460
rect 132470 687220 132560 687460
rect 132800 687220 132910 687460
rect 133150 687220 133570 687460
rect 133810 687220 133900 687460
rect 134140 687220 134230 687460
rect 134470 687220 134560 687460
rect 134800 687220 134910 687460
rect 135150 687220 135240 687460
rect 135480 687220 135570 687460
rect 135810 687220 135900 687460
rect 136140 687220 136250 687460
rect 136490 687220 136580 687460
rect 136820 687220 136910 687460
rect 137150 687220 137240 687460
rect 137480 687220 137590 687460
rect 137830 687220 137920 687460
rect 138160 687220 138250 687460
rect 138490 687220 138580 687460
rect 138820 687220 138930 687460
rect 139170 687220 139260 687460
rect 139500 687220 139590 687460
rect 139830 687220 139920 687460
rect 140160 687220 140270 687460
rect 140510 687220 140600 687460
rect 140840 687220 140930 687460
rect 141170 687220 141260 687460
rect 141500 687220 141610 687460
rect 141850 687220 141940 687460
rect 142180 687220 142270 687460
rect 142510 687220 142600 687460
rect 142840 687220 142950 687460
rect 143190 687220 143280 687460
rect 143520 687220 143610 687460
rect 143850 687220 143940 687460
rect 144180 687220 144290 687460
rect 144530 687220 144950 687460
rect 145190 687220 145280 687460
rect 145520 687220 145610 687460
rect 145850 687220 145940 687460
rect 146180 687220 146290 687460
rect 146530 687220 146620 687460
rect 146860 687220 146950 687460
rect 147190 687220 147280 687460
rect 147520 687220 147630 687460
rect 147870 687220 147960 687460
rect 148200 687220 148290 687460
rect 148530 687220 148620 687460
rect 148860 687220 148970 687460
rect 149210 687220 149300 687460
rect 149540 687220 149630 687460
rect 149870 687220 149960 687460
rect 150200 687220 150310 687460
rect 150550 687220 150640 687460
rect 150880 687220 150970 687460
rect 151210 687220 151300 687460
rect 151540 687220 151650 687460
rect 151890 687220 151980 687460
rect 152220 687220 152310 687460
rect 152550 687220 152640 687460
rect 152880 687220 152990 687460
rect 153230 687220 153320 687460
rect 153560 687220 153650 687460
rect 153890 687220 153980 687460
rect 154220 687220 154330 687460
rect 154570 687220 154660 687460
rect 154900 687220 154990 687460
rect 155230 687220 155320 687460
rect 155560 687220 155670 687460
rect 155910 687220 155960 687460
rect 110760 687130 155960 687220
rect 110760 686890 110810 687130
rect 111050 686890 111140 687130
rect 111380 686890 111470 687130
rect 111710 686890 111800 687130
rect 112040 686890 112150 687130
rect 112390 686890 112480 687130
rect 112720 686890 112810 687130
rect 113050 686890 113140 687130
rect 113380 686890 113490 687130
rect 113730 686890 113820 687130
rect 114060 686890 114150 687130
rect 114390 686890 114480 687130
rect 114720 686890 114830 687130
rect 115070 686890 115160 687130
rect 115400 686890 115490 687130
rect 115730 686890 115820 687130
rect 116060 686890 116170 687130
rect 116410 686890 116500 687130
rect 116740 686890 116830 687130
rect 117070 686890 117160 687130
rect 117400 686890 117510 687130
rect 117750 686890 117840 687130
rect 118080 686890 118170 687130
rect 118410 686890 118500 687130
rect 118740 686890 118850 687130
rect 119090 686890 119180 687130
rect 119420 686890 119510 687130
rect 119750 686890 119840 687130
rect 120080 686890 120190 687130
rect 120430 686890 120520 687130
rect 120760 686890 120850 687130
rect 121090 686890 121180 687130
rect 121420 686890 121530 687130
rect 121770 686890 122190 687130
rect 122430 686890 122520 687130
rect 122760 686890 122850 687130
rect 123090 686890 123180 687130
rect 123420 686890 123530 687130
rect 123770 686890 123860 687130
rect 124100 686890 124190 687130
rect 124430 686890 124520 687130
rect 124760 686890 124870 687130
rect 125110 686890 125200 687130
rect 125440 686890 125530 687130
rect 125770 686890 125860 687130
rect 126100 686890 126210 687130
rect 126450 686890 126540 687130
rect 126780 686890 126870 687130
rect 127110 686890 127200 687130
rect 127440 686890 127550 687130
rect 127790 686890 127880 687130
rect 128120 686890 128210 687130
rect 128450 686890 128540 687130
rect 128780 686890 128890 687130
rect 129130 686890 129220 687130
rect 129460 686890 129550 687130
rect 129790 686890 129880 687130
rect 130120 686890 130230 687130
rect 130470 686890 130560 687130
rect 130800 686890 130890 687130
rect 131130 686890 131220 687130
rect 131460 686890 131570 687130
rect 131810 686890 131900 687130
rect 132140 686890 132230 687130
rect 132470 686890 132560 687130
rect 132800 686890 132910 687130
rect 133150 686890 133570 687130
rect 133810 686890 133900 687130
rect 134140 686890 134230 687130
rect 134470 686890 134560 687130
rect 134800 686890 134910 687130
rect 135150 686890 135240 687130
rect 135480 686890 135570 687130
rect 135810 686890 135900 687130
rect 136140 686890 136250 687130
rect 136490 686890 136580 687130
rect 136820 686890 136910 687130
rect 137150 686890 137240 687130
rect 137480 686890 137590 687130
rect 137830 686890 137920 687130
rect 138160 686890 138250 687130
rect 138490 686890 138580 687130
rect 138820 686890 138930 687130
rect 139170 686890 139260 687130
rect 139500 686890 139590 687130
rect 139830 686890 139920 687130
rect 140160 686890 140270 687130
rect 140510 686890 140600 687130
rect 140840 686890 140930 687130
rect 141170 686890 141260 687130
rect 141500 686890 141610 687130
rect 141850 686890 141940 687130
rect 142180 686890 142270 687130
rect 142510 686890 142600 687130
rect 142840 686890 142950 687130
rect 143190 686890 143280 687130
rect 143520 686890 143610 687130
rect 143850 686890 143940 687130
rect 144180 686890 144290 687130
rect 144530 686890 144950 687130
rect 145190 686890 145280 687130
rect 145520 686890 145610 687130
rect 145850 686890 145940 687130
rect 146180 686890 146290 687130
rect 146530 686890 146620 687130
rect 146860 686890 146950 687130
rect 147190 686890 147280 687130
rect 147520 686890 147630 687130
rect 147870 686890 147960 687130
rect 148200 686890 148290 687130
rect 148530 686890 148620 687130
rect 148860 686890 148970 687130
rect 149210 686890 149300 687130
rect 149540 686890 149630 687130
rect 149870 686890 149960 687130
rect 150200 686890 150310 687130
rect 150550 686890 150640 687130
rect 150880 686890 150970 687130
rect 151210 686890 151300 687130
rect 151540 686890 151650 687130
rect 151890 686890 151980 687130
rect 152220 686890 152310 687130
rect 152550 686890 152640 687130
rect 152880 686890 152990 687130
rect 153230 686890 153320 687130
rect 153560 686890 153650 687130
rect 153890 686890 153980 687130
rect 154220 686890 154330 687130
rect 154570 686890 154660 687130
rect 154900 686890 154990 687130
rect 155230 686890 155320 687130
rect 155560 686890 155670 687130
rect 155910 686890 155960 687130
rect 110760 686800 155960 686890
rect 110760 686560 110810 686800
rect 111050 686560 111140 686800
rect 111380 686560 111470 686800
rect 111710 686560 111800 686800
rect 112040 686560 112150 686800
rect 112390 686560 112480 686800
rect 112720 686560 112810 686800
rect 113050 686560 113140 686800
rect 113380 686560 113490 686800
rect 113730 686560 113820 686800
rect 114060 686560 114150 686800
rect 114390 686560 114480 686800
rect 114720 686560 114830 686800
rect 115070 686560 115160 686800
rect 115400 686560 115490 686800
rect 115730 686560 115820 686800
rect 116060 686560 116170 686800
rect 116410 686560 116500 686800
rect 116740 686560 116830 686800
rect 117070 686560 117160 686800
rect 117400 686560 117510 686800
rect 117750 686560 117840 686800
rect 118080 686560 118170 686800
rect 118410 686560 118500 686800
rect 118740 686560 118850 686800
rect 119090 686560 119180 686800
rect 119420 686560 119510 686800
rect 119750 686560 119840 686800
rect 120080 686560 120190 686800
rect 120430 686560 120520 686800
rect 120760 686560 120850 686800
rect 121090 686560 121180 686800
rect 121420 686560 121530 686800
rect 121770 686560 122190 686800
rect 122430 686560 122520 686800
rect 122760 686560 122850 686800
rect 123090 686560 123180 686800
rect 123420 686560 123530 686800
rect 123770 686560 123860 686800
rect 124100 686560 124190 686800
rect 124430 686560 124520 686800
rect 124760 686560 124870 686800
rect 125110 686560 125200 686800
rect 125440 686560 125530 686800
rect 125770 686560 125860 686800
rect 126100 686560 126210 686800
rect 126450 686560 126540 686800
rect 126780 686560 126870 686800
rect 127110 686560 127200 686800
rect 127440 686560 127550 686800
rect 127790 686560 127880 686800
rect 128120 686560 128210 686800
rect 128450 686560 128540 686800
rect 128780 686560 128890 686800
rect 129130 686560 129220 686800
rect 129460 686560 129550 686800
rect 129790 686560 129880 686800
rect 130120 686560 130230 686800
rect 130470 686560 130560 686800
rect 130800 686560 130890 686800
rect 131130 686560 131220 686800
rect 131460 686560 131570 686800
rect 131810 686560 131900 686800
rect 132140 686560 132230 686800
rect 132470 686560 132560 686800
rect 132800 686560 132910 686800
rect 133150 686560 133570 686800
rect 133810 686560 133900 686800
rect 134140 686560 134230 686800
rect 134470 686560 134560 686800
rect 134800 686560 134910 686800
rect 135150 686560 135240 686800
rect 135480 686560 135570 686800
rect 135810 686560 135900 686800
rect 136140 686560 136250 686800
rect 136490 686560 136580 686800
rect 136820 686560 136910 686800
rect 137150 686560 137240 686800
rect 137480 686560 137590 686800
rect 137830 686560 137920 686800
rect 138160 686560 138250 686800
rect 138490 686560 138580 686800
rect 138820 686560 138930 686800
rect 139170 686560 139260 686800
rect 139500 686560 139590 686800
rect 139830 686560 139920 686800
rect 140160 686560 140270 686800
rect 140510 686560 140600 686800
rect 140840 686560 140930 686800
rect 141170 686560 141260 686800
rect 141500 686560 141610 686800
rect 141850 686560 141940 686800
rect 142180 686560 142270 686800
rect 142510 686560 142600 686800
rect 142840 686560 142950 686800
rect 143190 686560 143280 686800
rect 143520 686560 143610 686800
rect 143850 686560 143940 686800
rect 144180 686560 144290 686800
rect 144530 686560 144950 686800
rect 145190 686560 145280 686800
rect 145520 686560 145610 686800
rect 145850 686560 145940 686800
rect 146180 686560 146290 686800
rect 146530 686560 146620 686800
rect 146860 686560 146950 686800
rect 147190 686560 147280 686800
rect 147520 686560 147630 686800
rect 147870 686560 147960 686800
rect 148200 686560 148290 686800
rect 148530 686560 148620 686800
rect 148860 686560 148970 686800
rect 149210 686560 149300 686800
rect 149540 686560 149630 686800
rect 149870 686560 149960 686800
rect 150200 686560 150310 686800
rect 150550 686560 150640 686800
rect 150880 686560 150970 686800
rect 151210 686560 151300 686800
rect 151540 686560 151650 686800
rect 151890 686560 151980 686800
rect 152220 686560 152310 686800
rect 152550 686560 152640 686800
rect 152880 686560 152990 686800
rect 153230 686560 153320 686800
rect 153560 686560 153650 686800
rect 153890 686560 153980 686800
rect 154220 686560 154330 686800
rect 154570 686560 154660 686800
rect 154900 686560 154990 686800
rect 155230 686560 155320 686800
rect 155560 686560 155670 686800
rect 155910 686560 155960 686800
rect 110760 686450 155960 686560
rect 110760 686210 110810 686450
rect 111050 686210 111140 686450
rect 111380 686210 111470 686450
rect 111710 686210 111800 686450
rect 112040 686210 112150 686450
rect 112390 686210 112480 686450
rect 112720 686210 112810 686450
rect 113050 686210 113140 686450
rect 113380 686210 113490 686450
rect 113730 686210 113820 686450
rect 114060 686210 114150 686450
rect 114390 686210 114480 686450
rect 114720 686210 114830 686450
rect 115070 686210 115160 686450
rect 115400 686210 115490 686450
rect 115730 686210 115820 686450
rect 116060 686210 116170 686450
rect 116410 686210 116500 686450
rect 116740 686210 116830 686450
rect 117070 686210 117160 686450
rect 117400 686210 117510 686450
rect 117750 686210 117840 686450
rect 118080 686210 118170 686450
rect 118410 686210 118500 686450
rect 118740 686210 118850 686450
rect 119090 686210 119180 686450
rect 119420 686210 119510 686450
rect 119750 686210 119840 686450
rect 120080 686210 120190 686450
rect 120430 686210 120520 686450
rect 120760 686210 120850 686450
rect 121090 686210 121180 686450
rect 121420 686210 121530 686450
rect 121770 686210 122190 686450
rect 122430 686210 122520 686450
rect 122760 686210 122850 686450
rect 123090 686210 123180 686450
rect 123420 686210 123530 686450
rect 123770 686210 123860 686450
rect 124100 686210 124190 686450
rect 124430 686210 124520 686450
rect 124760 686210 124870 686450
rect 125110 686210 125200 686450
rect 125440 686210 125530 686450
rect 125770 686210 125860 686450
rect 126100 686210 126210 686450
rect 126450 686210 126540 686450
rect 126780 686210 126870 686450
rect 127110 686210 127200 686450
rect 127440 686210 127550 686450
rect 127790 686210 127880 686450
rect 128120 686210 128210 686450
rect 128450 686210 128540 686450
rect 128780 686210 128890 686450
rect 129130 686210 129220 686450
rect 129460 686210 129550 686450
rect 129790 686210 129880 686450
rect 130120 686210 130230 686450
rect 130470 686210 130560 686450
rect 130800 686210 130890 686450
rect 131130 686210 131220 686450
rect 131460 686210 131570 686450
rect 131810 686210 131900 686450
rect 132140 686210 132230 686450
rect 132470 686210 132560 686450
rect 132800 686210 132910 686450
rect 133150 686210 133570 686450
rect 133810 686210 133900 686450
rect 134140 686210 134230 686450
rect 134470 686210 134560 686450
rect 134800 686210 134910 686450
rect 135150 686210 135240 686450
rect 135480 686210 135570 686450
rect 135810 686210 135900 686450
rect 136140 686210 136250 686450
rect 136490 686210 136580 686450
rect 136820 686210 136910 686450
rect 137150 686210 137240 686450
rect 137480 686210 137590 686450
rect 137830 686210 137920 686450
rect 138160 686210 138250 686450
rect 138490 686210 138580 686450
rect 138820 686210 138930 686450
rect 139170 686210 139260 686450
rect 139500 686210 139590 686450
rect 139830 686210 139920 686450
rect 140160 686210 140270 686450
rect 140510 686210 140600 686450
rect 140840 686210 140930 686450
rect 141170 686210 141260 686450
rect 141500 686210 141610 686450
rect 141850 686210 141940 686450
rect 142180 686210 142270 686450
rect 142510 686210 142600 686450
rect 142840 686210 142950 686450
rect 143190 686210 143280 686450
rect 143520 686210 143610 686450
rect 143850 686210 143940 686450
rect 144180 686210 144290 686450
rect 144530 686210 144950 686450
rect 145190 686210 145280 686450
rect 145520 686210 145610 686450
rect 145850 686210 145940 686450
rect 146180 686210 146290 686450
rect 146530 686210 146620 686450
rect 146860 686210 146950 686450
rect 147190 686210 147280 686450
rect 147520 686210 147630 686450
rect 147870 686210 147960 686450
rect 148200 686210 148290 686450
rect 148530 686210 148620 686450
rect 148860 686210 148970 686450
rect 149210 686210 149300 686450
rect 149540 686210 149630 686450
rect 149870 686210 149960 686450
rect 150200 686210 150310 686450
rect 150550 686210 150640 686450
rect 150880 686210 150970 686450
rect 151210 686210 151300 686450
rect 151540 686210 151650 686450
rect 151890 686210 151980 686450
rect 152220 686210 152310 686450
rect 152550 686210 152640 686450
rect 152880 686210 152990 686450
rect 153230 686210 153320 686450
rect 153560 686210 153650 686450
rect 153890 686210 153980 686450
rect 154220 686210 154330 686450
rect 154570 686210 154660 686450
rect 154900 686210 154990 686450
rect 155230 686210 155320 686450
rect 155560 686210 155670 686450
rect 155910 686210 155960 686450
rect 110760 686120 155960 686210
rect 110760 685880 110810 686120
rect 111050 685880 111140 686120
rect 111380 685880 111470 686120
rect 111710 685880 111800 686120
rect 112040 685880 112150 686120
rect 112390 685880 112480 686120
rect 112720 685880 112810 686120
rect 113050 685880 113140 686120
rect 113380 685880 113490 686120
rect 113730 685880 113820 686120
rect 114060 685880 114150 686120
rect 114390 685880 114480 686120
rect 114720 685880 114830 686120
rect 115070 685880 115160 686120
rect 115400 685880 115490 686120
rect 115730 685880 115820 686120
rect 116060 685880 116170 686120
rect 116410 685880 116500 686120
rect 116740 685880 116830 686120
rect 117070 685880 117160 686120
rect 117400 685880 117510 686120
rect 117750 685880 117840 686120
rect 118080 685880 118170 686120
rect 118410 685880 118500 686120
rect 118740 685880 118850 686120
rect 119090 685880 119180 686120
rect 119420 685880 119510 686120
rect 119750 685880 119840 686120
rect 120080 685880 120190 686120
rect 120430 685880 120520 686120
rect 120760 685880 120850 686120
rect 121090 685880 121180 686120
rect 121420 685880 121530 686120
rect 121770 685880 122190 686120
rect 122430 685880 122520 686120
rect 122760 685880 122850 686120
rect 123090 685880 123180 686120
rect 123420 685880 123530 686120
rect 123770 685880 123860 686120
rect 124100 685880 124190 686120
rect 124430 685880 124520 686120
rect 124760 685880 124870 686120
rect 125110 685880 125200 686120
rect 125440 685880 125530 686120
rect 125770 685880 125860 686120
rect 126100 685880 126210 686120
rect 126450 685880 126540 686120
rect 126780 685880 126870 686120
rect 127110 685880 127200 686120
rect 127440 685880 127550 686120
rect 127790 685880 127880 686120
rect 128120 685880 128210 686120
rect 128450 685880 128540 686120
rect 128780 685880 128890 686120
rect 129130 685880 129220 686120
rect 129460 685880 129550 686120
rect 129790 685880 129880 686120
rect 130120 685880 130230 686120
rect 130470 685880 130560 686120
rect 130800 685880 130890 686120
rect 131130 685880 131220 686120
rect 131460 685880 131570 686120
rect 131810 685880 131900 686120
rect 132140 685880 132230 686120
rect 132470 685880 132560 686120
rect 132800 685880 132910 686120
rect 133150 685880 133570 686120
rect 133810 685880 133900 686120
rect 134140 685880 134230 686120
rect 134470 685880 134560 686120
rect 134800 685880 134910 686120
rect 135150 685880 135240 686120
rect 135480 685880 135570 686120
rect 135810 685880 135900 686120
rect 136140 685880 136250 686120
rect 136490 685880 136580 686120
rect 136820 685880 136910 686120
rect 137150 685880 137240 686120
rect 137480 685880 137590 686120
rect 137830 685880 137920 686120
rect 138160 685880 138250 686120
rect 138490 685880 138580 686120
rect 138820 685880 138930 686120
rect 139170 685880 139260 686120
rect 139500 685880 139590 686120
rect 139830 685880 139920 686120
rect 140160 685880 140270 686120
rect 140510 685880 140600 686120
rect 140840 685880 140930 686120
rect 141170 685880 141260 686120
rect 141500 685880 141610 686120
rect 141850 685880 141940 686120
rect 142180 685880 142270 686120
rect 142510 685880 142600 686120
rect 142840 685880 142950 686120
rect 143190 685880 143280 686120
rect 143520 685880 143610 686120
rect 143850 685880 143940 686120
rect 144180 685880 144290 686120
rect 144530 685880 144950 686120
rect 145190 685880 145280 686120
rect 145520 685880 145610 686120
rect 145850 685880 145940 686120
rect 146180 685880 146290 686120
rect 146530 685880 146620 686120
rect 146860 685880 146950 686120
rect 147190 685880 147280 686120
rect 147520 685880 147630 686120
rect 147870 685880 147960 686120
rect 148200 685880 148290 686120
rect 148530 685880 148620 686120
rect 148860 685880 148970 686120
rect 149210 685880 149300 686120
rect 149540 685880 149630 686120
rect 149870 685880 149960 686120
rect 150200 685880 150310 686120
rect 150550 685880 150640 686120
rect 150880 685880 150970 686120
rect 151210 685880 151300 686120
rect 151540 685880 151650 686120
rect 151890 685880 151980 686120
rect 152220 685880 152310 686120
rect 152550 685880 152640 686120
rect 152880 685880 152990 686120
rect 153230 685880 153320 686120
rect 153560 685880 153650 686120
rect 153890 685880 153980 686120
rect 154220 685880 154330 686120
rect 154570 685880 154660 686120
rect 154900 685880 154990 686120
rect 155230 685880 155320 686120
rect 155560 685880 155670 686120
rect 155910 685880 155960 686120
rect 110760 685790 155960 685880
rect 110760 685550 110810 685790
rect 111050 685550 111140 685790
rect 111380 685550 111470 685790
rect 111710 685550 111800 685790
rect 112040 685550 112150 685790
rect 112390 685550 112480 685790
rect 112720 685550 112810 685790
rect 113050 685550 113140 685790
rect 113380 685550 113490 685790
rect 113730 685550 113820 685790
rect 114060 685550 114150 685790
rect 114390 685550 114480 685790
rect 114720 685550 114830 685790
rect 115070 685550 115160 685790
rect 115400 685550 115490 685790
rect 115730 685550 115820 685790
rect 116060 685550 116170 685790
rect 116410 685550 116500 685790
rect 116740 685550 116830 685790
rect 117070 685550 117160 685790
rect 117400 685550 117510 685790
rect 117750 685550 117840 685790
rect 118080 685550 118170 685790
rect 118410 685550 118500 685790
rect 118740 685550 118850 685790
rect 119090 685550 119180 685790
rect 119420 685550 119510 685790
rect 119750 685550 119840 685790
rect 120080 685550 120190 685790
rect 120430 685550 120520 685790
rect 120760 685550 120850 685790
rect 121090 685550 121180 685790
rect 121420 685550 121530 685790
rect 121770 685550 122190 685790
rect 122430 685550 122520 685790
rect 122760 685550 122850 685790
rect 123090 685550 123180 685790
rect 123420 685550 123530 685790
rect 123770 685550 123860 685790
rect 124100 685550 124190 685790
rect 124430 685550 124520 685790
rect 124760 685550 124870 685790
rect 125110 685550 125200 685790
rect 125440 685550 125530 685790
rect 125770 685550 125860 685790
rect 126100 685550 126210 685790
rect 126450 685550 126540 685790
rect 126780 685550 126870 685790
rect 127110 685550 127200 685790
rect 127440 685550 127550 685790
rect 127790 685550 127880 685790
rect 128120 685550 128210 685790
rect 128450 685550 128540 685790
rect 128780 685550 128890 685790
rect 129130 685550 129220 685790
rect 129460 685550 129550 685790
rect 129790 685550 129880 685790
rect 130120 685550 130230 685790
rect 130470 685550 130560 685790
rect 130800 685550 130890 685790
rect 131130 685550 131220 685790
rect 131460 685550 131570 685790
rect 131810 685550 131900 685790
rect 132140 685550 132230 685790
rect 132470 685550 132560 685790
rect 132800 685550 132910 685790
rect 133150 685550 133570 685790
rect 133810 685550 133900 685790
rect 134140 685550 134230 685790
rect 134470 685550 134560 685790
rect 134800 685550 134910 685790
rect 135150 685550 135240 685790
rect 135480 685550 135570 685790
rect 135810 685550 135900 685790
rect 136140 685550 136250 685790
rect 136490 685550 136580 685790
rect 136820 685550 136910 685790
rect 137150 685550 137240 685790
rect 137480 685550 137590 685790
rect 137830 685550 137920 685790
rect 138160 685550 138250 685790
rect 138490 685550 138580 685790
rect 138820 685550 138930 685790
rect 139170 685550 139260 685790
rect 139500 685550 139590 685790
rect 139830 685550 139920 685790
rect 140160 685550 140270 685790
rect 140510 685550 140600 685790
rect 140840 685550 140930 685790
rect 141170 685550 141260 685790
rect 141500 685550 141610 685790
rect 141850 685550 141940 685790
rect 142180 685550 142270 685790
rect 142510 685550 142600 685790
rect 142840 685550 142950 685790
rect 143190 685550 143280 685790
rect 143520 685550 143610 685790
rect 143850 685550 143940 685790
rect 144180 685550 144290 685790
rect 144530 685550 144950 685790
rect 145190 685550 145280 685790
rect 145520 685550 145610 685790
rect 145850 685550 145940 685790
rect 146180 685550 146290 685790
rect 146530 685550 146620 685790
rect 146860 685550 146950 685790
rect 147190 685550 147280 685790
rect 147520 685550 147630 685790
rect 147870 685550 147960 685790
rect 148200 685550 148290 685790
rect 148530 685550 148620 685790
rect 148860 685550 148970 685790
rect 149210 685550 149300 685790
rect 149540 685550 149630 685790
rect 149870 685550 149960 685790
rect 150200 685550 150310 685790
rect 150550 685550 150640 685790
rect 150880 685550 150970 685790
rect 151210 685550 151300 685790
rect 151540 685550 151650 685790
rect 151890 685550 151980 685790
rect 152220 685550 152310 685790
rect 152550 685550 152640 685790
rect 152880 685550 152990 685790
rect 153230 685550 153320 685790
rect 153560 685550 153650 685790
rect 153890 685550 153980 685790
rect 154220 685550 154330 685790
rect 154570 685550 154660 685790
rect 154900 685550 154990 685790
rect 155230 685550 155320 685790
rect 155560 685550 155670 685790
rect 155910 685550 155960 685790
rect 110760 685460 155960 685550
rect 110760 685220 110810 685460
rect 111050 685220 111140 685460
rect 111380 685220 111470 685460
rect 111710 685220 111800 685460
rect 112040 685220 112150 685460
rect 112390 685220 112480 685460
rect 112720 685220 112810 685460
rect 113050 685220 113140 685460
rect 113380 685220 113490 685460
rect 113730 685220 113820 685460
rect 114060 685220 114150 685460
rect 114390 685220 114480 685460
rect 114720 685220 114830 685460
rect 115070 685220 115160 685460
rect 115400 685220 115490 685460
rect 115730 685220 115820 685460
rect 116060 685220 116170 685460
rect 116410 685220 116500 685460
rect 116740 685220 116830 685460
rect 117070 685220 117160 685460
rect 117400 685220 117510 685460
rect 117750 685220 117840 685460
rect 118080 685220 118170 685460
rect 118410 685220 118500 685460
rect 118740 685220 118850 685460
rect 119090 685220 119180 685460
rect 119420 685220 119510 685460
rect 119750 685220 119840 685460
rect 120080 685220 120190 685460
rect 120430 685220 120520 685460
rect 120760 685220 120850 685460
rect 121090 685220 121180 685460
rect 121420 685220 121530 685460
rect 121770 685220 122190 685460
rect 122430 685220 122520 685460
rect 122760 685220 122850 685460
rect 123090 685220 123180 685460
rect 123420 685220 123530 685460
rect 123770 685220 123860 685460
rect 124100 685220 124190 685460
rect 124430 685220 124520 685460
rect 124760 685220 124870 685460
rect 125110 685220 125200 685460
rect 125440 685220 125530 685460
rect 125770 685220 125860 685460
rect 126100 685220 126210 685460
rect 126450 685220 126540 685460
rect 126780 685220 126870 685460
rect 127110 685220 127200 685460
rect 127440 685220 127550 685460
rect 127790 685220 127880 685460
rect 128120 685220 128210 685460
rect 128450 685220 128540 685460
rect 128780 685220 128890 685460
rect 129130 685220 129220 685460
rect 129460 685220 129550 685460
rect 129790 685220 129880 685460
rect 130120 685220 130230 685460
rect 130470 685220 130560 685460
rect 130800 685220 130890 685460
rect 131130 685220 131220 685460
rect 131460 685220 131570 685460
rect 131810 685220 131900 685460
rect 132140 685220 132230 685460
rect 132470 685220 132560 685460
rect 132800 685220 132910 685460
rect 133150 685220 133570 685460
rect 133810 685220 133900 685460
rect 134140 685220 134230 685460
rect 134470 685220 134560 685460
rect 134800 685220 134910 685460
rect 135150 685220 135240 685460
rect 135480 685220 135570 685460
rect 135810 685220 135900 685460
rect 136140 685220 136250 685460
rect 136490 685220 136580 685460
rect 136820 685220 136910 685460
rect 137150 685220 137240 685460
rect 137480 685220 137590 685460
rect 137830 685220 137920 685460
rect 138160 685220 138250 685460
rect 138490 685220 138580 685460
rect 138820 685220 138930 685460
rect 139170 685220 139260 685460
rect 139500 685220 139590 685460
rect 139830 685220 139920 685460
rect 140160 685220 140270 685460
rect 140510 685220 140600 685460
rect 140840 685220 140930 685460
rect 141170 685220 141260 685460
rect 141500 685220 141610 685460
rect 141850 685220 141940 685460
rect 142180 685220 142270 685460
rect 142510 685220 142600 685460
rect 142840 685220 142950 685460
rect 143190 685220 143280 685460
rect 143520 685220 143610 685460
rect 143850 685220 143940 685460
rect 144180 685220 144290 685460
rect 144530 685220 144950 685460
rect 145190 685220 145280 685460
rect 145520 685220 145610 685460
rect 145850 685220 145940 685460
rect 146180 685220 146290 685460
rect 146530 685220 146620 685460
rect 146860 685220 146950 685460
rect 147190 685220 147280 685460
rect 147520 685220 147630 685460
rect 147870 685220 147960 685460
rect 148200 685220 148290 685460
rect 148530 685220 148620 685460
rect 148860 685220 148970 685460
rect 149210 685220 149300 685460
rect 149540 685220 149630 685460
rect 149870 685220 149960 685460
rect 150200 685220 150310 685460
rect 150550 685220 150640 685460
rect 150880 685220 150970 685460
rect 151210 685220 151300 685460
rect 151540 685220 151650 685460
rect 151890 685220 151980 685460
rect 152220 685220 152310 685460
rect 152550 685220 152640 685460
rect 152880 685220 152990 685460
rect 153230 685220 153320 685460
rect 153560 685220 153650 685460
rect 153890 685220 153980 685460
rect 154220 685220 154330 685460
rect 154570 685220 154660 685460
rect 154900 685220 154990 685460
rect 155230 685220 155320 685460
rect 155560 685220 155670 685460
rect 155910 685220 155960 685460
rect 110760 685110 155960 685220
rect 110760 684870 110810 685110
rect 111050 684870 111140 685110
rect 111380 684870 111470 685110
rect 111710 684870 111800 685110
rect 112040 684870 112150 685110
rect 112390 684870 112480 685110
rect 112720 684870 112810 685110
rect 113050 684870 113140 685110
rect 113380 684870 113490 685110
rect 113730 684870 113820 685110
rect 114060 684870 114150 685110
rect 114390 684870 114480 685110
rect 114720 684870 114830 685110
rect 115070 684870 115160 685110
rect 115400 684870 115490 685110
rect 115730 684870 115820 685110
rect 116060 684870 116170 685110
rect 116410 684870 116500 685110
rect 116740 684870 116830 685110
rect 117070 684870 117160 685110
rect 117400 684870 117510 685110
rect 117750 684870 117840 685110
rect 118080 684870 118170 685110
rect 118410 684870 118500 685110
rect 118740 684870 118850 685110
rect 119090 684870 119180 685110
rect 119420 684870 119510 685110
rect 119750 684870 119840 685110
rect 120080 684870 120190 685110
rect 120430 684870 120520 685110
rect 120760 684870 120850 685110
rect 121090 684870 121180 685110
rect 121420 684870 121530 685110
rect 121770 684870 122190 685110
rect 122430 684870 122520 685110
rect 122760 684870 122850 685110
rect 123090 684870 123180 685110
rect 123420 684870 123530 685110
rect 123770 684870 123860 685110
rect 124100 684870 124190 685110
rect 124430 684870 124520 685110
rect 124760 684870 124870 685110
rect 125110 684870 125200 685110
rect 125440 684870 125530 685110
rect 125770 684870 125860 685110
rect 126100 684870 126210 685110
rect 126450 684870 126540 685110
rect 126780 684870 126870 685110
rect 127110 684870 127200 685110
rect 127440 684870 127550 685110
rect 127790 684870 127880 685110
rect 128120 684870 128210 685110
rect 128450 684870 128540 685110
rect 128780 684870 128890 685110
rect 129130 684870 129220 685110
rect 129460 684870 129550 685110
rect 129790 684870 129880 685110
rect 130120 684870 130230 685110
rect 130470 684870 130560 685110
rect 130800 684870 130890 685110
rect 131130 684870 131220 685110
rect 131460 684870 131570 685110
rect 131810 684870 131900 685110
rect 132140 684870 132230 685110
rect 132470 684870 132560 685110
rect 132800 684870 132910 685110
rect 133150 684870 133570 685110
rect 133810 684870 133900 685110
rect 134140 684870 134230 685110
rect 134470 684870 134560 685110
rect 134800 684870 134910 685110
rect 135150 684870 135240 685110
rect 135480 684870 135570 685110
rect 135810 684870 135900 685110
rect 136140 684870 136250 685110
rect 136490 684870 136580 685110
rect 136820 684870 136910 685110
rect 137150 684870 137240 685110
rect 137480 684870 137590 685110
rect 137830 684870 137920 685110
rect 138160 684870 138250 685110
rect 138490 684870 138580 685110
rect 138820 684870 138930 685110
rect 139170 684870 139260 685110
rect 139500 684870 139590 685110
rect 139830 684870 139920 685110
rect 140160 684870 140270 685110
rect 140510 684870 140600 685110
rect 140840 684870 140930 685110
rect 141170 684870 141260 685110
rect 141500 684870 141610 685110
rect 141850 684870 141940 685110
rect 142180 684870 142270 685110
rect 142510 684870 142600 685110
rect 142840 684870 142950 685110
rect 143190 684870 143280 685110
rect 143520 684870 143610 685110
rect 143850 684870 143940 685110
rect 144180 684870 144290 685110
rect 144530 684870 144950 685110
rect 145190 684870 145280 685110
rect 145520 684870 145610 685110
rect 145850 684870 145940 685110
rect 146180 684870 146290 685110
rect 146530 684870 146620 685110
rect 146860 684870 146950 685110
rect 147190 684870 147280 685110
rect 147520 684870 147630 685110
rect 147870 684870 147960 685110
rect 148200 684870 148290 685110
rect 148530 684870 148620 685110
rect 148860 684870 148970 685110
rect 149210 684870 149300 685110
rect 149540 684870 149630 685110
rect 149870 684870 149960 685110
rect 150200 684870 150310 685110
rect 150550 684870 150640 685110
rect 150880 684870 150970 685110
rect 151210 684870 151300 685110
rect 151540 684870 151650 685110
rect 151890 684870 151980 685110
rect 152220 684870 152310 685110
rect 152550 684870 152640 685110
rect 152880 684870 152990 685110
rect 153230 684870 153320 685110
rect 153560 684870 153650 685110
rect 153890 684870 153980 685110
rect 154220 684870 154330 685110
rect 154570 684870 154660 685110
rect 154900 684870 154990 685110
rect 155230 684870 155320 685110
rect 155560 684870 155670 685110
rect 155910 684870 155960 685110
rect 110760 684780 155960 684870
rect 110760 684540 110810 684780
rect 111050 684540 111140 684780
rect 111380 684540 111470 684780
rect 111710 684540 111800 684780
rect 112040 684540 112150 684780
rect 112390 684540 112480 684780
rect 112720 684540 112810 684780
rect 113050 684540 113140 684780
rect 113380 684540 113490 684780
rect 113730 684540 113820 684780
rect 114060 684540 114150 684780
rect 114390 684540 114480 684780
rect 114720 684540 114830 684780
rect 115070 684540 115160 684780
rect 115400 684540 115490 684780
rect 115730 684540 115820 684780
rect 116060 684540 116170 684780
rect 116410 684540 116500 684780
rect 116740 684540 116830 684780
rect 117070 684540 117160 684780
rect 117400 684540 117510 684780
rect 117750 684540 117840 684780
rect 118080 684540 118170 684780
rect 118410 684540 118500 684780
rect 118740 684540 118850 684780
rect 119090 684540 119180 684780
rect 119420 684540 119510 684780
rect 119750 684540 119840 684780
rect 120080 684540 120190 684780
rect 120430 684540 120520 684780
rect 120760 684540 120850 684780
rect 121090 684540 121180 684780
rect 121420 684540 121530 684780
rect 121770 684540 122190 684780
rect 122430 684540 122520 684780
rect 122760 684540 122850 684780
rect 123090 684540 123180 684780
rect 123420 684540 123530 684780
rect 123770 684540 123860 684780
rect 124100 684540 124190 684780
rect 124430 684540 124520 684780
rect 124760 684540 124870 684780
rect 125110 684540 125200 684780
rect 125440 684540 125530 684780
rect 125770 684540 125860 684780
rect 126100 684540 126210 684780
rect 126450 684540 126540 684780
rect 126780 684540 126870 684780
rect 127110 684540 127200 684780
rect 127440 684540 127550 684780
rect 127790 684540 127880 684780
rect 128120 684540 128210 684780
rect 128450 684540 128540 684780
rect 128780 684540 128890 684780
rect 129130 684540 129220 684780
rect 129460 684540 129550 684780
rect 129790 684540 129880 684780
rect 130120 684540 130230 684780
rect 130470 684540 130560 684780
rect 130800 684540 130890 684780
rect 131130 684540 131220 684780
rect 131460 684540 131570 684780
rect 131810 684540 131900 684780
rect 132140 684540 132230 684780
rect 132470 684540 132560 684780
rect 132800 684540 132910 684780
rect 133150 684540 133570 684780
rect 133810 684540 133900 684780
rect 134140 684540 134230 684780
rect 134470 684540 134560 684780
rect 134800 684540 134910 684780
rect 135150 684540 135240 684780
rect 135480 684540 135570 684780
rect 135810 684540 135900 684780
rect 136140 684540 136250 684780
rect 136490 684540 136580 684780
rect 136820 684540 136910 684780
rect 137150 684540 137240 684780
rect 137480 684540 137590 684780
rect 137830 684540 137920 684780
rect 138160 684540 138250 684780
rect 138490 684540 138580 684780
rect 138820 684540 138930 684780
rect 139170 684540 139260 684780
rect 139500 684540 139590 684780
rect 139830 684540 139920 684780
rect 140160 684540 140270 684780
rect 140510 684540 140600 684780
rect 140840 684540 140930 684780
rect 141170 684540 141260 684780
rect 141500 684540 141610 684780
rect 141850 684540 141940 684780
rect 142180 684540 142270 684780
rect 142510 684540 142600 684780
rect 142840 684540 142950 684780
rect 143190 684540 143280 684780
rect 143520 684540 143610 684780
rect 143850 684540 143940 684780
rect 144180 684540 144290 684780
rect 144530 684540 144950 684780
rect 145190 684540 145280 684780
rect 145520 684540 145610 684780
rect 145850 684540 145940 684780
rect 146180 684540 146290 684780
rect 146530 684540 146620 684780
rect 146860 684540 146950 684780
rect 147190 684540 147280 684780
rect 147520 684540 147630 684780
rect 147870 684540 147960 684780
rect 148200 684540 148290 684780
rect 148530 684540 148620 684780
rect 148860 684540 148970 684780
rect 149210 684540 149300 684780
rect 149540 684540 149630 684780
rect 149870 684540 149960 684780
rect 150200 684540 150310 684780
rect 150550 684540 150640 684780
rect 150880 684540 150970 684780
rect 151210 684540 151300 684780
rect 151540 684540 151650 684780
rect 151890 684540 151980 684780
rect 152220 684540 152310 684780
rect 152550 684540 152640 684780
rect 152880 684540 152990 684780
rect 153230 684540 153320 684780
rect 153560 684540 153650 684780
rect 153890 684540 153980 684780
rect 154220 684540 154330 684780
rect 154570 684540 154660 684780
rect 154900 684540 154990 684780
rect 155230 684540 155320 684780
rect 155560 684540 155670 684780
rect 155910 684540 155960 684780
rect 110760 684450 155960 684540
rect 110760 684210 110810 684450
rect 111050 684210 111140 684450
rect 111380 684210 111470 684450
rect 111710 684210 111800 684450
rect 112040 684210 112150 684450
rect 112390 684210 112480 684450
rect 112720 684210 112810 684450
rect 113050 684210 113140 684450
rect 113380 684210 113490 684450
rect 113730 684210 113820 684450
rect 114060 684210 114150 684450
rect 114390 684210 114480 684450
rect 114720 684210 114830 684450
rect 115070 684210 115160 684450
rect 115400 684210 115490 684450
rect 115730 684210 115820 684450
rect 116060 684210 116170 684450
rect 116410 684210 116500 684450
rect 116740 684210 116830 684450
rect 117070 684210 117160 684450
rect 117400 684210 117510 684450
rect 117750 684210 117840 684450
rect 118080 684210 118170 684450
rect 118410 684210 118500 684450
rect 118740 684210 118850 684450
rect 119090 684210 119180 684450
rect 119420 684210 119510 684450
rect 119750 684210 119840 684450
rect 120080 684210 120190 684450
rect 120430 684210 120520 684450
rect 120760 684210 120850 684450
rect 121090 684210 121180 684450
rect 121420 684210 121530 684450
rect 121770 684210 122190 684450
rect 122430 684210 122520 684450
rect 122760 684210 122850 684450
rect 123090 684210 123180 684450
rect 123420 684210 123530 684450
rect 123770 684210 123860 684450
rect 124100 684210 124190 684450
rect 124430 684210 124520 684450
rect 124760 684210 124870 684450
rect 125110 684210 125200 684450
rect 125440 684210 125530 684450
rect 125770 684210 125860 684450
rect 126100 684210 126210 684450
rect 126450 684210 126540 684450
rect 126780 684210 126870 684450
rect 127110 684210 127200 684450
rect 127440 684210 127550 684450
rect 127790 684210 127880 684450
rect 128120 684210 128210 684450
rect 128450 684210 128540 684450
rect 128780 684210 128890 684450
rect 129130 684210 129220 684450
rect 129460 684210 129550 684450
rect 129790 684210 129880 684450
rect 130120 684210 130230 684450
rect 130470 684210 130560 684450
rect 130800 684210 130890 684450
rect 131130 684210 131220 684450
rect 131460 684210 131570 684450
rect 131810 684210 131900 684450
rect 132140 684210 132230 684450
rect 132470 684210 132560 684450
rect 132800 684210 132910 684450
rect 133150 684210 133570 684450
rect 133810 684210 133900 684450
rect 134140 684210 134230 684450
rect 134470 684210 134560 684450
rect 134800 684210 134910 684450
rect 135150 684210 135240 684450
rect 135480 684210 135570 684450
rect 135810 684210 135900 684450
rect 136140 684210 136250 684450
rect 136490 684210 136580 684450
rect 136820 684210 136910 684450
rect 137150 684210 137240 684450
rect 137480 684210 137590 684450
rect 137830 684210 137920 684450
rect 138160 684210 138250 684450
rect 138490 684210 138580 684450
rect 138820 684210 138930 684450
rect 139170 684210 139260 684450
rect 139500 684210 139590 684450
rect 139830 684210 139920 684450
rect 140160 684210 140270 684450
rect 140510 684210 140600 684450
rect 140840 684210 140930 684450
rect 141170 684210 141260 684450
rect 141500 684210 141610 684450
rect 141850 684210 141940 684450
rect 142180 684210 142270 684450
rect 142510 684210 142600 684450
rect 142840 684210 142950 684450
rect 143190 684210 143280 684450
rect 143520 684210 143610 684450
rect 143850 684210 143940 684450
rect 144180 684210 144290 684450
rect 144530 684210 144950 684450
rect 145190 684210 145280 684450
rect 145520 684210 145610 684450
rect 145850 684210 145940 684450
rect 146180 684210 146290 684450
rect 146530 684210 146620 684450
rect 146860 684210 146950 684450
rect 147190 684210 147280 684450
rect 147520 684210 147630 684450
rect 147870 684210 147960 684450
rect 148200 684210 148290 684450
rect 148530 684210 148620 684450
rect 148860 684210 148970 684450
rect 149210 684210 149300 684450
rect 149540 684210 149630 684450
rect 149870 684210 149960 684450
rect 150200 684210 150310 684450
rect 150550 684210 150640 684450
rect 150880 684210 150970 684450
rect 151210 684210 151300 684450
rect 151540 684210 151650 684450
rect 151890 684210 151980 684450
rect 152220 684210 152310 684450
rect 152550 684210 152640 684450
rect 152880 684210 152990 684450
rect 153230 684210 153320 684450
rect 153560 684210 153650 684450
rect 153890 684210 153980 684450
rect 154220 684210 154330 684450
rect 154570 684210 154660 684450
rect 154900 684210 154990 684450
rect 155230 684210 155320 684450
rect 155560 684210 155670 684450
rect 155910 684210 155960 684450
rect 110760 684120 155960 684210
rect 110760 683880 110810 684120
rect 111050 683880 111140 684120
rect 111380 683880 111470 684120
rect 111710 683880 111800 684120
rect 112040 683880 112150 684120
rect 112390 683880 112480 684120
rect 112720 683880 112810 684120
rect 113050 683880 113140 684120
rect 113380 683880 113490 684120
rect 113730 683880 113820 684120
rect 114060 683880 114150 684120
rect 114390 683880 114480 684120
rect 114720 683880 114830 684120
rect 115070 683880 115160 684120
rect 115400 683880 115490 684120
rect 115730 683880 115820 684120
rect 116060 683880 116170 684120
rect 116410 683880 116500 684120
rect 116740 683880 116830 684120
rect 117070 683880 117160 684120
rect 117400 683880 117510 684120
rect 117750 683880 117840 684120
rect 118080 683880 118170 684120
rect 118410 683880 118500 684120
rect 118740 683880 118850 684120
rect 119090 683880 119180 684120
rect 119420 683880 119510 684120
rect 119750 683880 119840 684120
rect 120080 683880 120190 684120
rect 120430 683880 120520 684120
rect 120760 683880 120850 684120
rect 121090 683880 121180 684120
rect 121420 683880 121530 684120
rect 121770 683880 122190 684120
rect 122430 683880 122520 684120
rect 122760 683880 122850 684120
rect 123090 683880 123180 684120
rect 123420 683880 123530 684120
rect 123770 683880 123860 684120
rect 124100 683880 124190 684120
rect 124430 683880 124520 684120
rect 124760 683880 124870 684120
rect 125110 683880 125200 684120
rect 125440 683880 125530 684120
rect 125770 683880 125860 684120
rect 126100 683880 126210 684120
rect 126450 683880 126540 684120
rect 126780 683880 126870 684120
rect 127110 683880 127200 684120
rect 127440 683880 127550 684120
rect 127790 683880 127880 684120
rect 128120 683880 128210 684120
rect 128450 683880 128540 684120
rect 128780 683880 128890 684120
rect 129130 683880 129220 684120
rect 129460 683880 129550 684120
rect 129790 683880 129880 684120
rect 130120 683880 130230 684120
rect 130470 683880 130560 684120
rect 130800 683880 130890 684120
rect 131130 683880 131220 684120
rect 131460 683880 131570 684120
rect 131810 683880 131900 684120
rect 132140 683880 132230 684120
rect 132470 683880 132560 684120
rect 132800 683880 132910 684120
rect 133150 683880 133570 684120
rect 133810 683880 133900 684120
rect 134140 683880 134230 684120
rect 134470 683880 134560 684120
rect 134800 683880 134910 684120
rect 135150 683880 135240 684120
rect 135480 683880 135570 684120
rect 135810 683880 135900 684120
rect 136140 683880 136250 684120
rect 136490 683880 136580 684120
rect 136820 683880 136910 684120
rect 137150 683880 137240 684120
rect 137480 683880 137590 684120
rect 137830 683880 137920 684120
rect 138160 683880 138250 684120
rect 138490 683880 138580 684120
rect 138820 683880 138930 684120
rect 139170 683880 139260 684120
rect 139500 683880 139590 684120
rect 139830 683880 139920 684120
rect 140160 683880 140270 684120
rect 140510 683880 140600 684120
rect 140840 683880 140930 684120
rect 141170 683880 141260 684120
rect 141500 683880 141610 684120
rect 141850 683880 141940 684120
rect 142180 683880 142270 684120
rect 142510 683880 142600 684120
rect 142840 683880 142950 684120
rect 143190 683880 143280 684120
rect 143520 683880 143610 684120
rect 143850 683880 143940 684120
rect 144180 683880 144290 684120
rect 144530 683880 144950 684120
rect 145190 683880 145280 684120
rect 145520 683880 145610 684120
rect 145850 683880 145940 684120
rect 146180 683880 146290 684120
rect 146530 683880 146620 684120
rect 146860 683880 146950 684120
rect 147190 683880 147280 684120
rect 147520 683880 147630 684120
rect 147870 683880 147960 684120
rect 148200 683880 148290 684120
rect 148530 683880 148620 684120
rect 148860 683880 148970 684120
rect 149210 683880 149300 684120
rect 149540 683880 149630 684120
rect 149870 683880 149960 684120
rect 150200 683880 150310 684120
rect 150550 683880 150640 684120
rect 150880 683880 150970 684120
rect 151210 683880 151300 684120
rect 151540 683880 151650 684120
rect 151890 683880 151980 684120
rect 152220 683880 152310 684120
rect 152550 683880 152640 684120
rect 152880 683880 152990 684120
rect 153230 683880 153320 684120
rect 153560 683880 153650 684120
rect 153890 683880 153980 684120
rect 154220 683880 154330 684120
rect 154570 683880 154660 684120
rect 154900 683880 154990 684120
rect 155230 683880 155320 684120
rect 155560 683880 155670 684120
rect 155910 683880 155960 684120
rect 110760 683700 155960 683880
rect 110760 683460 110890 683700
rect 111130 683460 111220 683700
rect 111460 683460 111550 683700
rect 111790 683460 111880 683700
rect 112120 683460 112210 683700
rect 112450 683460 112540 683700
rect 112780 683460 112870 683700
rect 113110 683460 113200 683700
rect 113440 683460 113530 683700
rect 113770 683460 113860 683700
rect 114100 683460 114190 683700
rect 114430 683460 114520 683700
rect 114760 683460 114850 683700
rect 115090 683460 115180 683700
rect 115420 683460 115510 683700
rect 115750 683460 115840 683700
rect 116080 683460 116170 683700
rect 116410 683460 116500 683700
rect 116740 683460 116830 683700
rect 117070 683460 117160 683700
rect 117400 683460 117490 683700
rect 117730 683460 117820 683700
rect 118060 683460 118150 683700
rect 118390 683460 118480 683700
rect 118720 683460 118810 683700
rect 119050 683460 119140 683700
rect 119380 683460 119470 683700
rect 119710 683460 119800 683700
rect 120040 683460 120130 683700
rect 120370 683460 120460 683700
rect 120700 683460 120790 683700
rect 121030 683460 121120 683700
rect 121360 683460 121450 683700
rect 121690 683460 122270 683700
rect 122510 683460 122600 683700
rect 122840 683460 122930 683700
rect 123170 683460 123260 683700
rect 123500 683460 123590 683700
rect 123830 683460 123920 683700
rect 124160 683460 124250 683700
rect 124490 683460 124580 683700
rect 124820 683460 124910 683700
rect 125150 683460 125240 683700
rect 125480 683460 125570 683700
rect 125810 683460 125900 683700
rect 126140 683460 126230 683700
rect 126470 683460 126560 683700
rect 126800 683460 126890 683700
rect 127130 683460 127220 683700
rect 127460 683460 127550 683700
rect 127790 683460 127880 683700
rect 128120 683460 128210 683700
rect 128450 683460 128540 683700
rect 128780 683460 128870 683700
rect 129110 683460 129200 683700
rect 129440 683460 129530 683700
rect 129770 683460 129860 683700
rect 130100 683460 130190 683700
rect 130430 683460 130520 683700
rect 130760 683460 130850 683700
rect 131090 683460 131180 683700
rect 131420 683460 131510 683700
rect 131750 683460 131840 683700
rect 132080 683460 132170 683700
rect 132410 683460 132500 683700
rect 132740 683460 132830 683700
rect 133070 683460 133650 683700
rect 133890 683460 133980 683700
rect 134220 683460 134310 683700
rect 134550 683460 134640 683700
rect 134880 683460 134970 683700
rect 135210 683460 135300 683700
rect 135540 683460 135630 683700
rect 135870 683460 135960 683700
rect 136200 683460 136290 683700
rect 136530 683460 136620 683700
rect 136860 683460 136950 683700
rect 137190 683460 137280 683700
rect 137520 683460 137610 683700
rect 137850 683460 137940 683700
rect 138180 683460 138270 683700
rect 138510 683460 138600 683700
rect 138840 683460 138930 683700
rect 139170 683460 139260 683700
rect 139500 683460 139590 683700
rect 139830 683460 139920 683700
rect 140160 683460 140250 683700
rect 140490 683460 140580 683700
rect 140820 683460 140910 683700
rect 141150 683460 141240 683700
rect 141480 683460 141570 683700
rect 141810 683460 141900 683700
rect 142140 683460 142230 683700
rect 142470 683460 142560 683700
rect 142800 683460 142890 683700
rect 143130 683460 143220 683700
rect 143460 683460 143550 683700
rect 143790 683460 143880 683700
rect 144120 683460 144210 683700
rect 144450 683460 145030 683700
rect 145270 683460 145360 683700
rect 145600 683460 145690 683700
rect 145930 683460 146020 683700
rect 146260 683460 146350 683700
rect 146590 683460 146680 683700
rect 146920 683460 147010 683700
rect 147250 683460 147340 683700
rect 147580 683460 147670 683700
rect 147910 683460 148000 683700
rect 148240 683460 148330 683700
rect 148570 683460 148660 683700
rect 148900 683460 148990 683700
rect 149230 683460 149320 683700
rect 149560 683460 149650 683700
rect 149890 683460 149980 683700
rect 150220 683460 150310 683700
rect 150550 683460 150640 683700
rect 150880 683460 150970 683700
rect 151210 683460 151300 683700
rect 151540 683460 151630 683700
rect 151870 683460 151960 683700
rect 152200 683460 152290 683700
rect 152530 683460 152620 683700
rect 152860 683460 152950 683700
rect 153190 683460 153280 683700
rect 153520 683460 153610 683700
rect 153850 683460 153940 683700
rect 154180 683460 154270 683700
rect 154510 683460 154600 683700
rect 154840 683460 154930 683700
rect 155170 683460 155260 683700
rect 155500 683460 155590 683700
rect 155830 683460 155960 683700
rect 110760 683280 155960 683460
rect 110760 683040 110810 683280
rect 111050 683040 111160 683280
rect 111400 683040 111490 683280
rect 111730 683040 111820 683280
rect 112060 683040 112150 683280
rect 112390 683040 112500 683280
rect 112740 683040 112830 683280
rect 113070 683040 113160 683280
rect 113400 683040 113490 683280
rect 113730 683040 113840 683280
rect 114080 683040 114170 683280
rect 114410 683040 114500 683280
rect 114740 683040 114830 683280
rect 115070 683040 115180 683280
rect 115420 683040 115510 683280
rect 115750 683040 115840 683280
rect 116080 683040 116170 683280
rect 116410 683040 116520 683280
rect 116760 683040 116850 683280
rect 117090 683040 117180 683280
rect 117420 683040 117510 683280
rect 117750 683040 117860 683280
rect 118100 683040 118190 683280
rect 118430 683040 118520 683280
rect 118760 683040 118850 683280
rect 119090 683040 119200 683280
rect 119440 683040 119530 683280
rect 119770 683040 119860 683280
rect 120100 683040 120190 683280
rect 120430 683040 120540 683280
rect 120780 683040 120870 683280
rect 121110 683040 121200 683280
rect 121440 683040 121530 683280
rect 121770 683040 122190 683280
rect 122430 683040 122540 683280
rect 122780 683040 122870 683280
rect 123110 683040 123200 683280
rect 123440 683040 123530 683280
rect 123770 683040 123880 683280
rect 124120 683040 124210 683280
rect 124450 683040 124540 683280
rect 124780 683040 124870 683280
rect 125110 683040 125220 683280
rect 125460 683040 125550 683280
rect 125790 683040 125880 683280
rect 126120 683040 126210 683280
rect 126450 683040 126560 683280
rect 126800 683040 126890 683280
rect 127130 683040 127220 683280
rect 127460 683040 127550 683280
rect 127790 683040 127900 683280
rect 128140 683040 128230 683280
rect 128470 683040 128560 683280
rect 128800 683040 128890 683280
rect 129130 683040 129240 683280
rect 129480 683040 129570 683280
rect 129810 683040 129900 683280
rect 130140 683040 130230 683280
rect 130470 683040 130580 683280
rect 130820 683040 130910 683280
rect 131150 683040 131240 683280
rect 131480 683040 131570 683280
rect 131810 683040 131920 683280
rect 132160 683040 132250 683280
rect 132490 683040 132580 683280
rect 132820 683040 132910 683280
rect 133150 683040 133570 683280
rect 133810 683040 133920 683280
rect 134160 683040 134250 683280
rect 134490 683040 134580 683280
rect 134820 683040 134910 683280
rect 135150 683040 135260 683280
rect 135500 683040 135590 683280
rect 135830 683040 135920 683280
rect 136160 683040 136250 683280
rect 136490 683040 136600 683280
rect 136840 683040 136930 683280
rect 137170 683040 137260 683280
rect 137500 683040 137590 683280
rect 137830 683040 137940 683280
rect 138180 683040 138270 683280
rect 138510 683040 138600 683280
rect 138840 683040 138930 683280
rect 139170 683040 139280 683280
rect 139520 683040 139610 683280
rect 139850 683040 139940 683280
rect 140180 683040 140270 683280
rect 140510 683040 140620 683280
rect 140860 683040 140950 683280
rect 141190 683040 141280 683280
rect 141520 683040 141610 683280
rect 141850 683040 141960 683280
rect 142200 683040 142290 683280
rect 142530 683040 142620 683280
rect 142860 683040 142950 683280
rect 143190 683040 143300 683280
rect 143540 683040 143630 683280
rect 143870 683040 143960 683280
rect 144200 683040 144290 683280
rect 144530 683040 144950 683280
rect 145190 683040 145300 683280
rect 145540 683040 145630 683280
rect 145870 683040 145960 683280
rect 146200 683040 146290 683280
rect 146530 683040 146640 683280
rect 146880 683040 146970 683280
rect 147210 683040 147300 683280
rect 147540 683040 147630 683280
rect 147870 683040 147980 683280
rect 148220 683040 148310 683280
rect 148550 683040 148640 683280
rect 148880 683040 148970 683280
rect 149210 683040 149320 683280
rect 149560 683040 149650 683280
rect 149890 683040 149980 683280
rect 150220 683040 150310 683280
rect 150550 683040 150660 683280
rect 150900 683040 150990 683280
rect 151230 683040 151320 683280
rect 151560 683040 151650 683280
rect 151890 683040 152000 683280
rect 152240 683040 152330 683280
rect 152570 683040 152660 683280
rect 152900 683040 152990 683280
rect 153230 683040 153340 683280
rect 153580 683040 153670 683280
rect 153910 683040 154000 683280
rect 154240 683040 154330 683280
rect 154570 683040 154680 683280
rect 154920 683040 155010 683280
rect 155250 683040 155340 683280
rect 155580 683040 155670 683280
rect 155910 683040 155960 683280
rect 110760 682950 155960 683040
rect 110760 682710 110810 682950
rect 111050 682710 111160 682950
rect 111400 682710 111490 682950
rect 111730 682710 111820 682950
rect 112060 682710 112150 682950
rect 112390 682710 112500 682950
rect 112740 682710 112830 682950
rect 113070 682710 113160 682950
rect 113400 682710 113490 682950
rect 113730 682710 113840 682950
rect 114080 682710 114170 682950
rect 114410 682710 114500 682950
rect 114740 682710 114830 682950
rect 115070 682710 115180 682950
rect 115420 682710 115510 682950
rect 115750 682710 115840 682950
rect 116080 682710 116170 682950
rect 116410 682710 116520 682950
rect 116760 682710 116850 682950
rect 117090 682710 117180 682950
rect 117420 682710 117510 682950
rect 117750 682710 117860 682950
rect 118100 682710 118190 682950
rect 118430 682710 118520 682950
rect 118760 682710 118850 682950
rect 119090 682710 119200 682950
rect 119440 682710 119530 682950
rect 119770 682710 119860 682950
rect 120100 682710 120190 682950
rect 120430 682710 120540 682950
rect 120780 682710 120870 682950
rect 121110 682710 121200 682950
rect 121440 682710 121530 682950
rect 121770 682710 122190 682950
rect 122430 682710 122540 682950
rect 122780 682710 122870 682950
rect 123110 682710 123200 682950
rect 123440 682710 123530 682950
rect 123770 682710 123880 682950
rect 124120 682710 124210 682950
rect 124450 682710 124540 682950
rect 124780 682710 124870 682950
rect 125110 682710 125220 682950
rect 125460 682710 125550 682950
rect 125790 682710 125880 682950
rect 126120 682710 126210 682950
rect 126450 682710 126560 682950
rect 126800 682710 126890 682950
rect 127130 682710 127220 682950
rect 127460 682710 127550 682950
rect 127790 682710 127900 682950
rect 128140 682710 128230 682950
rect 128470 682710 128560 682950
rect 128800 682710 128890 682950
rect 129130 682710 129240 682950
rect 129480 682710 129570 682950
rect 129810 682710 129900 682950
rect 130140 682710 130230 682950
rect 130470 682710 130580 682950
rect 130820 682710 130910 682950
rect 131150 682710 131240 682950
rect 131480 682710 131570 682950
rect 131810 682710 131920 682950
rect 132160 682710 132250 682950
rect 132490 682710 132580 682950
rect 132820 682710 132910 682950
rect 133150 682710 133570 682950
rect 133810 682710 133920 682950
rect 134160 682710 134250 682950
rect 134490 682710 134580 682950
rect 134820 682710 134910 682950
rect 135150 682710 135260 682950
rect 135500 682710 135590 682950
rect 135830 682710 135920 682950
rect 136160 682710 136250 682950
rect 136490 682710 136600 682950
rect 136840 682710 136930 682950
rect 137170 682710 137260 682950
rect 137500 682710 137590 682950
rect 137830 682710 137940 682950
rect 138180 682710 138270 682950
rect 138510 682710 138600 682950
rect 138840 682710 138930 682950
rect 139170 682710 139280 682950
rect 139520 682710 139610 682950
rect 139850 682710 139940 682950
rect 140180 682710 140270 682950
rect 140510 682710 140620 682950
rect 140860 682710 140950 682950
rect 141190 682710 141280 682950
rect 141520 682710 141610 682950
rect 141850 682710 141960 682950
rect 142200 682710 142290 682950
rect 142530 682710 142620 682950
rect 142860 682710 142950 682950
rect 143190 682710 143300 682950
rect 143540 682710 143630 682950
rect 143870 682710 143960 682950
rect 144200 682710 144290 682950
rect 144530 682710 144950 682950
rect 145190 682710 145300 682950
rect 145540 682710 145630 682950
rect 145870 682710 145960 682950
rect 146200 682710 146290 682950
rect 146530 682710 146640 682950
rect 146880 682710 146970 682950
rect 147210 682710 147300 682950
rect 147540 682710 147630 682950
rect 147870 682710 147980 682950
rect 148220 682710 148310 682950
rect 148550 682710 148640 682950
rect 148880 682710 148970 682950
rect 149210 682710 149320 682950
rect 149560 682710 149650 682950
rect 149890 682710 149980 682950
rect 150220 682710 150310 682950
rect 150550 682710 150660 682950
rect 150900 682710 150990 682950
rect 151230 682710 151320 682950
rect 151560 682710 151650 682950
rect 151890 682710 152000 682950
rect 152240 682710 152330 682950
rect 152570 682710 152660 682950
rect 152900 682710 152990 682950
rect 153230 682710 153340 682950
rect 153580 682710 153670 682950
rect 153910 682710 154000 682950
rect 154240 682710 154330 682950
rect 154570 682710 154680 682950
rect 154920 682710 155010 682950
rect 155250 682710 155340 682950
rect 155580 682710 155670 682950
rect 155910 682710 155960 682950
rect 110760 682620 155960 682710
rect 110760 682380 110810 682620
rect 111050 682380 111160 682620
rect 111400 682380 111490 682620
rect 111730 682380 111820 682620
rect 112060 682380 112150 682620
rect 112390 682380 112500 682620
rect 112740 682380 112830 682620
rect 113070 682380 113160 682620
rect 113400 682380 113490 682620
rect 113730 682380 113840 682620
rect 114080 682380 114170 682620
rect 114410 682380 114500 682620
rect 114740 682380 114830 682620
rect 115070 682380 115180 682620
rect 115420 682380 115510 682620
rect 115750 682380 115840 682620
rect 116080 682380 116170 682620
rect 116410 682380 116520 682620
rect 116760 682380 116850 682620
rect 117090 682380 117180 682620
rect 117420 682380 117510 682620
rect 117750 682380 117860 682620
rect 118100 682380 118190 682620
rect 118430 682380 118520 682620
rect 118760 682380 118850 682620
rect 119090 682380 119200 682620
rect 119440 682380 119530 682620
rect 119770 682380 119860 682620
rect 120100 682380 120190 682620
rect 120430 682380 120540 682620
rect 120780 682380 120870 682620
rect 121110 682380 121200 682620
rect 121440 682380 121530 682620
rect 121770 682380 122190 682620
rect 122430 682380 122540 682620
rect 122780 682380 122870 682620
rect 123110 682380 123200 682620
rect 123440 682380 123530 682620
rect 123770 682380 123880 682620
rect 124120 682380 124210 682620
rect 124450 682380 124540 682620
rect 124780 682380 124870 682620
rect 125110 682380 125220 682620
rect 125460 682380 125550 682620
rect 125790 682380 125880 682620
rect 126120 682380 126210 682620
rect 126450 682380 126560 682620
rect 126800 682380 126890 682620
rect 127130 682380 127220 682620
rect 127460 682380 127550 682620
rect 127790 682380 127900 682620
rect 128140 682380 128230 682620
rect 128470 682380 128560 682620
rect 128800 682380 128890 682620
rect 129130 682380 129240 682620
rect 129480 682380 129570 682620
rect 129810 682380 129900 682620
rect 130140 682380 130230 682620
rect 130470 682380 130580 682620
rect 130820 682380 130910 682620
rect 131150 682380 131240 682620
rect 131480 682380 131570 682620
rect 131810 682380 131920 682620
rect 132160 682380 132250 682620
rect 132490 682380 132580 682620
rect 132820 682380 132910 682620
rect 133150 682380 133570 682620
rect 133810 682380 133920 682620
rect 134160 682380 134250 682620
rect 134490 682380 134580 682620
rect 134820 682380 134910 682620
rect 135150 682380 135260 682620
rect 135500 682380 135590 682620
rect 135830 682380 135920 682620
rect 136160 682380 136250 682620
rect 136490 682380 136600 682620
rect 136840 682380 136930 682620
rect 137170 682380 137260 682620
rect 137500 682380 137590 682620
rect 137830 682380 137940 682620
rect 138180 682380 138270 682620
rect 138510 682380 138600 682620
rect 138840 682380 138930 682620
rect 139170 682380 139280 682620
rect 139520 682380 139610 682620
rect 139850 682380 139940 682620
rect 140180 682380 140270 682620
rect 140510 682380 140620 682620
rect 140860 682380 140950 682620
rect 141190 682380 141280 682620
rect 141520 682380 141610 682620
rect 141850 682380 141960 682620
rect 142200 682380 142290 682620
rect 142530 682380 142620 682620
rect 142860 682380 142950 682620
rect 143190 682380 143300 682620
rect 143540 682380 143630 682620
rect 143870 682380 143960 682620
rect 144200 682380 144290 682620
rect 144530 682380 144950 682620
rect 145190 682380 145300 682620
rect 145540 682380 145630 682620
rect 145870 682380 145960 682620
rect 146200 682380 146290 682620
rect 146530 682380 146640 682620
rect 146880 682380 146970 682620
rect 147210 682380 147300 682620
rect 147540 682380 147630 682620
rect 147870 682380 147980 682620
rect 148220 682380 148310 682620
rect 148550 682380 148640 682620
rect 148880 682380 148970 682620
rect 149210 682380 149320 682620
rect 149560 682380 149650 682620
rect 149890 682380 149980 682620
rect 150220 682380 150310 682620
rect 150550 682380 150660 682620
rect 150900 682380 150990 682620
rect 151230 682380 151320 682620
rect 151560 682380 151650 682620
rect 151890 682380 152000 682620
rect 152240 682380 152330 682620
rect 152570 682380 152660 682620
rect 152900 682380 152990 682620
rect 153230 682380 153340 682620
rect 153580 682380 153670 682620
rect 153910 682380 154000 682620
rect 154240 682380 154330 682620
rect 154570 682380 154680 682620
rect 154920 682380 155010 682620
rect 155250 682380 155340 682620
rect 155580 682380 155670 682620
rect 155910 682380 155960 682620
rect 110760 682290 155960 682380
rect 110760 682050 110810 682290
rect 111050 682050 111160 682290
rect 111400 682050 111490 682290
rect 111730 682050 111820 682290
rect 112060 682050 112150 682290
rect 112390 682050 112500 682290
rect 112740 682050 112830 682290
rect 113070 682050 113160 682290
rect 113400 682050 113490 682290
rect 113730 682050 113840 682290
rect 114080 682050 114170 682290
rect 114410 682050 114500 682290
rect 114740 682050 114830 682290
rect 115070 682050 115180 682290
rect 115420 682050 115510 682290
rect 115750 682050 115840 682290
rect 116080 682050 116170 682290
rect 116410 682050 116520 682290
rect 116760 682050 116850 682290
rect 117090 682050 117180 682290
rect 117420 682050 117510 682290
rect 117750 682050 117860 682290
rect 118100 682050 118190 682290
rect 118430 682050 118520 682290
rect 118760 682050 118850 682290
rect 119090 682050 119200 682290
rect 119440 682050 119530 682290
rect 119770 682050 119860 682290
rect 120100 682050 120190 682290
rect 120430 682050 120540 682290
rect 120780 682050 120870 682290
rect 121110 682050 121200 682290
rect 121440 682050 121530 682290
rect 121770 682050 122190 682290
rect 122430 682050 122540 682290
rect 122780 682050 122870 682290
rect 123110 682050 123200 682290
rect 123440 682050 123530 682290
rect 123770 682050 123880 682290
rect 124120 682050 124210 682290
rect 124450 682050 124540 682290
rect 124780 682050 124870 682290
rect 125110 682050 125220 682290
rect 125460 682050 125550 682290
rect 125790 682050 125880 682290
rect 126120 682050 126210 682290
rect 126450 682050 126560 682290
rect 126800 682050 126890 682290
rect 127130 682050 127220 682290
rect 127460 682050 127550 682290
rect 127790 682050 127900 682290
rect 128140 682050 128230 682290
rect 128470 682050 128560 682290
rect 128800 682050 128890 682290
rect 129130 682050 129240 682290
rect 129480 682050 129570 682290
rect 129810 682050 129900 682290
rect 130140 682050 130230 682290
rect 130470 682050 130580 682290
rect 130820 682050 130910 682290
rect 131150 682050 131240 682290
rect 131480 682050 131570 682290
rect 131810 682050 131920 682290
rect 132160 682050 132250 682290
rect 132490 682050 132580 682290
rect 132820 682050 132910 682290
rect 133150 682050 133570 682290
rect 133810 682050 133920 682290
rect 134160 682050 134250 682290
rect 134490 682050 134580 682290
rect 134820 682050 134910 682290
rect 135150 682050 135260 682290
rect 135500 682050 135590 682290
rect 135830 682050 135920 682290
rect 136160 682050 136250 682290
rect 136490 682050 136600 682290
rect 136840 682050 136930 682290
rect 137170 682050 137260 682290
rect 137500 682050 137590 682290
rect 137830 682050 137940 682290
rect 138180 682050 138270 682290
rect 138510 682050 138600 682290
rect 138840 682050 138930 682290
rect 139170 682050 139280 682290
rect 139520 682050 139610 682290
rect 139850 682050 139940 682290
rect 140180 682050 140270 682290
rect 140510 682050 140620 682290
rect 140860 682050 140950 682290
rect 141190 682050 141280 682290
rect 141520 682050 141610 682290
rect 141850 682050 141960 682290
rect 142200 682050 142290 682290
rect 142530 682050 142620 682290
rect 142860 682050 142950 682290
rect 143190 682050 143300 682290
rect 143540 682050 143630 682290
rect 143870 682050 143960 682290
rect 144200 682050 144290 682290
rect 144530 682050 144950 682290
rect 145190 682050 145300 682290
rect 145540 682050 145630 682290
rect 145870 682050 145960 682290
rect 146200 682050 146290 682290
rect 146530 682050 146640 682290
rect 146880 682050 146970 682290
rect 147210 682050 147300 682290
rect 147540 682050 147630 682290
rect 147870 682050 147980 682290
rect 148220 682050 148310 682290
rect 148550 682050 148640 682290
rect 148880 682050 148970 682290
rect 149210 682050 149320 682290
rect 149560 682050 149650 682290
rect 149890 682050 149980 682290
rect 150220 682050 150310 682290
rect 150550 682050 150660 682290
rect 150900 682050 150990 682290
rect 151230 682050 151320 682290
rect 151560 682050 151650 682290
rect 151890 682050 152000 682290
rect 152240 682050 152330 682290
rect 152570 682050 152660 682290
rect 152900 682050 152990 682290
rect 153230 682050 153340 682290
rect 153580 682050 153670 682290
rect 153910 682050 154000 682290
rect 154240 682050 154330 682290
rect 154570 682050 154680 682290
rect 154920 682050 155010 682290
rect 155250 682050 155340 682290
rect 155580 682050 155670 682290
rect 155910 682050 155960 682290
rect 110760 681940 155960 682050
rect 110760 681700 110810 681940
rect 111050 681700 111160 681940
rect 111400 681700 111490 681940
rect 111730 681700 111820 681940
rect 112060 681700 112150 681940
rect 112390 681700 112500 681940
rect 112740 681700 112830 681940
rect 113070 681700 113160 681940
rect 113400 681700 113490 681940
rect 113730 681700 113840 681940
rect 114080 681700 114170 681940
rect 114410 681700 114500 681940
rect 114740 681700 114830 681940
rect 115070 681700 115180 681940
rect 115420 681700 115510 681940
rect 115750 681700 115840 681940
rect 116080 681700 116170 681940
rect 116410 681700 116520 681940
rect 116760 681700 116850 681940
rect 117090 681700 117180 681940
rect 117420 681700 117510 681940
rect 117750 681700 117860 681940
rect 118100 681700 118190 681940
rect 118430 681700 118520 681940
rect 118760 681700 118850 681940
rect 119090 681700 119200 681940
rect 119440 681700 119530 681940
rect 119770 681700 119860 681940
rect 120100 681700 120190 681940
rect 120430 681700 120540 681940
rect 120780 681700 120870 681940
rect 121110 681700 121200 681940
rect 121440 681700 121530 681940
rect 121770 681700 122190 681940
rect 122430 681700 122540 681940
rect 122780 681700 122870 681940
rect 123110 681700 123200 681940
rect 123440 681700 123530 681940
rect 123770 681700 123880 681940
rect 124120 681700 124210 681940
rect 124450 681700 124540 681940
rect 124780 681700 124870 681940
rect 125110 681700 125220 681940
rect 125460 681700 125550 681940
rect 125790 681700 125880 681940
rect 126120 681700 126210 681940
rect 126450 681700 126560 681940
rect 126800 681700 126890 681940
rect 127130 681700 127220 681940
rect 127460 681700 127550 681940
rect 127790 681700 127900 681940
rect 128140 681700 128230 681940
rect 128470 681700 128560 681940
rect 128800 681700 128890 681940
rect 129130 681700 129240 681940
rect 129480 681700 129570 681940
rect 129810 681700 129900 681940
rect 130140 681700 130230 681940
rect 130470 681700 130580 681940
rect 130820 681700 130910 681940
rect 131150 681700 131240 681940
rect 131480 681700 131570 681940
rect 131810 681700 131920 681940
rect 132160 681700 132250 681940
rect 132490 681700 132580 681940
rect 132820 681700 132910 681940
rect 133150 681700 133570 681940
rect 133810 681700 133920 681940
rect 134160 681700 134250 681940
rect 134490 681700 134580 681940
rect 134820 681700 134910 681940
rect 135150 681700 135260 681940
rect 135500 681700 135590 681940
rect 135830 681700 135920 681940
rect 136160 681700 136250 681940
rect 136490 681700 136600 681940
rect 136840 681700 136930 681940
rect 137170 681700 137260 681940
rect 137500 681700 137590 681940
rect 137830 681700 137940 681940
rect 138180 681700 138270 681940
rect 138510 681700 138600 681940
rect 138840 681700 138930 681940
rect 139170 681700 139280 681940
rect 139520 681700 139610 681940
rect 139850 681700 139940 681940
rect 140180 681700 140270 681940
rect 140510 681700 140620 681940
rect 140860 681700 140950 681940
rect 141190 681700 141280 681940
rect 141520 681700 141610 681940
rect 141850 681700 141960 681940
rect 142200 681700 142290 681940
rect 142530 681700 142620 681940
rect 142860 681700 142950 681940
rect 143190 681700 143300 681940
rect 143540 681700 143630 681940
rect 143870 681700 143960 681940
rect 144200 681700 144290 681940
rect 144530 681700 144950 681940
rect 145190 681700 145300 681940
rect 145540 681700 145630 681940
rect 145870 681700 145960 681940
rect 146200 681700 146290 681940
rect 146530 681700 146640 681940
rect 146880 681700 146970 681940
rect 147210 681700 147300 681940
rect 147540 681700 147630 681940
rect 147870 681700 147980 681940
rect 148220 681700 148310 681940
rect 148550 681700 148640 681940
rect 148880 681700 148970 681940
rect 149210 681700 149320 681940
rect 149560 681700 149650 681940
rect 149890 681700 149980 681940
rect 150220 681700 150310 681940
rect 150550 681700 150660 681940
rect 150900 681700 150990 681940
rect 151230 681700 151320 681940
rect 151560 681700 151650 681940
rect 151890 681700 152000 681940
rect 152240 681700 152330 681940
rect 152570 681700 152660 681940
rect 152900 681700 152990 681940
rect 153230 681700 153340 681940
rect 153580 681700 153670 681940
rect 153910 681700 154000 681940
rect 154240 681700 154330 681940
rect 154570 681700 154680 681940
rect 154920 681700 155010 681940
rect 155250 681700 155340 681940
rect 155580 681700 155670 681940
rect 155910 681700 155960 681940
rect 110760 681610 155960 681700
rect 110760 681370 110810 681610
rect 111050 681370 111160 681610
rect 111400 681370 111490 681610
rect 111730 681370 111820 681610
rect 112060 681370 112150 681610
rect 112390 681370 112500 681610
rect 112740 681370 112830 681610
rect 113070 681370 113160 681610
rect 113400 681370 113490 681610
rect 113730 681370 113840 681610
rect 114080 681370 114170 681610
rect 114410 681370 114500 681610
rect 114740 681370 114830 681610
rect 115070 681370 115180 681610
rect 115420 681370 115510 681610
rect 115750 681370 115840 681610
rect 116080 681370 116170 681610
rect 116410 681370 116520 681610
rect 116760 681370 116850 681610
rect 117090 681370 117180 681610
rect 117420 681370 117510 681610
rect 117750 681370 117860 681610
rect 118100 681370 118190 681610
rect 118430 681370 118520 681610
rect 118760 681370 118850 681610
rect 119090 681370 119200 681610
rect 119440 681370 119530 681610
rect 119770 681370 119860 681610
rect 120100 681370 120190 681610
rect 120430 681370 120540 681610
rect 120780 681370 120870 681610
rect 121110 681370 121200 681610
rect 121440 681370 121530 681610
rect 121770 681370 122190 681610
rect 122430 681370 122540 681610
rect 122780 681370 122870 681610
rect 123110 681370 123200 681610
rect 123440 681370 123530 681610
rect 123770 681370 123880 681610
rect 124120 681370 124210 681610
rect 124450 681370 124540 681610
rect 124780 681370 124870 681610
rect 125110 681370 125220 681610
rect 125460 681370 125550 681610
rect 125790 681370 125880 681610
rect 126120 681370 126210 681610
rect 126450 681370 126560 681610
rect 126800 681370 126890 681610
rect 127130 681370 127220 681610
rect 127460 681370 127550 681610
rect 127790 681370 127900 681610
rect 128140 681370 128230 681610
rect 128470 681370 128560 681610
rect 128800 681370 128890 681610
rect 129130 681370 129240 681610
rect 129480 681370 129570 681610
rect 129810 681370 129900 681610
rect 130140 681370 130230 681610
rect 130470 681370 130580 681610
rect 130820 681370 130910 681610
rect 131150 681370 131240 681610
rect 131480 681370 131570 681610
rect 131810 681370 131920 681610
rect 132160 681370 132250 681610
rect 132490 681370 132580 681610
rect 132820 681370 132910 681610
rect 133150 681370 133570 681610
rect 133810 681370 133920 681610
rect 134160 681370 134250 681610
rect 134490 681370 134580 681610
rect 134820 681370 134910 681610
rect 135150 681370 135260 681610
rect 135500 681370 135590 681610
rect 135830 681370 135920 681610
rect 136160 681370 136250 681610
rect 136490 681370 136600 681610
rect 136840 681370 136930 681610
rect 137170 681370 137260 681610
rect 137500 681370 137590 681610
rect 137830 681370 137940 681610
rect 138180 681370 138270 681610
rect 138510 681370 138600 681610
rect 138840 681370 138930 681610
rect 139170 681370 139280 681610
rect 139520 681370 139610 681610
rect 139850 681370 139940 681610
rect 140180 681370 140270 681610
rect 140510 681370 140620 681610
rect 140860 681370 140950 681610
rect 141190 681370 141280 681610
rect 141520 681370 141610 681610
rect 141850 681370 141960 681610
rect 142200 681370 142290 681610
rect 142530 681370 142620 681610
rect 142860 681370 142950 681610
rect 143190 681370 143300 681610
rect 143540 681370 143630 681610
rect 143870 681370 143960 681610
rect 144200 681370 144290 681610
rect 144530 681370 144950 681610
rect 145190 681370 145300 681610
rect 145540 681370 145630 681610
rect 145870 681370 145960 681610
rect 146200 681370 146290 681610
rect 146530 681370 146640 681610
rect 146880 681370 146970 681610
rect 147210 681370 147300 681610
rect 147540 681370 147630 681610
rect 147870 681370 147980 681610
rect 148220 681370 148310 681610
rect 148550 681370 148640 681610
rect 148880 681370 148970 681610
rect 149210 681370 149320 681610
rect 149560 681370 149650 681610
rect 149890 681370 149980 681610
rect 150220 681370 150310 681610
rect 150550 681370 150660 681610
rect 150900 681370 150990 681610
rect 151230 681370 151320 681610
rect 151560 681370 151650 681610
rect 151890 681370 152000 681610
rect 152240 681370 152330 681610
rect 152570 681370 152660 681610
rect 152900 681370 152990 681610
rect 153230 681370 153340 681610
rect 153580 681370 153670 681610
rect 153910 681370 154000 681610
rect 154240 681370 154330 681610
rect 154570 681370 154680 681610
rect 154920 681370 155010 681610
rect 155250 681370 155340 681610
rect 155580 681370 155670 681610
rect 155910 681370 155960 681610
rect 110760 681280 155960 681370
rect 110760 681040 110810 681280
rect 111050 681040 111160 681280
rect 111400 681040 111490 681280
rect 111730 681040 111820 681280
rect 112060 681040 112150 681280
rect 112390 681040 112500 681280
rect 112740 681040 112830 681280
rect 113070 681040 113160 681280
rect 113400 681040 113490 681280
rect 113730 681040 113840 681280
rect 114080 681040 114170 681280
rect 114410 681040 114500 681280
rect 114740 681040 114830 681280
rect 115070 681040 115180 681280
rect 115420 681040 115510 681280
rect 115750 681040 115840 681280
rect 116080 681040 116170 681280
rect 116410 681040 116520 681280
rect 116760 681040 116850 681280
rect 117090 681040 117180 681280
rect 117420 681040 117510 681280
rect 117750 681040 117860 681280
rect 118100 681040 118190 681280
rect 118430 681040 118520 681280
rect 118760 681040 118850 681280
rect 119090 681040 119200 681280
rect 119440 681040 119530 681280
rect 119770 681040 119860 681280
rect 120100 681040 120190 681280
rect 120430 681040 120540 681280
rect 120780 681040 120870 681280
rect 121110 681040 121200 681280
rect 121440 681040 121530 681280
rect 121770 681040 122190 681280
rect 122430 681040 122540 681280
rect 122780 681040 122870 681280
rect 123110 681040 123200 681280
rect 123440 681040 123530 681280
rect 123770 681040 123880 681280
rect 124120 681040 124210 681280
rect 124450 681040 124540 681280
rect 124780 681040 124870 681280
rect 125110 681040 125220 681280
rect 125460 681040 125550 681280
rect 125790 681040 125880 681280
rect 126120 681040 126210 681280
rect 126450 681040 126560 681280
rect 126800 681040 126890 681280
rect 127130 681040 127220 681280
rect 127460 681040 127550 681280
rect 127790 681040 127900 681280
rect 128140 681040 128230 681280
rect 128470 681040 128560 681280
rect 128800 681040 128890 681280
rect 129130 681040 129240 681280
rect 129480 681040 129570 681280
rect 129810 681040 129900 681280
rect 130140 681040 130230 681280
rect 130470 681040 130580 681280
rect 130820 681040 130910 681280
rect 131150 681040 131240 681280
rect 131480 681040 131570 681280
rect 131810 681040 131920 681280
rect 132160 681040 132250 681280
rect 132490 681040 132580 681280
rect 132820 681040 132910 681280
rect 133150 681040 133570 681280
rect 133810 681040 133920 681280
rect 134160 681040 134250 681280
rect 134490 681040 134580 681280
rect 134820 681040 134910 681280
rect 135150 681040 135260 681280
rect 135500 681040 135590 681280
rect 135830 681040 135920 681280
rect 136160 681040 136250 681280
rect 136490 681040 136600 681280
rect 136840 681040 136930 681280
rect 137170 681040 137260 681280
rect 137500 681040 137590 681280
rect 137830 681040 137940 681280
rect 138180 681040 138270 681280
rect 138510 681040 138600 681280
rect 138840 681040 138930 681280
rect 139170 681040 139280 681280
rect 139520 681040 139610 681280
rect 139850 681040 139940 681280
rect 140180 681040 140270 681280
rect 140510 681040 140620 681280
rect 140860 681040 140950 681280
rect 141190 681040 141280 681280
rect 141520 681040 141610 681280
rect 141850 681040 141960 681280
rect 142200 681040 142290 681280
rect 142530 681040 142620 681280
rect 142860 681040 142950 681280
rect 143190 681040 143300 681280
rect 143540 681040 143630 681280
rect 143870 681040 143960 681280
rect 144200 681040 144290 681280
rect 144530 681040 144950 681280
rect 145190 681040 145300 681280
rect 145540 681040 145630 681280
rect 145870 681040 145960 681280
rect 146200 681040 146290 681280
rect 146530 681040 146640 681280
rect 146880 681040 146970 681280
rect 147210 681040 147300 681280
rect 147540 681040 147630 681280
rect 147870 681040 147980 681280
rect 148220 681040 148310 681280
rect 148550 681040 148640 681280
rect 148880 681040 148970 681280
rect 149210 681040 149320 681280
rect 149560 681040 149650 681280
rect 149890 681040 149980 681280
rect 150220 681040 150310 681280
rect 150550 681040 150660 681280
rect 150900 681040 150990 681280
rect 151230 681040 151320 681280
rect 151560 681040 151650 681280
rect 151890 681040 152000 681280
rect 152240 681040 152330 681280
rect 152570 681040 152660 681280
rect 152900 681040 152990 681280
rect 153230 681040 153340 681280
rect 153580 681040 153670 681280
rect 153910 681040 154000 681280
rect 154240 681040 154330 681280
rect 154570 681040 154680 681280
rect 154920 681040 155010 681280
rect 155250 681040 155340 681280
rect 155580 681040 155670 681280
rect 155910 681040 155960 681280
rect 110760 680950 155960 681040
rect 110760 680710 110810 680950
rect 111050 680710 111160 680950
rect 111400 680710 111490 680950
rect 111730 680710 111820 680950
rect 112060 680710 112150 680950
rect 112390 680710 112500 680950
rect 112740 680710 112830 680950
rect 113070 680710 113160 680950
rect 113400 680710 113490 680950
rect 113730 680710 113840 680950
rect 114080 680710 114170 680950
rect 114410 680710 114500 680950
rect 114740 680710 114830 680950
rect 115070 680710 115180 680950
rect 115420 680710 115510 680950
rect 115750 680710 115840 680950
rect 116080 680710 116170 680950
rect 116410 680710 116520 680950
rect 116760 680710 116850 680950
rect 117090 680710 117180 680950
rect 117420 680710 117510 680950
rect 117750 680710 117860 680950
rect 118100 680710 118190 680950
rect 118430 680710 118520 680950
rect 118760 680710 118850 680950
rect 119090 680710 119200 680950
rect 119440 680710 119530 680950
rect 119770 680710 119860 680950
rect 120100 680710 120190 680950
rect 120430 680710 120540 680950
rect 120780 680710 120870 680950
rect 121110 680710 121200 680950
rect 121440 680710 121530 680950
rect 121770 680710 122190 680950
rect 122430 680710 122540 680950
rect 122780 680710 122870 680950
rect 123110 680710 123200 680950
rect 123440 680710 123530 680950
rect 123770 680710 123880 680950
rect 124120 680710 124210 680950
rect 124450 680710 124540 680950
rect 124780 680710 124870 680950
rect 125110 680710 125220 680950
rect 125460 680710 125550 680950
rect 125790 680710 125880 680950
rect 126120 680710 126210 680950
rect 126450 680710 126560 680950
rect 126800 680710 126890 680950
rect 127130 680710 127220 680950
rect 127460 680710 127550 680950
rect 127790 680710 127900 680950
rect 128140 680710 128230 680950
rect 128470 680710 128560 680950
rect 128800 680710 128890 680950
rect 129130 680710 129240 680950
rect 129480 680710 129570 680950
rect 129810 680710 129900 680950
rect 130140 680710 130230 680950
rect 130470 680710 130580 680950
rect 130820 680710 130910 680950
rect 131150 680710 131240 680950
rect 131480 680710 131570 680950
rect 131810 680710 131920 680950
rect 132160 680710 132250 680950
rect 132490 680710 132580 680950
rect 132820 680710 132910 680950
rect 133150 680710 133570 680950
rect 133810 680710 133920 680950
rect 134160 680710 134250 680950
rect 134490 680710 134580 680950
rect 134820 680710 134910 680950
rect 135150 680710 135260 680950
rect 135500 680710 135590 680950
rect 135830 680710 135920 680950
rect 136160 680710 136250 680950
rect 136490 680710 136600 680950
rect 136840 680710 136930 680950
rect 137170 680710 137260 680950
rect 137500 680710 137590 680950
rect 137830 680710 137940 680950
rect 138180 680710 138270 680950
rect 138510 680710 138600 680950
rect 138840 680710 138930 680950
rect 139170 680710 139280 680950
rect 139520 680710 139610 680950
rect 139850 680710 139940 680950
rect 140180 680710 140270 680950
rect 140510 680710 140620 680950
rect 140860 680710 140950 680950
rect 141190 680710 141280 680950
rect 141520 680710 141610 680950
rect 141850 680710 141960 680950
rect 142200 680710 142290 680950
rect 142530 680710 142620 680950
rect 142860 680710 142950 680950
rect 143190 680710 143300 680950
rect 143540 680710 143630 680950
rect 143870 680710 143960 680950
rect 144200 680710 144290 680950
rect 144530 680710 144950 680950
rect 145190 680710 145300 680950
rect 145540 680710 145630 680950
rect 145870 680710 145960 680950
rect 146200 680710 146290 680950
rect 146530 680710 146640 680950
rect 146880 680710 146970 680950
rect 147210 680710 147300 680950
rect 147540 680710 147630 680950
rect 147870 680710 147980 680950
rect 148220 680710 148310 680950
rect 148550 680710 148640 680950
rect 148880 680710 148970 680950
rect 149210 680710 149320 680950
rect 149560 680710 149650 680950
rect 149890 680710 149980 680950
rect 150220 680710 150310 680950
rect 150550 680710 150660 680950
rect 150900 680710 150990 680950
rect 151230 680710 151320 680950
rect 151560 680710 151650 680950
rect 151890 680710 152000 680950
rect 152240 680710 152330 680950
rect 152570 680710 152660 680950
rect 152900 680710 152990 680950
rect 153230 680710 153340 680950
rect 153580 680710 153670 680950
rect 153910 680710 154000 680950
rect 154240 680710 154330 680950
rect 154570 680710 154680 680950
rect 154920 680710 155010 680950
rect 155250 680710 155340 680950
rect 155580 680710 155670 680950
rect 155910 680710 155960 680950
rect 110760 680600 155960 680710
rect 110760 680360 110810 680600
rect 111050 680360 111160 680600
rect 111400 680360 111490 680600
rect 111730 680360 111820 680600
rect 112060 680360 112150 680600
rect 112390 680360 112500 680600
rect 112740 680360 112830 680600
rect 113070 680360 113160 680600
rect 113400 680360 113490 680600
rect 113730 680360 113840 680600
rect 114080 680360 114170 680600
rect 114410 680360 114500 680600
rect 114740 680360 114830 680600
rect 115070 680360 115180 680600
rect 115420 680360 115510 680600
rect 115750 680360 115840 680600
rect 116080 680360 116170 680600
rect 116410 680360 116520 680600
rect 116760 680360 116850 680600
rect 117090 680360 117180 680600
rect 117420 680360 117510 680600
rect 117750 680360 117860 680600
rect 118100 680360 118190 680600
rect 118430 680360 118520 680600
rect 118760 680360 118850 680600
rect 119090 680360 119200 680600
rect 119440 680360 119530 680600
rect 119770 680360 119860 680600
rect 120100 680360 120190 680600
rect 120430 680360 120540 680600
rect 120780 680360 120870 680600
rect 121110 680360 121200 680600
rect 121440 680360 121530 680600
rect 121770 680360 122190 680600
rect 122430 680360 122540 680600
rect 122780 680360 122870 680600
rect 123110 680360 123200 680600
rect 123440 680360 123530 680600
rect 123770 680360 123880 680600
rect 124120 680360 124210 680600
rect 124450 680360 124540 680600
rect 124780 680360 124870 680600
rect 125110 680360 125220 680600
rect 125460 680360 125550 680600
rect 125790 680360 125880 680600
rect 126120 680360 126210 680600
rect 126450 680360 126560 680600
rect 126800 680360 126890 680600
rect 127130 680360 127220 680600
rect 127460 680360 127550 680600
rect 127790 680360 127900 680600
rect 128140 680360 128230 680600
rect 128470 680360 128560 680600
rect 128800 680360 128890 680600
rect 129130 680360 129240 680600
rect 129480 680360 129570 680600
rect 129810 680360 129900 680600
rect 130140 680360 130230 680600
rect 130470 680360 130580 680600
rect 130820 680360 130910 680600
rect 131150 680360 131240 680600
rect 131480 680360 131570 680600
rect 131810 680360 131920 680600
rect 132160 680360 132250 680600
rect 132490 680360 132580 680600
rect 132820 680360 132910 680600
rect 133150 680360 133570 680600
rect 133810 680360 133920 680600
rect 134160 680360 134250 680600
rect 134490 680360 134580 680600
rect 134820 680360 134910 680600
rect 135150 680360 135260 680600
rect 135500 680360 135590 680600
rect 135830 680360 135920 680600
rect 136160 680360 136250 680600
rect 136490 680360 136600 680600
rect 136840 680360 136930 680600
rect 137170 680360 137260 680600
rect 137500 680360 137590 680600
rect 137830 680360 137940 680600
rect 138180 680360 138270 680600
rect 138510 680360 138600 680600
rect 138840 680360 138930 680600
rect 139170 680360 139280 680600
rect 139520 680360 139610 680600
rect 139850 680360 139940 680600
rect 140180 680360 140270 680600
rect 140510 680360 140620 680600
rect 140860 680360 140950 680600
rect 141190 680360 141280 680600
rect 141520 680360 141610 680600
rect 141850 680360 141960 680600
rect 142200 680360 142290 680600
rect 142530 680360 142620 680600
rect 142860 680360 142950 680600
rect 143190 680360 143300 680600
rect 143540 680360 143630 680600
rect 143870 680360 143960 680600
rect 144200 680360 144290 680600
rect 144530 680360 144950 680600
rect 145190 680360 145300 680600
rect 145540 680360 145630 680600
rect 145870 680360 145960 680600
rect 146200 680360 146290 680600
rect 146530 680360 146640 680600
rect 146880 680360 146970 680600
rect 147210 680360 147300 680600
rect 147540 680360 147630 680600
rect 147870 680360 147980 680600
rect 148220 680360 148310 680600
rect 148550 680360 148640 680600
rect 148880 680360 148970 680600
rect 149210 680360 149320 680600
rect 149560 680360 149650 680600
rect 149890 680360 149980 680600
rect 150220 680360 150310 680600
rect 150550 680360 150660 680600
rect 150900 680360 150990 680600
rect 151230 680360 151320 680600
rect 151560 680360 151650 680600
rect 151890 680360 152000 680600
rect 152240 680360 152330 680600
rect 152570 680360 152660 680600
rect 152900 680360 152990 680600
rect 153230 680360 153340 680600
rect 153580 680360 153670 680600
rect 153910 680360 154000 680600
rect 154240 680360 154330 680600
rect 154570 680360 154680 680600
rect 154920 680360 155010 680600
rect 155250 680360 155340 680600
rect 155580 680360 155670 680600
rect 155910 680360 155960 680600
rect 110760 680270 155960 680360
rect 110760 680030 110810 680270
rect 111050 680030 111160 680270
rect 111400 680030 111490 680270
rect 111730 680030 111820 680270
rect 112060 680030 112150 680270
rect 112390 680030 112500 680270
rect 112740 680030 112830 680270
rect 113070 680030 113160 680270
rect 113400 680030 113490 680270
rect 113730 680030 113840 680270
rect 114080 680030 114170 680270
rect 114410 680030 114500 680270
rect 114740 680030 114830 680270
rect 115070 680030 115180 680270
rect 115420 680030 115510 680270
rect 115750 680030 115840 680270
rect 116080 680030 116170 680270
rect 116410 680030 116520 680270
rect 116760 680030 116850 680270
rect 117090 680030 117180 680270
rect 117420 680030 117510 680270
rect 117750 680030 117860 680270
rect 118100 680030 118190 680270
rect 118430 680030 118520 680270
rect 118760 680030 118850 680270
rect 119090 680030 119200 680270
rect 119440 680030 119530 680270
rect 119770 680030 119860 680270
rect 120100 680030 120190 680270
rect 120430 680030 120540 680270
rect 120780 680030 120870 680270
rect 121110 680030 121200 680270
rect 121440 680030 121530 680270
rect 121770 680030 122190 680270
rect 122430 680030 122540 680270
rect 122780 680030 122870 680270
rect 123110 680030 123200 680270
rect 123440 680030 123530 680270
rect 123770 680030 123880 680270
rect 124120 680030 124210 680270
rect 124450 680030 124540 680270
rect 124780 680030 124870 680270
rect 125110 680030 125220 680270
rect 125460 680030 125550 680270
rect 125790 680030 125880 680270
rect 126120 680030 126210 680270
rect 126450 680030 126560 680270
rect 126800 680030 126890 680270
rect 127130 680030 127220 680270
rect 127460 680030 127550 680270
rect 127790 680030 127900 680270
rect 128140 680030 128230 680270
rect 128470 680030 128560 680270
rect 128800 680030 128890 680270
rect 129130 680030 129240 680270
rect 129480 680030 129570 680270
rect 129810 680030 129900 680270
rect 130140 680030 130230 680270
rect 130470 680030 130580 680270
rect 130820 680030 130910 680270
rect 131150 680030 131240 680270
rect 131480 680030 131570 680270
rect 131810 680030 131920 680270
rect 132160 680030 132250 680270
rect 132490 680030 132580 680270
rect 132820 680030 132910 680270
rect 133150 680030 133570 680270
rect 133810 680030 133920 680270
rect 134160 680030 134250 680270
rect 134490 680030 134580 680270
rect 134820 680030 134910 680270
rect 135150 680030 135260 680270
rect 135500 680030 135590 680270
rect 135830 680030 135920 680270
rect 136160 680030 136250 680270
rect 136490 680030 136600 680270
rect 136840 680030 136930 680270
rect 137170 680030 137260 680270
rect 137500 680030 137590 680270
rect 137830 680030 137940 680270
rect 138180 680030 138270 680270
rect 138510 680030 138600 680270
rect 138840 680030 138930 680270
rect 139170 680030 139280 680270
rect 139520 680030 139610 680270
rect 139850 680030 139940 680270
rect 140180 680030 140270 680270
rect 140510 680030 140620 680270
rect 140860 680030 140950 680270
rect 141190 680030 141280 680270
rect 141520 680030 141610 680270
rect 141850 680030 141960 680270
rect 142200 680030 142290 680270
rect 142530 680030 142620 680270
rect 142860 680030 142950 680270
rect 143190 680030 143300 680270
rect 143540 680030 143630 680270
rect 143870 680030 143960 680270
rect 144200 680030 144290 680270
rect 144530 680030 144950 680270
rect 145190 680030 145300 680270
rect 145540 680030 145630 680270
rect 145870 680030 145960 680270
rect 146200 680030 146290 680270
rect 146530 680030 146640 680270
rect 146880 680030 146970 680270
rect 147210 680030 147300 680270
rect 147540 680030 147630 680270
rect 147870 680030 147980 680270
rect 148220 680030 148310 680270
rect 148550 680030 148640 680270
rect 148880 680030 148970 680270
rect 149210 680030 149320 680270
rect 149560 680030 149650 680270
rect 149890 680030 149980 680270
rect 150220 680030 150310 680270
rect 150550 680030 150660 680270
rect 150900 680030 150990 680270
rect 151230 680030 151320 680270
rect 151560 680030 151650 680270
rect 151890 680030 152000 680270
rect 152240 680030 152330 680270
rect 152570 680030 152660 680270
rect 152900 680030 152990 680270
rect 153230 680030 153340 680270
rect 153580 680030 153670 680270
rect 153910 680030 154000 680270
rect 154240 680030 154330 680270
rect 154570 680030 154680 680270
rect 154920 680030 155010 680270
rect 155250 680030 155340 680270
rect 155580 680030 155670 680270
rect 155910 680030 155960 680270
rect 110760 679940 155960 680030
rect 110760 679700 110810 679940
rect 111050 679700 111160 679940
rect 111400 679700 111490 679940
rect 111730 679700 111820 679940
rect 112060 679700 112150 679940
rect 112390 679700 112500 679940
rect 112740 679700 112830 679940
rect 113070 679700 113160 679940
rect 113400 679700 113490 679940
rect 113730 679700 113840 679940
rect 114080 679700 114170 679940
rect 114410 679700 114500 679940
rect 114740 679700 114830 679940
rect 115070 679700 115180 679940
rect 115420 679700 115510 679940
rect 115750 679700 115840 679940
rect 116080 679700 116170 679940
rect 116410 679700 116520 679940
rect 116760 679700 116850 679940
rect 117090 679700 117180 679940
rect 117420 679700 117510 679940
rect 117750 679700 117860 679940
rect 118100 679700 118190 679940
rect 118430 679700 118520 679940
rect 118760 679700 118850 679940
rect 119090 679700 119200 679940
rect 119440 679700 119530 679940
rect 119770 679700 119860 679940
rect 120100 679700 120190 679940
rect 120430 679700 120540 679940
rect 120780 679700 120870 679940
rect 121110 679700 121200 679940
rect 121440 679700 121530 679940
rect 121770 679700 122190 679940
rect 122430 679700 122540 679940
rect 122780 679700 122870 679940
rect 123110 679700 123200 679940
rect 123440 679700 123530 679940
rect 123770 679700 123880 679940
rect 124120 679700 124210 679940
rect 124450 679700 124540 679940
rect 124780 679700 124870 679940
rect 125110 679700 125220 679940
rect 125460 679700 125550 679940
rect 125790 679700 125880 679940
rect 126120 679700 126210 679940
rect 126450 679700 126560 679940
rect 126800 679700 126890 679940
rect 127130 679700 127220 679940
rect 127460 679700 127550 679940
rect 127790 679700 127900 679940
rect 128140 679700 128230 679940
rect 128470 679700 128560 679940
rect 128800 679700 128890 679940
rect 129130 679700 129240 679940
rect 129480 679700 129570 679940
rect 129810 679700 129900 679940
rect 130140 679700 130230 679940
rect 130470 679700 130580 679940
rect 130820 679700 130910 679940
rect 131150 679700 131240 679940
rect 131480 679700 131570 679940
rect 131810 679700 131920 679940
rect 132160 679700 132250 679940
rect 132490 679700 132580 679940
rect 132820 679700 132910 679940
rect 133150 679700 133570 679940
rect 133810 679700 133920 679940
rect 134160 679700 134250 679940
rect 134490 679700 134580 679940
rect 134820 679700 134910 679940
rect 135150 679700 135260 679940
rect 135500 679700 135590 679940
rect 135830 679700 135920 679940
rect 136160 679700 136250 679940
rect 136490 679700 136600 679940
rect 136840 679700 136930 679940
rect 137170 679700 137260 679940
rect 137500 679700 137590 679940
rect 137830 679700 137940 679940
rect 138180 679700 138270 679940
rect 138510 679700 138600 679940
rect 138840 679700 138930 679940
rect 139170 679700 139280 679940
rect 139520 679700 139610 679940
rect 139850 679700 139940 679940
rect 140180 679700 140270 679940
rect 140510 679700 140620 679940
rect 140860 679700 140950 679940
rect 141190 679700 141280 679940
rect 141520 679700 141610 679940
rect 141850 679700 141960 679940
rect 142200 679700 142290 679940
rect 142530 679700 142620 679940
rect 142860 679700 142950 679940
rect 143190 679700 143300 679940
rect 143540 679700 143630 679940
rect 143870 679700 143960 679940
rect 144200 679700 144290 679940
rect 144530 679700 144950 679940
rect 145190 679700 145300 679940
rect 145540 679700 145630 679940
rect 145870 679700 145960 679940
rect 146200 679700 146290 679940
rect 146530 679700 146640 679940
rect 146880 679700 146970 679940
rect 147210 679700 147300 679940
rect 147540 679700 147630 679940
rect 147870 679700 147980 679940
rect 148220 679700 148310 679940
rect 148550 679700 148640 679940
rect 148880 679700 148970 679940
rect 149210 679700 149320 679940
rect 149560 679700 149650 679940
rect 149890 679700 149980 679940
rect 150220 679700 150310 679940
rect 150550 679700 150660 679940
rect 150900 679700 150990 679940
rect 151230 679700 151320 679940
rect 151560 679700 151650 679940
rect 151890 679700 152000 679940
rect 152240 679700 152330 679940
rect 152570 679700 152660 679940
rect 152900 679700 152990 679940
rect 153230 679700 153340 679940
rect 153580 679700 153670 679940
rect 153910 679700 154000 679940
rect 154240 679700 154330 679940
rect 154570 679700 154680 679940
rect 154920 679700 155010 679940
rect 155250 679700 155340 679940
rect 155580 679700 155670 679940
rect 155910 679700 155960 679940
rect 110760 679610 155960 679700
rect 110760 679370 110810 679610
rect 111050 679370 111160 679610
rect 111400 679370 111490 679610
rect 111730 679370 111820 679610
rect 112060 679370 112150 679610
rect 112390 679370 112500 679610
rect 112740 679370 112830 679610
rect 113070 679370 113160 679610
rect 113400 679370 113490 679610
rect 113730 679370 113840 679610
rect 114080 679370 114170 679610
rect 114410 679370 114500 679610
rect 114740 679370 114830 679610
rect 115070 679370 115180 679610
rect 115420 679370 115510 679610
rect 115750 679370 115840 679610
rect 116080 679370 116170 679610
rect 116410 679370 116520 679610
rect 116760 679370 116850 679610
rect 117090 679370 117180 679610
rect 117420 679370 117510 679610
rect 117750 679370 117860 679610
rect 118100 679370 118190 679610
rect 118430 679370 118520 679610
rect 118760 679370 118850 679610
rect 119090 679370 119200 679610
rect 119440 679370 119530 679610
rect 119770 679370 119860 679610
rect 120100 679370 120190 679610
rect 120430 679370 120540 679610
rect 120780 679370 120870 679610
rect 121110 679370 121200 679610
rect 121440 679370 121530 679610
rect 121770 679370 122190 679610
rect 122430 679370 122540 679610
rect 122780 679370 122870 679610
rect 123110 679370 123200 679610
rect 123440 679370 123530 679610
rect 123770 679370 123880 679610
rect 124120 679370 124210 679610
rect 124450 679370 124540 679610
rect 124780 679370 124870 679610
rect 125110 679370 125220 679610
rect 125460 679370 125550 679610
rect 125790 679370 125880 679610
rect 126120 679370 126210 679610
rect 126450 679370 126560 679610
rect 126800 679370 126890 679610
rect 127130 679370 127220 679610
rect 127460 679370 127550 679610
rect 127790 679370 127900 679610
rect 128140 679370 128230 679610
rect 128470 679370 128560 679610
rect 128800 679370 128890 679610
rect 129130 679370 129240 679610
rect 129480 679370 129570 679610
rect 129810 679370 129900 679610
rect 130140 679370 130230 679610
rect 130470 679370 130580 679610
rect 130820 679370 130910 679610
rect 131150 679370 131240 679610
rect 131480 679370 131570 679610
rect 131810 679370 131920 679610
rect 132160 679370 132250 679610
rect 132490 679370 132580 679610
rect 132820 679370 132910 679610
rect 133150 679370 133570 679610
rect 133810 679370 133920 679610
rect 134160 679370 134250 679610
rect 134490 679370 134580 679610
rect 134820 679370 134910 679610
rect 135150 679370 135260 679610
rect 135500 679370 135590 679610
rect 135830 679370 135920 679610
rect 136160 679370 136250 679610
rect 136490 679370 136600 679610
rect 136840 679370 136930 679610
rect 137170 679370 137260 679610
rect 137500 679370 137590 679610
rect 137830 679370 137940 679610
rect 138180 679370 138270 679610
rect 138510 679370 138600 679610
rect 138840 679370 138930 679610
rect 139170 679370 139280 679610
rect 139520 679370 139610 679610
rect 139850 679370 139940 679610
rect 140180 679370 140270 679610
rect 140510 679370 140620 679610
rect 140860 679370 140950 679610
rect 141190 679370 141280 679610
rect 141520 679370 141610 679610
rect 141850 679370 141960 679610
rect 142200 679370 142290 679610
rect 142530 679370 142620 679610
rect 142860 679370 142950 679610
rect 143190 679370 143300 679610
rect 143540 679370 143630 679610
rect 143870 679370 143960 679610
rect 144200 679370 144290 679610
rect 144530 679370 144950 679610
rect 145190 679370 145300 679610
rect 145540 679370 145630 679610
rect 145870 679370 145960 679610
rect 146200 679370 146290 679610
rect 146530 679370 146640 679610
rect 146880 679370 146970 679610
rect 147210 679370 147300 679610
rect 147540 679370 147630 679610
rect 147870 679370 147980 679610
rect 148220 679370 148310 679610
rect 148550 679370 148640 679610
rect 148880 679370 148970 679610
rect 149210 679370 149320 679610
rect 149560 679370 149650 679610
rect 149890 679370 149980 679610
rect 150220 679370 150310 679610
rect 150550 679370 150660 679610
rect 150900 679370 150990 679610
rect 151230 679370 151320 679610
rect 151560 679370 151650 679610
rect 151890 679370 152000 679610
rect 152240 679370 152330 679610
rect 152570 679370 152660 679610
rect 152900 679370 152990 679610
rect 153230 679370 153340 679610
rect 153580 679370 153670 679610
rect 153910 679370 154000 679610
rect 154240 679370 154330 679610
rect 154570 679370 154680 679610
rect 154920 679370 155010 679610
rect 155250 679370 155340 679610
rect 155580 679370 155670 679610
rect 155910 679370 155960 679610
rect 110760 679260 155960 679370
rect 16197 678980 108640 679147
rect 16197 678740 107220 678980
rect 107480 678740 107580 678980
rect 107840 678740 107940 678980
rect 108200 678740 108300 678980
rect 108560 678740 108640 678980
rect 16197 678640 108640 678740
rect 16197 678400 107220 678640
rect 107480 678400 107580 678640
rect 107840 678400 107940 678640
rect 108200 678400 108300 678640
rect 108560 678400 108640 678640
rect 16197 678300 108640 678400
rect 16197 678060 107220 678300
rect 107480 678060 107580 678300
rect 107840 678060 107940 678300
rect 108200 678060 108300 678300
rect 108560 678060 108640 678300
rect 16197 677960 108640 678060
rect 16197 677720 107220 677960
rect 107480 677720 107580 677960
rect 107840 677720 107940 677960
rect 108200 677720 108300 677960
rect 108560 677720 108640 677960
rect 16197 677620 108640 677720
rect 16197 677380 107220 677620
rect 107480 677380 107580 677620
rect 107840 677380 107940 677620
rect 108200 677380 108300 677620
rect 108560 677380 108640 677620
rect 16197 677280 108640 677380
rect 16197 677040 107220 677280
rect 107480 677040 107580 677280
rect 107840 677040 107940 677280
rect 108200 677040 108300 677280
rect 108560 677040 108640 677280
rect 16197 676940 108640 677040
rect 16197 676700 107220 676940
rect 107480 676700 107580 676940
rect 107840 676700 107940 676940
rect 108200 676700 108300 676940
rect 108560 676700 108640 676940
rect 16197 676600 108640 676700
rect 16197 676360 107220 676600
rect 107480 676360 107580 676600
rect 107840 676360 107940 676600
rect 108200 676360 108300 676600
rect 108560 676360 108640 676600
rect 16197 676260 108640 676360
rect 16197 676020 107220 676260
rect 107480 676020 107580 676260
rect 107840 676020 107940 676260
rect 108200 676020 108300 676260
rect 108560 676020 108640 676260
rect 16197 675920 108640 676020
rect 16197 675680 107220 675920
rect 107480 675680 107580 675920
rect 107840 675680 107940 675920
rect 108200 675680 108300 675920
rect 108560 675680 108640 675920
rect 16197 675580 108640 675680
rect 16197 675340 107220 675580
rect 107480 675340 107580 675580
rect 107840 675340 107940 675580
rect 108200 675340 108300 675580
rect 108560 675340 108640 675580
rect 16197 675240 108640 675340
rect 16197 675000 107220 675240
rect 107480 675000 107580 675240
rect 107840 675000 107940 675240
rect 108200 675000 108300 675240
rect 108560 675000 108640 675240
rect 16197 674900 108640 675000
rect 16197 674660 107220 674900
rect 107480 674660 107580 674900
rect 107840 674660 107940 674900
rect 108200 674660 108300 674900
rect 108560 674660 108640 674900
rect 16197 674560 108640 674660
rect 16197 674320 107220 674560
rect 107480 674320 107580 674560
rect 107840 674320 107940 674560
rect 108200 674320 108300 674560
rect 108560 674320 108640 674560
rect 16197 674152 108640 674320
rect 110760 679020 110810 679260
rect 111050 679020 111160 679260
rect 111400 679020 111490 679260
rect 111730 679020 111820 679260
rect 112060 679020 112150 679260
rect 112390 679020 112500 679260
rect 112740 679020 112830 679260
rect 113070 679020 113160 679260
rect 113400 679020 113490 679260
rect 113730 679020 113840 679260
rect 114080 679020 114170 679260
rect 114410 679020 114500 679260
rect 114740 679020 114830 679260
rect 115070 679020 115180 679260
rect 115420 679020 115510 679260
rect 115750 679020 115840 679260
rect 116080 679020 116170 679260
rect 116410 679020 116520 679260
rect 116760 679020 116850 679260
rect 117090 679020 117180 679260
rect 117420 679020 117510 679260
rect 117750 679020 117860 679260
rect 118100 679020 118190 679260
rect 118430 679020 118520 679260
rect 118760 679020 118850 679260
rect 119090 679020 119200 679260
rect 119440 679020 119530 679260
rect 119770 679020 119860 679260
rect 120100 679020 120190 679260
rect 120430 679020 120540 679260
rect 120780 679020 120870 679260
rect 121110 679020 121200 679260
rect 121440 679020 121530 679260
rect 121770 679020 122190 679260
rect 122430 679020 122540 679260
rect 122780 679020 122870 679260
rect 123110 679020 123200 679260
rect 123440 679020 123530 679260
rect 123770 679020 123880 679260
rect 124120 679020 124210 679260
rect 124450 679020 124540 679260
rect 124780 679020 124870 679260
rect 125110 679020 125220 679260
rect 125460 679020 125550 679260
rect 125790 679020 125880 679260
rect 126120 679020 126210 679260
rect 126450 679020 126560 679260
rect 126800 679020 126890 679260
rect 127130 679020 127220 679260
rect 127460 679020 127550 679260
rect 127790 679020 127900 679260
rect 128140 679020 128230 679260
rect 128470 679020 128560 679260
rect 128800 679020 128890 679260
rect 129130 679020 129240 679260
rect 129480 679020 129570 679260
rect 129810 679020 129900 679260
rect 130140 679020 130230 679260
rect 130470 679020 130580 679260
rect 130820 679020 130910 679260
rect 131150 679020 131240 679260
rect 131480 679020 131570 679260
rect 131810 679020 131920 679260
rect 132160 679020 132250 679260
rect 132490 679020 132580 679260
rect 132820 679020 132910 679260
rect 133150 679020 133570 679260
rect 133810 679020 133920 679260
rect 134160 679020 134250 679260
rect 134490 679020 134580 679260
rect 134820 679020 134910 679260
rect 135150 679020 135260 679260
rect 135500 679020 135590 679260
rect 135830 679020 135920 679260
rect 136160 679020 136250 679260
rect 136490 679020 136600 679260
rect 136840 679020 136930 679260
rect 137170 679020 137260 679260
rect 137500 679020 137590 679260
rect 137830 679020 137940 679260
rect 138180 679020 138270 679260
rect 138510 679020 138600 679260
rect 138840 679020 138930 679260
rect 139170 679020 139280 679260
rect 139520 679020 139610 679260
rect 139850 679020 139940 679260
rect 140180 679020 140270 679260
rect 140510 679020 140620 679260
rect 140860 679020 140950 679260
rect 141190 679020 141280 679260
rect 141520 679020 141610 679260
rect 141850 679020 141960 679260
rect 142200 679020 142290 679260
rect 142530 679020 142620 679260
rect 142860 679020 142950 679260
rect 143190 679020 143300 679260
rect 143540 679020 143630 679260
rect 143870 679020 143960 679260
rect 144200 679020 144290 679260
rect 144530 679020 144950 679260
rect 145190 679020 145300 679260
rect 145540 679020 145630 679260
rect 145870 679020 145960 679260
rect 146200 679020 146290 679260
rect 146530 679020 146640 679260
rect 146880 679020 146970 679260
rect 147210 679020 147300 679260
rect 147540 679020 147630 679260
rect 147870 679020 147980 679260
rect 148220 679020 148310 679260
rect 148550 679020 148640 679260
rect 148880 679020 148970 679260
rect 149210 679020 149320 679260
rect 149560 679020 149650 679260
rect 149890 679020 149980 679260
rect 150220 679020 150310 679260
rect 150550 679020 150660 679260
rect 150900 679020 150990 679260
rect 151230 679020 151320 679260
rect 151560 679020 151650 679260
rect 151890 679020 152000 679260
rect 152240 679020 152330 679260
rect 152570 679020 152660 679260
rect 152900 679020 152990 679260
rect 153230 679020 153340 679260
rect 153580 679020 153670 679260
rect 153910 679020 154000 679260
rect 154240 679020 154330 679260
rect 154570 679020 154680 679260
rect 154920 679020 155010 679260
rect 155250 679020 155340 679260
rect 155580 679020 155670 679260
rect 155910 679020 155960 679260
rect 110760 678930 155960 679020
rect 110760 678690 110810 678930
rect 111050 678690 111160 678930
rect 111400 678690 111490 678930
rect 111730 678690 111820 678930
rect 112060 678690 112150 678930
rect 112390 678690 112500 678930
rect 112740 678690 112830 678930
rect 113070 678690 113160 678930
rect 113400 678690 113490 678930
rect 113730 678690 113840 678930
rect 114080 678690 114170 678930
rect 114410 678690 114500 678930
rect 114740 678690 114830 678930
rect 115070 678690 115180 678930
rect 115420 678690 115510 678930
rect 115750 678690 115840 678930
rect 116080 678690 116170 678930
rect 116410 678690 116520 678930
rect 116760 678690 116850 678930
rect 117090 678690 117180 678930
rect 117420 678690 117510 678930
rect 117750 678690 117860 678930
rect 118100 678690 118190 678930
rect 118430 678690 118520 678930
rect 118760 678690 118850 678930
rect 119090 678690 119200 678930
rect 119440 678690 119530 678930
rect 119770 678690 119860 678930
rect 120100 678690 120190 678930
rect 120430 678690 120540 678930
rect 120780 678690 120870 678930
rect 121110 678690 121200 678930
rect 121440 678690 121530 678930
rect 121770 678690 122190 678930
rect 122430 678690 122540 678930
rect 122780 678690 122870 678930
rect 123110 678690 123200 678930
rect 123440 678690 123530 678930
rect 123770 678690 123880 678930
rect 124120 678690 124210 678930
rect 124450 678690 124540 678930
rect 124780 678690 124870 678930
rect 125110 678690 125220 678930
rect 125460 678690 125550 678930
rect 125790 678690 125880 678930
rect 126120 678690 126210 678930
rect 126450 678690 126560 678930
rect 126800 678690 126890 678930
rect 127130 678690 127220 678930
rect 127460 678690 127550 678930
rect 127790 678690 127900 678930
rect 128140 678690 128230 678930
rect 128470 678690 128560 678930
rect 128800 678690 128890 678930
rect 129130 678690 129240 678930
rect 129480 678690 129570 678930
rect 129810 678690 129900 678930
rect 130140 678690 130230 678930
rect 130470 678690 130580 678930
rect 130820 678690 130910 678930
rect 131150 678690 131240 678930
rect 131480 678690 131570 678930
rect 131810 678690 131920 678930
rect 132160 678690 132250 678930
rect 132490 678690 132580 678930
rect 132820 678690 132910 678930
rect 133150 678690 133570 678930
rect 133810 678690 133920 678930
rect 134160 678690 134250 678930
rect 134490 678690 134580 678930
rect 134820 678690 134910 678930
rect 135150 678690 135260 678930
rect 135500 678690 135590 678930
rect 135830 678690 135920 678930
rect 136160 678690 136250 678930
rect 136490 678690 136600 678930
rect 136840 678690 136930 678930
rect 137170 678690 137260 678930
rect 137500 678690 137590 678930
rect 137830 678690 137940 678930
rect 138180 678690 138270 678930
rect 138510 678690 138600 678930
rect 138840 678690 138930 678930
rect 139170 678690 139280 678930
rect 139520 678690 139610 678930
rect 139850 678690 139940 678930
rect 140180 678690 140270 678930
rect 140510 678690 140620 678930
rect 140860 678690 140950 678930
rect 141190 678690 141280 678930
rect 141520 678690 141610 678930
rect 141850 678690 141960 678930
rect 142200 678690 142290 678930
rect 142530 678690 142620 678930
rect 142860 678690 142950 678930
rect 143190 678690 143300 678930
rect 143540 678690 143630 678930
rect 143870 678690 143960 678930
rect 144200 678690 144290 678930
rect 144530 678690 144950 678930
rect 145190 678690 145300 678930
rect 145540 678690 145630 678930
rect 145870 678690 145960 678930
rect 146200 678690 146290 678930
rect 146530 678690 146640 678930
rect 146880 678690 146970 678930
rect 147210 678690 147300 678930
rect 147540 678690 147630 678930
rect 147870 678690 147980 678930
rect 148220 678690 148310 678930
rect 148550 678690 148640 678930
rect 148880 678690 148970 678930
rect 149210 678690 149320 678930
rect 149560 678690 149650 678930
rect 149890 678690 149980 678930
rect 150220 678690 150310 678930
rect 150550 678690 150660 678930
rect 150900 678690 150990 678930
rect 151230 678690 151320 678930
rect 151560 678690 151650 678930
rect 151890 678690 152000 678930
rect 152240 678690 152330 678930
rect 152570 678690 152660 678930
rect 152900 678690 152990 678930
rect 153230 678690 153340 678930
rect 153580 678690 153670 678930
rect 153910 678690 154000 678930
rect 154240 678690 154330 678930
rect 154570 678690 154680 678930
rect 154920 678690 155010 678930
rect 155250 678690 155340 678930
rect 155580 678690 155670 678930
rect 155910 678690 155960 678930
rect 110760 678600 155960 678690
rect 110760 678360 110810 678600
rect 111050 678360 111160 678600
rect 111400 678360 111490 678600
rect 111730 678360 111820 678600
rect 112060 678360 112150 678600
rect 112390 678360 112500 678600
rect 112740 678360 112830 678600
rect 113070 678360 113160 678600
rect 113400 678360 113490 678600
rect 113730 678360 113840 678600
rect 114080 678360 114170 678600
rect 114410 678360 114500 678600
rect 114740 678360 114830 678600
rect 115070 678360 115180 678600
rect 115420 678360 115510 678600
rect 115750 678360 115840 678600
rect 116080 678360 116170 678600
rect 116410 678360 116520 678600
rect 116760 678360 116850 678600
rect 117090 678360 117180 678600
rect 117420 678360 117510 678600
rect 117750 678360 117860 678600
rect 118100 678360 118190 678600
rect 118430 678360 118520 678600
rect 118760 678360 118850 678600
rect 119090 678360 119200 678600
rect 119440 678360 119530 678600
rect 119770 678360 119860 678600
rect 120100 678360 120190 678600
rect 120430 678360 120540 678600
rect 120780 678360 120870 678600
rect 121110 678360 121200 678600
rect 121440 678360 121530 678600
rect 121770 678360 122190 678600
rect 122430 678360 122540 678600
rect 122780 678360 122870 678600
rect 123110 678360 123200 678600
rect 123440 678360 123530 678600
rect 123770 678360 123880 678600
rect 124120 678360 124210 678600
rect 124450 678360 124540 678600
rect 124780 678360 124870 678600
rect 125110 678360 125220 678600
rect 125460 678360 125550 678600
rect 125790 678360 125880 678600
rect 126120 678360 126210 678600
rect 126450 678360 126560 678600
rect 126800 678360 126890 678600
rect 127130 678360 127220 678600
rect 127460 678360 127550 678600
rect 127790 678360 127900 678600
rect 128140 678360 128230 678600
rect 128470 678360 128560 678600
rect 128800 678360 128890 678600
rect 129130 678360 129240 678600
rect 129480 678360 129570 678600
rect 129810 678360 129900 678600
rect 130140 678360 130230 678600
rect 130470 678360 130580 678600
rect 130820 678360 130910 678600
rect 131150 678360 131240 678600
rect 131480 678360 131570 678600
rect 131810 678360 131920 678600
rect 132160 678360 132250 678600
rect 132490 678360 132580 678600
rect 132820 678360 132910 678600
rect 133150 678360 133570 678600
rect 133810 678360 133920 678600
rect 134160 678360 134250 678600
rect 134490 678360 134580 678600
rect 134820 678360 134910 678600
rect 135150 678360 135260 678600
rect 135500 678360 135590 678600
rect 135830 678360 135920 678600
rect 136160 678360 136250 678600
rect 136490 678360 136600 678600
rect 136840 678360 136930 678600
rect 137170 678360 137260 678600
rect 137500 678360 137590 678600
rect 137830 678360 137940 678600
rect 138180 678360 138270 678600
rect 138510 678360 138600 678600
rect 138840 678360 138930 678600
rect 139170 678360 139280 678600
rect 139520 678360 139610 678600
rect 139850 678360 139940 678600
rect 140180 678360 140270 678600
rect 140510 678360 140620 678600
rect 140860 678360 140950 678600
rect 141190 678360 141280 678600
rect 141520 678360 141610 678600
rect 141850 678360 141960 678600
rect 142200 678360 142290 678600
rect 142530 678360 142620 678600
rect 142860 678360 142950 678600
rect 143190 678360 143300 678600
rect 143540 678360 143630 678600
rect 143870 678360 143960 678600
rect 144200 678360 144290 678600
rect 144530 678360 144950 678600
rect 145190 678360 145300 678600
rect 145540 678360 145630 678600
rect 145870 678360 145960 678600
rect 146200 678360 146290 678600
rect 146530 678360 146640 678600
rect 146880 678360 146970 678600
rect 147210 678360 147300 678600
rect 147540 678360 147630 678600
rect 147870 678360 147980 678600
rect 148220 678360 148310 678600
rect 148550 678360 148640 678600
rect 148880 678360 148970 678600
rect 149210 678360 149320 678600
rect 149560 678360 149650 678600
rect 149890 678360 149980 678600
rect 150220 678360 150310 678600
rect 150550 678360 150660 678600
rect 150900 678360 150990 678600
rect 151230 678360 151320 678600
rect 151560 678360 151650 678600
rect 151890 678360 152000 678600
rect 152240 678360 152330 678600
rect 152570 678360 152660 678600
rect 152900 678360 152990 678600
rect 153230 678360 153340 678600
rect 153580 678360 153670 678600
rect 153910 678360 154000 678600
rect 154240 678360 154330 678600
rect 154570 678360 154680 678600
rect 154920 678360 155010 678600
rect 155250 678360 155340 678600
rect 155580 678360 155670 678600
rect 155910 678360 155960 678600
rect 110760 678270 155960 678360
rect 110760 678030 110810 678270
rect 111050 678030 111160 678270
rect 111400 678030 111490 678270
rect 111730 678030 111820 678270
rect 112060 678030 112150 678270
rect 112390 678030 112500 678270
rect 112740 678030 112830 678270
rect 113070 678030 113160 678270
rect 113400 678030 113490 678270
rect 113730 678030 113840 678270
rect 114080 678030 114170 678270
rect 114410 678030 114500 678270
rect 114740 678030 114830 678270
rect 115070 678030 115180 678270
rect 115420 678030 115510 678270
rect 115750 678030 115840 678270
rect 116080 678030 116170 678270
rect 116410 678030 116520 678270
rect 116760 678030 116850 678270
rect 117090 678030 117180 678270
rect 117420 678030 117510 678270
rect 117750 678030 117860 678270
rect 118100 678030 118190 678270
rect 118430 678030 118520 678270
rect 118760 678030 118850 678270
rect 119090 678030 119200 678270
rect 119440 678030 119530 678270
rect 119770 678030 119860 678270
rect 120100 678030 120190 678270
rect 120430 678030 120540 678270
rect 120780 678030 120870 678270
rect 121110 678030 121200 678270
rect 121440 678030 121530 678270
rect 121770 678030 122190 678270
rect 122430 678030 122540 678270
rect 122780 678030 122870 678270
rect 123110 678030 123200 678270
rect 123440 678030 123530 678270
rect 123770 678030 123880 678270
rect 124120 678030 124210 678270
rect 124450 678030 124540 678270
rect 124780 678030 124870 678270
rect 125110 678030 125220 678270
rect 125460 678030 125550 678270
rect 125790 678030 125880 678270
rect 126120 678030 126210 678270
rect 126450 678030 126560 678270
rect 126800 678030 126890 678270
rect 127130 678030 127220 678270
rect 127460 678030 127550 678270
rect 127790 678030 127900 678270
rect 128140 678030 128230 678270
rect 128470 678030 128560 678270
rect 128800 678030 128890 678270
rect 129130 678030 129240 678270
rect 129480 678030 129570 678270
rect 129810 678030 129900 678270
rect 130140 678030 130230 678270
rect 130470 678030 130580 678270
rect 130820 678030 130910 678270
rect 131150 678030 131240 678270
rect 131480 678030 131570 678270
rect 131810 678030 131920 678270
rect 132160 678030 132250 678270
rect 132490 678030 132580 678270
rect 132820 678030 132910 678270
rect 133150 678030 133570 678270
rect 133810 678030 133920 678270
rect 134160 678030 134250 678270
rect 134490 678030 134580 678270
rect 134820 678030 134910 678270
rect 135150 678030 135260 678270
rect 135500 678030 135590 678270
rect 135830 678030 135920 678270
rect 136160 678030 136250 678270
rect 136490 678030 136600 678270
rect 136840 678030 136930 678270
rect 137170 678030 137260 678270
rect 137500 678030 137590 678270
rect 137830 678030 137940 678270
rect 138180 678030 138270 678270
rect 138510 678030 138600 678270
rect 138840 678030 138930 678270
rect 139170 678030 139280 678270
rect 139520 678030 139610 678270
rect 139850 678030 139940 678270
rect 140180 678030 140270 678270
rect 140510 678030 140620 678270
rect 140860 678030 140950 678270
rect 141190 678030 141280 678270
rect 141520 678030 141610 678270
rect 141850 678030 141960 678270
rect 142200 678030 142290 678270
rect 142530 678030 142620 678270
rect 142860 678030 142950 678270
rect 143190 678030 143300 678270
rect 143540 678030 143630 678270
rect 143870 678030 143960 678270
rect 144200 678030 144290 678270
rect 144530 678030 144950 678270
rect 145190 678030 145300 678270
rect 145540 678030 145630 678270
rect 145870 678030 145960 678270
rect 146200 678030 146290 678270
rect 146530 678030 146640 678270
rect 146880 678030 146970 678270
rect 147210 678030 147300 678270
rect 147540 678030 147630 678270
rect 147870 678030 147980 678270
rect 148220 678030 148310 678270
rect 148550 678030 148640 678270
rect 148880 678030 148970 678270
rect 149210 678030 149320 678270
rect 149560 678030 149650 678270
rect 149890 678030 149980 678270
rect 150220 678030 150310 678270
rect 150550 678030 150660 678270
rect 150900 678030 150990 678270
rect 151230 678030 151320 678270
rect 151560 678030 151650 678270
rect 151890 678030 152000 678270
rect 152240 678030 152330 678270
rect 152570 678030 152660 678270
rect 152900 678030 152990 678270
rect 153230 678030 153340 678270
rect 153580 678030 153670 678270
rect 153910 678030 154000 678270
rect 154240 678030 154330 678270
rect 154570 678030 154680 678270
rect 154920 678030 155010 678270
rect 155250 678030 155340 678270
rect 155580 678030 155670 678270
rect 155910 678030 155960 678270
rect 110760 677920 155960 678030
rect 110760 677680 110810 677920
rect 111050 677680 111160 677920
rect 111400 677680 111490 677920
rect 111730 677680 111820 677920
rect 112060 677680 112150 677920
rect 112390 677680 112500 677920
rect 112740 677680 112830 677920
rect 113070 677680 113160 677920
rect 113400 677680 113490 677920
rect 113730 677680 113840 677920
rect 114080 677680 114170 677920
rect 114410 677680 114500 677920
rect 114740 677680 114830 677920
rect 115070 677680 115180 677920
rect 115420 677680 115510 677920
rect 115750 677680 115840 677920
rect 116080 677680 116170 677920
rect 116410 677680 116520 677920
rect 116760 677680 116850 677920
rect 117090 677680 117180 677920
rect 117420 677680 117510 677920
rect 117750 677680 117860 677920
rect 118100 677680 118190 677920
rect 118430 677680 118520 677920
rect 118760 677680 118850 677920
rect 119090 677680 119200 677920
rect 119440 677680 119530 677920
rect 119770 677680 119860 677920
rect 120100 677680 120190 677920
rect 120430 677680 120540 677920
rect 120780 677680 120870 677920
rect 121110 677680 121200 677920
rect 121440 677680 121530 677920
rect 121770 677680 122190 677920
rect 122430 677680 122540 677920
rect 122780 677680 122870 677920
rect 123110 677680 123200 677920
rect 123440 677680 123530 677920
rect 123770 677680 123880 677920
rect 124120 677680 124210 677920
rect 124450 677680 124540 677920
rect 124780 677680 124870 677920
rect 125110 677680 125220 677920
rect 125460 677680 125550 677920
rect 125790 677680 125880 677920
rect 126120 677680 126210 677920
rect 126450 677680 126560 677920
rect 126800 677680 126890 677920
rect 127130 677680 127220 677920
rect 127460 677680 127550 677920
rect 127790 677680 127900 677920
rect 128140 677680 128230 677920
rect 128470 677680 128560 677920
rect 128800 677680 128890 677920
rect 129130 677680 129240 677920
rect 129480 677680 129570 677920
rect 129810 677680 129900 677920
rect 130140 677680 130230 677920
rect 130470 677680 130580 677920
rect 130820 677680 130910 677920
rect 131150 677680 131240 677920
rect 131480 677680 131570 677920
rect 131810 677680 131920 677920
rect 132160 677680 132250 677920
rect 132490 677680 132580 677920
rect 132820 677680 132910 677920
rect 133150 677680 133570 677920
rect 133810 677680 133920 677920
rect 134160 677680 134250 677920
rect 134490 677680 134580 677920
rect 134820 677680 134910 677920
rect 135150 677680 135260 677920
rect 135500 677680 135590 677920
rect 135830 677680 135920 677920
rect 136160 677680 136250 677920
rect 136490 677680 136600 677920
rect 136840 677680 136930 677920
rect 137170 677680 137260 677920
rect 137500 677680 137590 677920
rect 137830 677680 137940 677920
rect 138180 677680 138270 677920
rect 138510 677680 138600 677920
rect 138840 677680 138930 677920
rect 139170 677680 139280 677920
rect 139520 677680 139610 677920
rect 139850 677680 139940 677920
rect 140180 677680 140270 677920
rect 140510 677680 140620 677920
rect 140860 677680 140950 677920
rect 141190 677680 141280 677920
rect 141520 677680 141610 677920
rect 141850 677680 141960 677920
rect 142200 677680 142290 677920
rect 142530 677680 142620 677920
rect 142860 677680 142950 677920
rect 143190 677680 143300 677920
rect 143540 677680 143630 677920
rect 143870 677680 143960 677920
rect 144200 677680 144290 677920
rect 144530 677680 144950 677920
rect 145190 677680 145300 677920
rect 145540 677680 145630 677920
rect 145870 677680 145960 677920
rect 146200 677680 146290 677920
rect 146530 677680 146640 677920
rect 146880 677680 146970 677920
rect 147210 677680 147300 677920
rect 147540 677680 147630 677920
rect 147870 677680 147980 677920
rect 148220 677680 148310 677920
rect 148550 677680 148640 677920
rect 148880 677680 148970 677920
rect 149210 677680 149320 677920
rect 149560 677680 149650 677920
rect 149890 677680 149980 677920
rect 150220 677680 150310 677920
rect 150550 677680 150660 677920
rect 150900 677680 150990 677920
rect 151230 677680 151320 677920
rect 151560 677680 151650 677920
rect 151890 677680 152000 677920
rect 152240 677680 152330 677920
rect 152570 677680 152660 677920
rect 152900 677680 152990 677920
rect 153230 677680 153340 677920
rect 153580 677680 153670 677920
rect 153910 677680 154000 677920
rect 154240 677680 154330 677920
rect 154570 677680 154680 677920
rect 154920 677680 155010 677920
rect 155250 677680 155340 677920
rect 155580 677680 155670 677920
rect 155910 677680 155960 677920
rect 110760 677590 155960 677680
rect 110760 677350 110810 677590
rect 111050 677350 111160 677590
rect 111400 677350 111490 677590
rect 111730 677350 111820 677590
rect 112060 677350 112150 677590
rect 112390 677350 112500 677590
rect 112740 677350 112830 677590
rect 113070 677350 113160 677590
rect 113400 677350 113490 677590
rect 113730 677350 113840 677590
rect 114080 677350 114170 677590
rect 114410 677350 114500 677590
rect 114740 677350 114830 677590
rect 115070 677350 115180 677590
rect 115420 677350 115510 677590
rect 115750 677350 115840 677590
rect 116080 677350 116170 677590
rect 116410 677350 116520 677590
rect 116760 677350 116850 677590
rect 117090 677350 117180 677590
rect 117420 677350 117510 677590
rect 117750 677350 117860 677590
rect 118100 677350 118190 677590
rect 118430 677350 118520 677590
rect 118760 677350 118850 677590
rect 119090 677350 119200 677590
rect 119440 677350 119530 677590
rect 119770 677350 119860 677590
rect 120100 677350 120190 677590
rect 120430 677350 120540 677590
rect 120780 677350 120870 677590
rect 121110 677350 121200 677590
rect 121440 677350 121530 677590
rect 121770 677350 122190 677590
rect 122430 677350 122540 677590
rect 122780 677350 122870 677590
rect 123110 677350 123200 677590
rect 123440 677350 123530 677590
rect 123770 677350 123880 677590
rect 124120 677350 124210 677590
rect 124450 677350 124540 677590
rect 124780 677350 124870 677590
rect 125110 677350 125220 677590
rect 125460 677350 125550 677590
rect 125790 677350 125880 677590
rect 126120 677350 126210 677590
rect 126450 677350 126560 677590
rect 126800 677350 126890 677590
rect 127130 677350 127220 677590
rect 127460 677350 127550 677590
rect 127790 677350 127900 677590
rect 128140 677350 128230 677590
rect 128470 677350 128560 677590
rect 128800 677350 128890 677590
rect 129130 677350 129240 677590
rect 129480 677350 129570 677590
rect 129810 677350 129900 677590
rect 130140 677350 130230 677590
rect 130470 677350 130580 677590
rect 130820 677350 130910 677590
rect 131150 677350 131240 677590
rect 131480 677350 131570 677590
rect 131810 677350 131920 677590
rect 132160 677350 132250 677590
rect 132490 677350 132580 677590
rect 132820 677350 132910 677590
rect 133150 677350 133570 677590
rect 133810 677350 133920 677590
rect 134160 677350 134250 677590
rect 134490 677350 134580 677590
rect 134820 677350 134910 677590
rect 135150 677350 135260 677590
rect 135500 677350 135590 677590
rect 135830 677350 135920 677590
rect 136160 677350 136250 677590
rect 136490 677350 136600 677590
rect 136840 677350 136930 677590
rect 137170 677350 137260 677590
rect 137500 677350 137590 677590
rect 137830 677350 137940 677590
rect 138180 677350 138270 677590
rect 138510 677350 138600 677590
rect 138840 677350 138930 677590
rect 139170 677350 139280 677590
rect 139520 677350 139610 677590
rect 139850 677350 139940 677590
rect 140180 677350 140270 677590
rect 140510 677350 140620 677590
rect 140860 677350 140950 677590
rect 141190 677350 141280 677590
rect 141520 677350 141610 677590
rect 141850 677350 141960 677590
rect 142200 677350 142290 677590
rect 142530 677350 142620 677590
rect 142860 677350 142950 677590
rect 143190 677350 143300 677590
rect 143540 677350 143630 677590
rect 143870 677350 143960 677590
rect 144200 677350 144290 677590
rect 144530 677350 144950 677590
rect 145190 677350 145300 677590
rect 145540 677350 145630 677590
rect 145870 677350 145960 677590
rect 146200 677350 146290 677590
rect 146530 677350 146640 677590
rect 146880 677350 146970 677590
rect 147210 677350 147300 677590
rect 147540 677350 147630 677590
rect 147870 677350 147980 677590
rect 148220 677350 148310 677590
rect 148550 677350 148640 677590
rect 148880 677350 148970 677590
rect 149210 677350 149320 677590
rect 149560 677350 149650 677590
rect 149890 677350 149980 677590
rect 150220 677350 150310 677590
rect 150550 677350 150660 677590
rect 150900 677350 150990 677590
rect 151230 677350 151320 677590
rect 151560 677350 151650 677590
rect 151890 677350 152000 677590
rect 152240 677350 152330 677590
rect 152570 677350 152660 677590
rect 152900 677350 152990 677590
rect 153230 677350 153340 677590
rect 153580 677350 153670 677590
rect 153910 677350 154000 677590
rect 154240 677350 154330 677590
rect 154570 677350 154680 677590
rect 154920 677350 155010 677590
rect 155250 677350 155340 677590
rect 155580 677350 155670 677590
rect 155910 677350 155960 677590
rect 110760 677260 155960 677350
rect 110760 677020 110810 677260
rect 111050 677020 111160 677260
rect 111400 677020 111490 677260
rect 111730 677020 111820 677260
rect 112060 677020 112150 677260
rect 112390 677020 112500 677260
rect 112740 677020 112830 677260
rect 113070 677020 113160 677260
rect 113400 677020 113490 677260
rect 113730 677020 113840 677260
rect 114080 677020 114170 677260
rect 114410 677020 114500 677260
rect 114740 677020 114830 677260
rect 115070 677020 115180 677260
rect 115420 677020 115510 677260
rect 115750 677020 115840 677260
rect 116080 677020 116170 677260
rect 116410 677020 116520 677260
rect 116760 677020 116850 677260
rect 117090 677020 117180 677260
rect 117420 677020 117510 677260
rect 117750 677020 117860 677260
rect 118100 677020 118190 677260
rect 118430 677020 118520 677260
rect 118760 677020 118850 677260
rect 119090 677020 119200 677260
rect 119440 677020 119530 677260
rect 119770 677020 119860 677260
rect 120100 677020 120190 677260
rect 120430 677020 120540 677260
rect 120780 677020 120870 677260
rect 121110 677020 121200 677260
rect 121440 677020 121530 677260
rect 121770 677020 122190 677260
rect 122430 677020 122540 677260
rect 122780 677020 122870 677260
rect 123110 677020 123200 677260
rect 123440 677020 123530 677260
rect 123770 677020 123880 677260
rect 124120 677020 124210 677260
rect 124450 677020 124540 677260
rect 124780 677020 124870 677260
rect 125110 677020 125220 677260
rect 125460 677020 125550 677260
rect 125790 677020 125880 677260
rect 126120 677020 126210 677260
rect 126450 677020 126560 677260
rect 126800 677020 126890 677260
rect 127130 677020 127220 677260
rect 127460 677020 127550 677260
rect 127790 677020 127900 677260
rect 128140 677020 128230 677260
rect 128470 677020 128560 677260
rect 128800 677020 128890 677260
rect 129130 677020 129240 677260
rect 129480 677020 129570 677260
rect 129810 677020 129900 677260
rect 130140 677020 130230 677260
rect 130470 677020 130580 677260
rect 130820 677020 130910 677260
rect 131150 677020 131240 677260
rect 131480 677020 131570 677260
rect 131810 677020 131920 677260
rect 132160 677020 132250 677260
rect 132490 677020 132580 677260
rect 132820 677020 132910 677260
rect 133150 677020 133570 677260
rect 133810 677020 133920 677260
rect 134160 677020 134250 677260
rect 134490 677020 134580 677260
rect 134820 677020 134910 677260
rect 135150 677020 135260 677260
rect 135500 677020 135590 677260
rect 135830 677020 135920 677260
rect 136160 677020 136250 677260
rect 136490 677020 136600 677260
rect 136840 677020 136930 677260
rect 137170 677020 137260 677260
rect 137500 677020 137590 677260
rect 137830 677020 137940 677260
rect 138180 677020 138270 677260
rect 138510 677020 138600 677260
rect 138840 677020 138930 677260
rect 139170 677020 139280 677260
rect 139520 677020 139610 677260
rect 139850 677020 139940 677260
rect 140180 677020 140270 677260
rect 140510 677020 140620 677260
rect 140860 677020 140950 677260
rect 141190 677020 141280 677260
rect 141520 677020 141610 677260
rect 141850 677020 141960 677260
rect 142200 677020 142290 677260
rect 142530 677020 142620 677260
rect 142860 677020 142950 677260
rect 143190 677020 143300 677260
rect 143540 677020 143630 677260
rect 143870 677020 143960 677260
rect 144200 677020 144290 677260
rect 144530 677020 144950 677260
rect 145190 677020 145300 677260
rect 145540 677020 145630 677260
rect 145870 677020 145960 677260
rect 146200 677020 146290 677260
rect 146530 677020 146640 677260
rect 146880 677020 146970 677260
rect 147210 677020 147300 677260
rect 147540 677020 147630 677260
rect 147870 677020 147980 677260
rect 148220 677020 148310 677260
rect 148550 677020 148640 677260
rect 148880 677020 148970 677260
rect 149210 677020 149320 677260
rect 149560 677020 149650 677260
rect 149890 677020 149980 677260
rect 150220 677020 150310 677260
rect 150550 677020 150660 677260
rect 150900 677020 150990 677260
rect 151230 677020 151320 677260
rect 151560 677020 151650 677260
rect 151890 677020 152000 677260
rect 152240 677020 152330 677260
rect 152570 677020 152660 677260
rect 152900 677020 152990 677260
rect 153230 677020 153340 677260
rect 153580 677020 153670 677260
rect 153910 677020 154000 677260
rect 154240 677020 154330 677260
rect 154570 677020 154680 677260
rect 154920 677020 155010 677260
rect 155250 677020 155340 677260
rect 155580 677020 155670 677260
rect 155910 677020 155960 677260
rect 110760 676930 155960 677020
rect 110760 676690 110810 676930
rect 111050 676690 111160 676930
rect 111400 676690 111490 676930
rect 111730 676690 111820 676930
rect 112060 676690 112150 676930
rect 112390 676690 112500 676930
rect 112740 676690 112830 676930
rect 113070 676690 113160 676930
rect 113400 676690 113490 676930
rect 113730 676690 113840 676930
rect 114080 676690 114170 676930
rect 114410 676690 114500 676930
rect 114740 676690 114830 676930
rect 115070 676690 115180 676930
rect 115420 676690 115510 676930
rect 115750 676690 115840 676930
rect 116080 676690 116170 676930
rect 116410 676690 116520 676930
rect 116760 676690 116850 676930
rect 117090 676690 117180 676930
rect 117420 676690 117510 676930
rect 117750 676690 117860 676930
rect 118100 676690 118190 676930
rect 118430 676690 118520 676930
rect 118760 676690 118850 676930
rect 119090 676690 119200 676930
rect 119440 676690 119530 676930
rect 119770 676690 119860 676930
rect 120100 676690 120190 676930
rect 120430 676690 120540 676930
rect 120780 676690 120870 676930
rect 121110 676690 121200 676930
rect 121440 676690 121530 676930
rect 121770 676690 122190 676930
rect 122430 676690 122540 676930
rect 122780 676690 122870 676930
rect 123110 676690 123200 676930
rect 123440 676690 123530 676930
rect 123770 676690 123880 676930
rect 124120 676690 124210 676930
rect 124450 676690 124540 676930
rect 124780 676690 124870 676930
rect 125110 676690 125220 676930
rect 125460 676690 125550 676930
rect 125790 676690 125880 676930
rect 126120 676690 126210 676930
rect 126450 676690 126560 676930
rect 126800 676690 126890 676930
rect 127130 676690 127220 676930
rect 127460 676690 127550 676930
rect 127790 676690 127900 676930
rect 128140 676690 128230 676930
rect 128470 676690 128560 676930
rect 128800 676690 128890 676930
rect 129130 676690 129240 676930
rect 129480 676690 129570 676930
rect 129810 676690 129900 676930
rect 130140 676690 130230 676930
rect 130470 676690 130580 676930
rect 130820 676690 130910 676930
rect 131150 676690 131240 676930
rect 131480 676690 131570 676930
rect 131810 676690 131920 676930
rect 132160 676690 132250 676930
rect 132490 676690 132580 676930
rect 132820 676690 132910 676930
rect 133150 676690 133570 676930
rect 133810 676690 133920 676930
rect 134160 676690 134250 676930
rect 134490 676690 134580 676930
rect 134820 676690 134910 676930
rect 135150 676690 135260 676930
rect 135500 676690 135590 676930
rect 135830 676690 135920 676930
rect 136160 676690 136250 676930
rect 136490 676690 136600 676930
rect 136840 676690 136930 676930
rect 137170 676690 137260 676930
rect 137500 676690 137590 676930
rect 137830 676690 137940 676930
rect 138180 676690 138270 676930
rect 138510 676690 138600 676930
rect 138840 676690 138930 676930
rect 139170 676690 139280 676930
rect 139520 676690 139610 676930
rect 139850 676690 139940 676930
rect 140180 676690 140270 676930
rect 140510 676690 140620 676930
rect 140860 676690 140950 676930
rect 141190 676690 141280 676930
rect 141520 676690 141610 676930
rect 141850 676690 141960 676930
rect 142200 676690 142290 676930
rect 142530 676690 142620 676930
rect 142860 676690 142950 676930
rect 143190 676690 143300 676930
rect 143540 676690 143630 676930
rect 143870 676690 143960 676930
rect 144200 676690 144290 676930
rect 144530 676690 144950 676930
rect 145190 676690 145300 676930
rect 145540 676690 145630 676930
rect 145870 676690 145960 676930
rect 146200 676690 146290 676930
rect 146530 676690 146640 676930
rect 146880 676690 146970 676930
rect 147210 676690 147300 676930
rect 147540 676690 147630 676930
rect 147870 676690 147980 676930
rect 148220 676690 148310 676930
rect 148550 676690 148640 676930
rect 148880 676690 148970 676930
rect 149210 676690 149320 676930
rect 149560 676690 149650 676930
rect 149890 676690 149980 676930
rect 150220 676690 150310 676930
rect 150550 676690 150660 676930
rect 150900 676690 150990 676930
rect 151230 676690 151320 676930
rect 151560 676690 151650 676930
rect 151890 676690 152000 676930
rect 152240 676690 152330 676930
rect 152570 676690 152660 676930
rect 152900 676690 152990 676930
rect 153230 676690 153340 676930
rect 153580 676690 153670 676930
rect 153910 676690 154000 676930
rect 154240 676690 154330 676930
rect 154570 676690 154680 676930
rect 154920 676690 155010 676930
rect 155250 676690 155340 676930
rect 155580 676690 155670 676930
rect 155910 676690 155960 676930
rect 110760 676580 155960 676690
rect 110760 676340 110810 676580
rect 111050 676340 111160 676580
rect 111400 676340 111490 676580
rect 111730 676340 111820 676580
rect 112060 676340 112150 676580
rect 112390 676340 112500 676580
rect 112740 676340 112830 676580
rect 113070 676340 113160 676580
rect 113400 676340 113490 676580
rect 113730 676340 113840 676580
rect 114080 676340 114170 676580
rect 114410 676340 114500 676580
rect 114740 676340 114830 676580
rect 115070 676340 115180 676580
rect 115420 676340 115510 676580
rect 115750 676340 115840 676580
rect 116080 676340 116170 676580
rect 116410 676340 116520 676580
rect 116760 676340 116850 676580
rect 117090 676340 117180 676580
rect 117420 676340 117510 676580
rect 117750 676340 117860 676580
rect 118100 676340 118190 676580
rect 118430 676340 118520 676580
rect 118760 676340 118850 676580
rect 119090 676340 119200 676580
rect 119440 676340 119530 676580
rect 119770 676340 119860 676580
rect 120100 676340 120190 676580
rect 120430 676340 120540 676580
rect 120780 676340 120870 676580
rect 121110 676340 121200 676580
rect 121440 676340 121530 676580
rect 121770 676340 122190 676580
rect 122430 676340 122540 676580
rect 122780 676340 122870 676580
rect 123110 676340 123200 676580
rect 123440 676340 123530 676580
rect 123770 676340 123880 676580
rect 124120 676340 124210 676580
rect 124450 676340 124540 676580
rect 124780 676340 124870 676580
rect 125110 676340 125220 676580
rect 125460 676340 125550 676580
rect 125790 676340 125880 676580
rect 126120 676340 126210 676580
rect 126450 676340 126560 676580
rect 126800 676340 126890 676580
rect 127130 676340 127220 676580
rect 127460 676340 127550 676580
rect 127790 676340 127900 676580
rect 128140 676340 128230 676580
rect 128470 676340 128560 676580
rect 128800 676340 128890 676580
rect 129130 676340 129240 676580
rect 129480 676340 129570 676580
rect 129810 676340 129900 676580
rect 130140 676340 130230 676580
rect 130470 676340 130580 676580
rect 130820 676340 130910 676580
rect 131150 676340 131240 676580
rect 131480 676340 131570 676580
rect 131810 676340 131920 676580
rect 132160 676340 132250 676580
rect 132490 676340 132580 676580
rect 132820 676340 132910 676580
rect 133150 676340 133570 676580
rect 133810 676340 133920 676580
rect 134160 676340 134250 676580
rect 134490 676340 134580 676580
rect 134820 676340 134910 676580
rect 135150 676340 135260 676580
rect 135500 676340 135590 676580
rect 135830 676340 135920 676580
rect 136160 676340 136250 676580
rect 136490 676340 136600 676580
rect 136840 676340 136930 676580
rect 137170 676340 137260 676580
rect 137500 676340 137590 676580
rect 137830 676340 137940 676580
rect 138180 676340 138270 676580
rect 138510 676340 138600 676580
rect 138840 676340 138930 676580
rect 139170 676340 139280 676580
rect 139520 676340 139610 676580
rect 139850 676340 139940 676580
rect 140180 676340 140270 676580
rect 140510 676340 140620 676580
rect 140860 676340 140950 676580
rect 141190 676340 141280 676580
rect 141520 676340 141610 676580
rect 141850 676340 141960 676580
rect 142200 676340 142290 676580
rect 142530 676340 142620 676580
rect 142860 676340 142950 676580
rect 143190 676340 143300 676580
rect 143540 676340 143630 676580
rect 143870 676340 143960 676580
rect 144200 676340 144290 676580
rect 144530 676340 144950 676580
rect 145190 676340 145300 676580
rect 145540 676340 145630 676580
rect 145870 676340 145960 676580
rect 146200 676340 146290 676580
rect 146530 676340 146640 676580
rect 146880 676340 146970 676580
rect 147210 676340 147300 676580
rect 147540 676340 147630 676580
rect 147870 676340 147980 676580
rect 148220 676340 148310 676580
rect 148550 676340 148640 676580
rect 148880 676340 148970 676580
rect 149210 676340 149320 676580
rect 149560 676340 149650 676580
rect 149890 676340 149980 676580
rect 150220 676340 150310 676580
rect 150550 676340 150660 676580
rect 150900 676340 150990 676580
rect 151230 676340 151320 676580
rect 151560 676340 151650 676580
rect 151890 676340 152000 676580
rect 152240 676340 152330 676580
rect 152570 676340 152660 676580
rect 152900 676340 152990 676580
rect 153230 676340 153340 676580
rect 153580 676340 153670 676580
rect 153910 676340 154000 676580
rect 154240 676340 154330 676580
rect 154570 676340 154680 676580
rect 154920 676340 155010 676580
rect 155250 676340 155340 676580
rect 155580 676340 155670 676580
rect 155910 676340 155960 676580
rect 110760 676250 155960 676340
rect 110760 676010 110810 676250
rect 111050 676010 111160 676250
rect 111400 676010 111490 676250
rect 111730 676010 111820 676250
rect 112060 676010 112150 676250
rect 112390 676010 112500 676250
rect 112740 676010 112830 676250
rect 113070 676010 113160 676250
rect 113400 676010 113490 676250
rect 113730 676010 113840 676250
rect 114080 676010 114170 676250
rect 114410 676010 114500 676250
rect 114740 676010 114830 676250
rect 115070 676010 115180 676250
rect 115420 676010 115510 676250
rect 115750 676010 115840 676250
rect 116080 676010 116170 676250
rect 116410 676010 116520 676250
rect 116760 676010 116850 676250
rect 117090 676010 117180 676250
rect 117420 676010 117510 676250
rect 117750 676010 117860 676250
rect 118100 676010 118190 676250
rect 118430 676010 118520 676250
rect 118760 676010 118850 676250
rect 119090 676010 119200 676250
rect 119440 676010 119530 676250
rect 119770 676010 119860 676250
rect 120100 676010 120190 676250
rect 120430 676010 120540 676250
rect 120780 676010 120870 676250
rect 121110 676010 121200 676250
rect 121440 676010 121530 676250
rect 121770 676010 122190 676250
rect 122430 676010 122540 676250
rect 122780 676010 122870 676250
rect 123110 676010 123200 676250
rect 123440 676010 123530 676250
rect 123770 676010 123880 676250
rect 124120 676010 124210 676250
rect 124450 676010 124540 676250
rect 124780 676010 124870 676250
rect 125110 676010 125220 676250
rect 125460 676010 125550 676250
rect 125790 676010 125880 676250
rect 126120 676010 126210 676250
rect 126450 676010 126560 676250
rect 126800 676010 126890 676250
rect 127130 676010 127220 676250
rect 127460 676010 127550 676250
rect 127790 676010 127900 676250
rect 128140 676010 128230 676250
rect 128470 676010 128560 676250
rect 128800 676010 128890 676250
rect 129130 676010 129240 676250
rect 129480 676010 129570 676250
rect 129810 676010 129900 676250
rect 130140 676010 130230 676250
rect 130470 676010 130580 676250
rect 130820 676010 130910 676250
rect 131150 676010 131240 676250
rect 131480 676010 131570 676250
rect 131810 676010 131920 676250
rect 132160 676010 132250 676250
rect 132490 676010 132580 676250
rect 132820 676010 132910 676250
rect 133150 676010 133570 676250
rect 133810 676010 133920 676250
rect 134160 676010 134250 676250
rect 134490 676010 134580 676250
rect 134820 676010 134910 676250
rect 135150 676010 135260 676250
rect 135500 676010 135590 676250
rect 135830 676010 135920 676250
rect 136160 676010 136250 676250
rect 136490 676010 136600 676250
rect 136840 676010 136930 676250
rect 137170 676010 137260 676250
rect 137500 676010 137590 676250
rect 137830 676010 137940 676250
rect 138180 676010 138270 676250
rect 138510 676010 138600 676250
rect 138840 676010 138930 676250
rect 139170 676010 139280 676250
rect 139520 676010 139610 676250
rect 139850 676010 139940 676250
rect 140180 676010 140270 676250
rect 140510 676010 140620 676250
rect 140860 676010 140950 676250
rect 141190 676010 141280 676250
rect 141520 676010 141610 676250
rect 141850 676010 141960 676250
rect 142200 676010 142290 676250
rect 142530 676010 142620 676250
rect 142860 676010 142950 676250
rect 143190 676010 143300 676250
rect 143540 676010 143630 676250
rect 143870 676010 143960 676250
rect 144200 676010 144290 676250
rect 144530 676010 144950 676250
rect 145190 676010 145300 676250
rect 145540 676010 145630 676250
rect 145870 676010 145960 676250
rect 146200 676010 146290 676250
rect 146530 676010 146640 676250
rect 146880 676010 146970 676250
rect 147210 676010 147300 676250
rect 147540 676010 147630 676250
rect 147870 676010 147980 676250
rect 148220 676010 148310 676250
rect 148550 676010 148640 676250
rect 148880 676010 148970 676250
rect 149210 676010 149320 676250
rect 149560 676010 149650 676250
rect 149890 676010 149980 676250
rect 150220 676010 150310 676250
rect 150550 676010 150660 676250
rect 150900 676010 150990 676250
rect 151230 676010 151320 676250
rect 151560 676010 151650 676250
rect 151890 676010 152000 676250
rect 152240 676010 152330 676250
rect 152570 676010 152660 676250
rect 152900 676010 152990 676250
rect 153230 676010 153340 676250
rect 153580 676010 153670 676250
rect 153910 676010 154000 676250
rect 154240 676010 154330 676250
rect 154570 676010 154680 676250
rect 154920 676010 155010 676250
rect 155250 676010 155340 676250
rect 155580 676010 155670 676250
rect 155910 676010 155960 676250
rect 110760 675920 155960 676010
rect 110760 675680 110810 675920
rect 111050 675680 111160 675920
rect 111400 675680 111490 675920
rect 111730 675680 111820 675920
rect 112060 675680 112150 675920
rect 112390 675680 112500 675920
rect 112740 675680 112830 675920
rect 113070 675680 113160 675920
rect 113400 675680 113490 675920
rect 113730 675680 113840 675920
rect 114080 675680 114170 675920
rect 114410 675680 114500 675920
rect 114740 675680 114830 675920
rect 115070 675680 115180 675920
rect 115420 675680 115510 675920
rect 115750 675680 115840 675920
rect 116080 675680 116170 675920
rect 116410 675680 116520 675920
rect 116760 675680 116850 675920
rect 117090 675680 117180 675920
rect 117420 675680 117510 675920
rect 117750 675680 117860 675920
rect 118100 675680 118190 675920
rect 118430 675680 118520 675920
rect 118760 675680 118850 675920
rect 119090 675680 119200 675920
rect 119440 675680 119530 675920
rect 119770 675680 119860 675920
rect 120100 675680 120190 675920
rect 120430 675680 120540 675920
rect 120780 675680 120870 675920
rect 121110 675680 121200 675920
rect 121440 675680 121530 675920
rect 121770 675680 122190 675920
rect 122430 675680 122540 675920
rect 122780 675680 122870 675920
rect 123110 675680 123200 675920
rect 123440 675680 123530 675920
rect 123770 675680 123880 675920
rect 124120 675680 124210 675920
rect 124450 675680 124540 675920
rect 124780 675680 124870 675920
rect 125110 675680 125220 675920
rect 125460 675680 125550 675920
rect 125790 675680 125880 675920
rect 126120 675680 126210 675920
rect 126450 675680 126560 675920
rect 126800 675680 126890 675920
rect 127130 675680 127220 675920
rect 127460 675680 127550 675920
rect 127790 675680 127900 675920
rect 128140 675680 128230 675920
rect 128470 675680 128560 675920
rect 128800 675680 128890 675920
rect 129130 675680 129240 675920
rect 129480 675680 129570 675920
rect 129810 675680 129900 675920
rect 130140 675680 130230 675920
rect 130470 675680 130580 675920
rect 130820 675680 130910 675920
rect 131150 675680 131240 675920
rect 131480 675680 131570 675920
rect 131810 675680 131920 675920
rect 132160 675680 132250 675920
rect 132490 675680 132580 675920
rect 132820 675680 132910 675920
rect 133150 675680 133570 675920
rect 133810 675680 133920 675920
rect 134160 675680 134250 675920
rect 134490 675680 134580 675920
rect 134820 675680 134910 675920
rect 135150 675680 135260 675920
rect 135500 675680 135590 675920
rect 135830 675680 135920 675920
rect 136160 675680 136250 675920
rect 136490 675680 136600 675920
rect 136840 675680 136930 675920
rect 137170 675680 137260 675920
rect 137500 675680 137590 675920
rect 137830 675680 137940 675920
rect 138180 675680 138270 675920
rect 138510 675680 138600 675920
rect 138840 675680 138930 675920
rect 139170 675680 139280 675920
rect 139520 675680 139610 675920
rect 139850 675680 139940 675920
rect 140180 675680 140270 675920
rect 140510 675680 140620 675920
rect 140860 675680 140950 675920
rect 141190 675680 141280 675920
rect 141520 675680 141610 675920
rect 141850 675680 141960 675920
rect 142200 675680 142290 675920
rect 142530 675680 142620 675920
rect 142860 675680 142950 675920
rect 143190 675680 143300 675920
rect 143540 675680 143630 675920
rect 143870 675680 143960 675920
rect 144200 675680 144290 675920
rect 144530 675680 144950 675920
rect 145190 675680 145300 675920
rect 145540 675680 145630 675920
rect 145870 675680 145960 675920
rect 146200 675680 146290 675920
rect 146530 675680 146640 675920
rect 146880 675680 146970 675920
rect 147210 675680 147300 675920
rect 147540 675680 147630 675920
rect 147870 675680 147980 675920
rect 148220 675680 148310 675920
rect 148550 675680 148640 675920
rect 148880 675680 148970 675920
rect 149210 675680 149320 675920
rect 149560 675680 149650 675920
rect 149890 675680 149980 675920
rect 150220 675680 150310 675920
rect 150550 675680 150660 675920
rect 150900 675680 150990 675920
rect 151230 675680 151320 675920
rect 151560 675680 151650 675920
rect 151890 675680 152000 675920
rect 152240 675680 152330 675920
rect 152570 675680 152660 675920
rect 152900 675680 152990 675920
rect 153230 675680 153340 675920
rect 153580 675680 153670 675920
rect 153910 675680 154000 675920
rect 154240 675680 154330 675920
rect 154570 675680 154680 675920
rect 154920 675680 155010 675920
rect 155250 675680 155340 675920
rect 155580 675680 155670 675920
rect 155910 675680 155960 675920
rect 110760 675590 155960 675680
rect 110760 675350 110810 675590
rect 111050 675350 111160 675590
rect 111400 675350 111490 675590
rect 111730 675350 111820 675590
rect 112060 675350 112150 675590
rect 112390 675350 112500 675590
rect 112740 675350 112830 675590
rect 113070 675350 113160 675590
rect 113400 675350 113490 675590
rect 113730 675350 113840 675590
rect 114080 675350 114170 675590
rect 114410 675350 114500 675590
rect 114740 675350 114830 675590
rect 115070 675350 115180 675590
rect 115420 675350 115510 675590
rect 115750 675350 115840 675590
rect 116080 675350 116170 675590
rect 116410 675350 116520 675590
rect 116760 675350 116850 675590
rect 117090 675350 117180 675590
rect 117420 675350 117510 675590
rect 117750 675350 117860 675590
rect 118100 675350 118190 675590
rect 118430 675350 118520 675590
rect 118760 675350 118850 675590
rect 119090 675350 119200 675590
rect 119440 675350 119530 675590
rect 119770 675350 119860 675590
rect 120100 675350 120190 675590
rect 120430 675350 120540 675590
rect 120780 675350 120870 675590
rect 121110 675350 121200 675590
rect 121440 675350 121530 675590
rect 121770 675350 122190 675590
rect 122430 675350 122540 675590
rect 122780 675350 122870 675590
rect 123110 675350 123200 675590
rect 123440 675350 123530 675590
rect 123770 675350 123880 675590
rect 124120 675350 124210 675590
rect 124450 675350 124540 675590
rect 124780 675350 124870 675590
rect 125110 675350 125220 675590
rect 125460 675350 125550 675590
rect 125790 675350 125880 675590
rect 126120 675350 126210 675590
rect 126450 675350 126560 675590
rect 126800 675350 126890 675590
rect 127130 675350 127220 675590
rect 127460 675350 127550 675590
rect 127790 675350 127900 675590
rect 128140 675350 128230 675590
rect 128470 675350 128560 675590
rect 128800 675350 128890 675590
rect 129130 675350 129240 675590
rect 129480 675350 129570 675590
rect 129810 675350 129900 675590
rect 130140 675350 130230 675590
rect 130470 675350 130580 675590
rect 130820 675350 130910 675590
rect 131150 675350 131240 675590
rect 131480 675350 131570 675590
rect 131810 675350 131920 675590
rect 132160 675350 132250 675590
rect 132490 675350 132580 675590
rect 132820 675350 132910 675590
rect 133150 675350 133570 675590
rect 133810 675350 133920 675590
rect 134160 675350 134250 675590
rect 134490 675350 134580 675590
rect 134820 675350 134910 675590
rect 135150 675350 135260 675590
rect 135500 675350 135590 675590
rect 135830 675350 135920 675590
rect 136160 675350 136250 675590
rect 136490 675350 136600 675590
rect 136840 675350 136930 675590
rect 137170 675350 137260 675590
rect 137500 675350 137590 675590
rect 137830 675350 137940 675590
rect 138180 675350 138270 675590
rect 138510 675350 138600 675590
rect 138840 675350 138930 675590
rect 139170 675350 139280 675590
rect 139520 675350 139610 675590
rect 139850 675350 139940 675590
rect 140180 675350 140270 675590
rect 140510 675350 140620 675590
rect 140860 675350 140950 675590
rect 141190 675350 141280 675590
rect 141520 675350 141610 675590
rect 141850 675350 141960 675590
rect 142200 675350 142290 675590
rect 142530 675350 142620 675590
rect 142860 675350 142950 675590
rect 143190 675350 143300 675590
rect 143540 675350 143630 675590
rect 143870 675350 143960 675590
rect 144200 675350 144290 675590
rect 144530 675350 144950 675590
rect 145190 675350 145300 675590
rect 145540 675350 145630 675590
rect 145870 675350 145960 675590
rect 146200 675350 146290 675590
rect 146530 675350 146640 675590
rect 146880 675350 146970 675590
rect 147210 675350 147300 675590
rect 147540 675350 147630 675590
rect 147870 675350 147980 675590
rect 148220 675350 148310 675590
rect 148550 675350 148640 675590
rect 148880 675350 148970 675590
rect 149210 675350 149320 675590
rect 149560 675350 149650 675590
rect 149890 675350 149980 675590
rect 150220 675350 150310 675590
rect 150550 675350 150660 675590
rect 150900 675350 150990 675590
rect 151230 675350 151320 675590
rect 151560 675350 151650 675590
rect 151890 675350 152000 675590
rect 152240 675350 152330 675590
rect 152570 675350 152660 675590
rect 152900 675350 152990 675590
rect 153230 675350 153340 675590
rect 153580 675350 153670 675590
rect 153910 675350 154000 675590
rect 154240 675350 154330 675590
rect 154570 675350 154680 675590
rect 154920 675350 155010 675590
rect 155250 675350 155340 675590
rect 155580 675350 155670 675590
rect 155910 675350 155960 675590
rect 110760 675240 155960 675350
rect 110760 675000 110810 675240
rect 111050 675000 111160 675240
rect 111400 675000 111490 675240
rect 111730 675000 111820 675240
rect 112060 675000 112150 675240
rect 112390 675000 112500 675240
rect 112740 675000 112830 675240
rect 113070 675000 113160 675240
rect 113400 675000 113490 675240
rect 113730 675000 113840 675240
rect 114080 675000 114170 675240
rect 114410 675000 114500 675240
rect 114740 675000 114830 675240
rect 115070 675000 115180 675240
rect 115420 675000 115510 675240
rect 115750 675000 115840 675240
rect 116080 675000 116170 675240
rect 116410 675000 116520 675240
rect 116760 675000 116850 675240
rect 117090 675000 117180 675240
rect 117420 675000 117510 675240
rect 117750 675000 117860 675240
rect 118100 675000 118190 675240
rect 118430 675000 118520 675240
rect 118760 675000 118850 675240
rect 119090 675000 119200 675240
rect 119440 675000 119530 675240
rect 119770 675000 119860 675240
rect 120100 675000 120190 675240
rect 120430 675000 120540 675240
rect 120780 675000 120870 675240
rect 121110 675000 121200 675240
rect 121440 675000 121530 675240
rect 121770 675000 122190 675240
rect 122430 675000 122540 675240
rect 122780 675000 122870 675240
rect 123110 675000 123200 675240
rect 123440 675000 123530 675240
rect 123770 675000 123880 675240
rect 124120 675000 124210 675240
rect 124450 675000 124540 675240
rect 124780 675000 124870 675240
rect 125110 675000 125220 675240
rect 125460 675000 125550 675240
rect 125790 675000 125880 675240
rect 126120 675000 126210 675240
rect 126450 675000 126560 675240
rect 126800 675000 126890 675240
rect 127130 675000 127220 675240
rect 127460 675000 127550 675240
rect 127790 675000 127900 675240
rect 128140 675000 128230 675240
rect 128470 675000 128560 675240
rect 128800 675000 128890 675240
rect 129130 675000 129240 675240
rect 129480 675000 129570 675240
rect 129810 675000 129900 675240
rect 130140 675000 130230 675240
rect 130470 675000 130580 675240
rect 130820 675000 130910 675240
rect 131150 675000 131240 675240
rect 131480 675000 131570 675240
rect 131810 675000 131920 675240
rect 132160 675000 132250 675240
rect 132490 675000 132580 675240
rect 132820 675000 132910 675240
rect 133150 675000 133570 675240
rect 133810 675000 133920 675240
rect 134160 675000 134250 675240
rect 134490 675000 134580 675240
rect 134820 675000 134910 675240
rect 135150 675000 135260 675240
rect 135500 675000 135590 675240
rect 135830 675000 135920 675240
rect 136160 675000 136250 675240
rect 136490 675000 136600 675240
rect 136840 675000 136930 675240
rect 137170 675000 137260 675240
rect 137500 675000 137590 675240
rect 137830 675000 137940 675240
rect 138180 675000 138270 675240
rect 138510 675000 138600 675240
rect 138840 675000 138930 675240
rect 139170 675000 139280 675240
rect 139520 675000 139610 675240
rect 139850 675000 139940 675240
rect 140180 675000 140270 675240
rect 140510 675000 140620 675240
rect 140860 675000 140950 675240
rect 141190 675000 141280 675240
rect 141520 675000 141610 675240
rect 141850 675000 141960 675240
rect 142200 675000 142290 675240
rect 142530 675000 142620 675240
rect 142860 675000 142950 675240
rect 143190 675000 143300 675240
rect 143540 675000 143630 675240
rect 143870 675000 143960 675240
rect 144200 675000 144290 675240
rect 144530 675000 144950 675240
rect 145190 675000 145300 675240
rect 145540 675000 145630 675240
rect 145870 675000 145960 675240
rect 146200 675000 146290 675240
rect 146530 675000 146640 675240
rect 146880 675000 146970 675240
rect 147210 675000 147300 675240
rect 147540 675000 147630 675240
rect 147870 675000 147980 675240
rect 148220 675000 148310 675240
rect 148550 675000 148640 675240
rect 148880 675000 148970 675240
rect 149210 675000 149320 675240
rect 149560 675000 149650 675240
rect 149890 675000 149980 675240
rect 150220 675000 150310 675240
rect 150550 675000 150660 675240
rect 150900 675000 150990 675240
rect 151230 675000 151320 675240
rect 151560 675000 151650 675240
rect 151890 675000 152000 675240
rect 152240 675000 152330 675240
rect 152570 675000 152660 675240
rect 152900 675000 152990 675240
rect 153230 675000 153340 675240
rect 153580 675000 153670 675240
rect 153910 675000 154000 675240
rect 154240 675000 154330 675240
rect 154570 675000 154680 675240
rect 154920 675000 155010 675240
rect 155250 675000 155340 675240
rect 155580 675000 155670 675240
rect 155910 675000 155960 675240
rect 110760 674910 155960 675000
rect 110760 674670 110810 674910
rect 111050 674670 111160 674910
rect 111400 674670 111490 674910
rect 111730 674670 111820 674910
rect 112060 674670 112150 674910
rect 112390 674670 112500 674910
rect 112740 674670 112830 674910
rect 113070 674670 113160 674910
rect 113400 674670 113490 674910
rect 113730 674670 113840 674910
rect 114080 674670 114170 674910
rect 114410 674670 114500 674910
rect 114740 674670 114830 674910
rect 115070 674670 115180 674910
rect 115420 674670 115510 674910
rect 115750 674670 115840 674910
rect 116080 674670 116170 674910
rect 116410 674670 116520 674910
rect 116760 674670 116850 674910
rect 117090 674670 117180 674910
rect 117420 674670 117510 674910
rect 117750 674670 117860 674910
rect 118100 674670 118190 674910
rect 118430 674670 118520 674910
rect 118760 674670 118850 674910
rect 119090 674670 119200 674910
rect 119440 674670 119530 674910
rect 119770 674670 119860 674910
rect 120100 674670 120190 674910
rect 120430 674670 120540 674910
rect 120780 674670 120870 674910
rect 121110 674670 121200 674910
rect 121440 674670 121530 674910
rect 121770 674670 122190 674910
rect 122430 674670 122540 674910
rect 122780 674670 122870 674910
rect 123110 674670 123200 674910
rect 123440 674670 123530 674910
rect 123770 674670 123880 674910
rect 124120 674670 124210 674910
rect 124450 674670 124540 674910
rect 124780 674670 124870 674910
rect 125110 674670 125220 674910
rect 125460 674670 125550 674910
rect 125790 674670 125880 674910
rect 126120 674670 126210 674910
rect 126450 674670 126560 674910
rect 126800 674670 126890 674910
rect 127130 674670 127220 674910
rect 127460 674670 127550 674910
rect 127790 674670 127900 674910
rect 128140 674670 128230 674910
rect 128470 674670 128560 674910
rect 128800 674670 128890 674910
rect 129130 674670 129240 674910
rect 129480 674670 129570 674910
rect 129810 674670 129900 674910
rect 130140 674670 130230 674910
rect 130470 674670 130580 674910
rect 130820 674670 130910 674910
rect 131150 674670 131240 674910
rect 131480 674670 131570 674910
rect 131810 674670 131920 674910
rect 132160 674670 132250 674910
rect 132490 674670 132580 674910
rect 132820 674670 132910 674910
rect 133150 674670 133570 674910
rect 133810 674670 133920 674910
rect 134160 674670 134250 674910
rect 134490 674670 134580 674910
rect 134820 674670 134910 674910
rect 135150 674670 135260 674910
rect 135500 674670 135590 674910
rect 135830 674670 135920 674910
rect 136160 674670 136250 674910
rect 136490 674670 136600 674910
rect 136840 674670 136930 674910
rect 137170 674670 137260 674910
rect 137500 674670 137590 674910
rect 137830 674670 137940 674910
rect 138180 674670 138270 674910
rect 138510 674670 138600 674910
rect 138840 674670 138930 674910
rect 139170 674670 139280 674910
rect 139520 674670 139610 674910
rect 139850 674670 139940 674910
rect 140180 674670 140270 674910
rect 140510 674670 140620 674910
rect 140860 674670 140950 674910
rect 141190 674670 141280 674910
rect 141520 674670 141610 674910
rect 141850 674670 141960 674910
rect 142200 674670 142290 674910
rect 142530 674670 142620 674910
rect 142860 674670 142950 674910
rect 143190 674670 143300 674910
rect 143540 674670 143630 674910
rect 143870 674670 143960 674910
rect 144200 674670 144290 674910
rect 144530 674670 144950 674910
rect 145190 674670 145300 674910
rect 145540 674670 145630 674910
rect 145870 674670 145960 674910
rect 146200 674670 146290 674910
rect 146530 674670 146640 674910
rect 146880 674670 146970 674910
rect 147210 674670 147300 674910
rect 147540 674670 147630 674910
rect 147870 674670 147980 674910
rect 148220 674670 148310 674910
rect 148550 674670 148640 674910
rect 148880 674670 148970 674910
rect 149210 674670 149320 674910
rect 149560 674670 149650 674910
rect 149890 674670 149980 674910
rect 150220 674670 150310 674910
rect 150550 674670 150660 674910
rect 150900 674670 150990 674910
rect 151230 674670 151320 674910
rect 151560 674670 151650 674910
rect 151890 674670 152000 674910
rect 152240 674670 152330 674910
rect 152570 674670 152660 674910
rect 152900 674670 152990 674910
rect 153230 674670 153340 674910
rect 153580 674670 153670 674910
rect 153910 674670 154000 674910
rect 154240 674670 154330 674910
rect 154570 674670 154680 674910
rect 154920 674670 155010 674910
rect 155250 674670 155340 674910
rect 155580 674670 155670 674910
rect 155910 674670 155960 674910
rect 110760 674580 155960 674670
rect 110760 674340 110810 674580
rect 111050 674340 111160 674580
rect 111400 674340 111490 674580
rect 111730 674340 111820 674580
rect 112060 674340 112150 674580
rect 112390 674340 112500 674580
rect 112740 674340 112830 674580
rect 113070 674340 113160 674580
rect 113400 674340 113490 674580
rect 113730 674340 113840 674580
rect 114080 674340 114170 674580
rect 114410 674340 114500 674580
rect 114740 674340 114830 674580
rect 115070 674340 115180 674580
rect 115420 674340 115510 674580
rect 115750 674340 115840 674580
rect 116080 674340 116170 674580
rect 116410 674340 116520 674580
rect 116760 674340 116850 674580
rect 117090 674340 117180 674580
rect 117420 674340 117510 674580
rect 117750 674340 117860 674580
rect 118100 674340 118190 674580
rect 118430 674340 118520 674580
rect 118760 674340 118850 674580
rect 119090 674340 119200 674580
rect 119440 674340 119530 674580
rect 119770 674340 119860 674580
rect 120100 674340 120190 674580
rect 120430 674340 120540 674580
rect 120780 674340 120870 674580
rect 121110 674340 121200 674580
rect 121440 674340 121530 674580
rect 121770 674340 122190 674580
rect 122430 674340 122540 674580
rect 122780 674340 122870 674580
rect 123110 674340 123200 674580
rect 123440 674340 123530 674580
rect 123770 674340 123880 674580
rect 124120 674340 124210 674580
rect 124450 674340 124540 674580
rect 124780 674340 124870 674580
rect 125110 674340 125220 674580
rect 125460 674340 125550 674580
rect 125790 674340 125880 674580
rect 126120 674340 126210 674580
rect 126450 674340 126560 674580
rect 126800 674340 126890 674580
rect 127130 674340 127220 674580
rect 127460 674340 127550 674580
rect 127790 674340 127900 674580
rect 128140 674340 128230 674580
rect 128470 674340 128560 674580
rect 128800 674340 128890 674580
rect 129130 674340 129240 674580
rect 129480 674340 129570 674580
rect 129810 674340 129900 674580
rect 130140 674340 130230 674580
rect 130470 674340 130580 674580
rect 130820 674340 130910 674580
rect 131150 674340 131240 674580
rect 131480 674340 131570 674580
rect 131810 674340 131920 674580
rect 132160 674340 132250 674580
rect 132490 674340 132580 674580
rect 132820 674340 132910 674580
rect 133150 674340 133570 674580
rect 133810 674340 133920 674580
rect 134160 674340 134250 674580
rect 134490 674340 134580 674580
rect 134820 674340 134910 674580
rect 135150 674340 135260 674580
rect 135500 674340 135590 674580
rect 135830 674340 135920 674580
rect 136160 674340 136250 674580
rect 136490 674340 136600 674580
rect 136840 674340 136930 674580
rect 137170 674340 137260 674580
rect 137500 674340 137590 674580
rect 137830 674340 137940 674580
rect 138180 674340 138270 674580
rect 138510 674340 138600 674580
rect 138840 674340 138930 674580
rect 139170 674340 139280 674580
rect 139520 674340 139610 674580
rect 139850 674340 139940 674580
rect 140180 674340 140270 674580
rect 140510 674340 140620 674580
rect 140860 674340 140950 674580
rect 141190 674340 141280 674580
rect 141520 674340 141610 674580
rect 141850 674340 141960 674580
rect 142200 674340 142290 674580
rect 142530 674340 142620 674580
rect 142860 674340 142950 674580
rect 143190 674340 143300 674580
rect 143540 674340 143630 674580
rect 143870 674340 143960 674580
rect 144200 674340 144290 674580
rect 144530 674340 144950 674580
rect 145190 674340 145300 674580
rect 145540 674340 145630 674580
rect 145870 674340 145960 674580
rect 146200 674340 146290 674580
rect 146530 674340 146640 674580
rect 146880 674340 146970 674580
rect 147210 674340 147300 674580
rect 147540 674340 147630 674580
rect 147870 674340 147980 674580
rect 148220 674340 148310 674580
rect 148550 674340 148640 674580
rect 148880 674340 148970 674580
rect 149210 674340 149320 674580
rect 149560 674340 149650 674580
rect 149890 674340 149980 674580
rect 150220 674340 150310 674580
rect 150550 674340 150660 674580
rect 150900 674340 150990 674580
rect 151230 674340 151320 674580
rect 151560 674340 151650 674580
rect 151890 674340 152000 674580
rect 152240 674340 152330 674580
rect 152570 674340 152660 674580
rect 152900 674340 152990 674580
rect 153230 674340 153340 674580
rect 153580 674340 153670 674580
rect 153910 674340 154000 674580
rect 154240 674340 154330 674580
rect 154570 674340 154680 674580
rect 154920 674340 155010 674580
rect 155250 674340 155340 674580
rect 155580 674340 155670 674580
rect 155910 674340 155960 674580
rect 110760 674250 155960 674340
rect 110760 674010 110810 674250
rect 111050 674010 111160 674250
rect 111400 674010 111490 674250
rect 111730 674010 111820 674250
rect 112060 674010 112150 674250
rect 112390 674010 112500 674250
rect 112740 674010 112830 674250
rect 113070 674010 113160 674250
rect 113400 674010 113490 674250
rect 113730 674010 113840 674250
rect 114080 674010 114170 674250
rect 114410 674010 114500 674250
rect 114740 674010 114830 674250
rect 115070 674010 115180 674250
rect 115420 674010 115510 674250
rect 115750 674010 115840 674250
rect 116080 674010 116170 674250
rect 116410 674010 116520 674250
rect 116760 674010 116850 674250
rect 117090 674010 117180 674250
rect 117420 674010 117510 674250
rect 117750 674010 117860 674250
rect 118100 674010 118190 674250
rect 118430 674010 118520 674250
rect 118760 674010 118850 674250
rect 119090 674010 119200 674250
rect 119440 674010 119530 674250
rect 119770 674010 119860 674250
rect 120100 674010 120190 674250
rect 120430 674010 120540 674250
rect 120780 674010 120870 674250
rect 121110 674010 121200 674250
rect 121440 674010 121530 674250
rect 121770 674010 122190 674250
rect 122430 674010 122540 674250
rect 122780 674010 122870 674250
rect 123110 674010 123200 674250
rect 123440 674010 123530 674250
rect 123770 674010 123880 674250
rect 124120 674010 124210 674250
rect 124450 674010 124540 674250
rect 124780 674010 124870 674250
rect 125110 674010 125220 674250
rect 125460 674010 125550 674250
rect 125790 674010 125880 674250
rect 126120 674010 126210 674250
rect 126450 674010 126560 674250
rect 126800 674010 126890 674250
rect 127130 674010 127220 674250
rect 127460 674010 127550 674250
rect 127790 674010 127900 674250
rect 128140 674010 128230 674250
rect 128470 674010 128560 674250
rect 128800 674010 128890 674250
rect 129130 674010 129240 674250
rect 129480 674010 129570 674250
rect 129810 674010 129900 674250
rect 130140 674010 130230 674250
rect 130470 674010 130580 674250
rect 130820 674010 130910 674250
rect 131150 674010 131240 674250
rect 131480 674010 131570 674250
rect 131810 674010 131920 674250
rect 132160 674010 132250 674250
rect 132490 674010 132580 674250
rect 132820 674010 132910 674250
rect 133150 674010 133570 674250
rect 133810 674010 133920 674250
rect 134160 674010 134250 674250
rect 134490 674010 134580 674250
rect 134820 674010 134910 674250
rect 135150 674010 135260 674250
rect 135500 674010 135590 674250
rect 135830 674010 135920 674250
rect 136160 674010 136250 674250
rect 136490 674010 136600 674250
rect 136840 674010 136930 674250
rect 137170 674010 137260 674250
rect 137500 674010 137590 674250
rect 137830 674010 137940 674250
rect 138180 674010 138270 674250
rect 138510 674010 138600 674250
rect 138840 674010 138930 674250
rect 139170 674010 139280 674250
rect 139520 674010 139610 674250
rect 139850 674010 139940 674250
rect 140180 674010 140270 674250
rect 140510 674010 140620 674250
rect 140860 674010 140950 674250
rect 141190 674010 141280 674250
rect 141520 674010 141610 674250
rect 141850 674010 141960 674250
rect 142200 674010 142290 674250
rect 142530 674010 142620 674250
rect 142860 674010 142950 674250
rect 143190 674010 143300 674250
rect 143540 674010 143630 674250
rect 143870 674010 143960 674250
rect 144200 674010 144290 674250
rect 144530 674010 144950 674250
rect 145190 674010 145300 674250
rect 145540 674010 145630 674250
rect 145870 674010 145960 674250
rect 146200 674010 146290 674250
rect 146530 674010 146640 674250
rect 146880 674010 146970 674250
rect 147210 674010 147300 674250
rect 147540 674010 147630 674250
rect 147870 674010 147980 674250
rect 148220 674010 148310 674250
rect 148550 674010 148640 674250
rect 148880 674010 148970 674250
rect 149210 674010 149320 674250
rect 149560 674010 149650 674250
rect 149890 674010 149980 674250
rect 150220 674010 150310 674250
rect 150550 674010 150660 674250
rect 150900 674010 150990 674250
rect 151230 674010 151320 674250
rect 151560 674010 151650 674250
rect 151890 674010 152000 674250
rect 152240 674010 152330 674250
rect 152570 674010 152660 674250
rect 152900 674010 152990 674250
rect 153230 674010 153340 674250
rect 153580 674010 153670 674250
rect 153910 674010 154000 674250
rect 154240 674010 154330 674250
rect 154570 674010 154680 674250
rect 154920 674010 155010 674250
rect 155250 674010 155340 674250
rect 155580 674010 155670 674250
rect 155910 674010 155960 674250
rect 157440 678979 186713 679147
rect 157440 678739 157520 678979
rect 157780 678739 157880 678979
rect 158140 678739 158240 678979
rect 158500 678739 158600 678979
rect 158860 678739 186713 678979
rect 157440 678639 186713 678739
rect 157440 678399 157520 678639
rect 157780 678399 157880 678639
rect 158140 678399 158240 678639
rect 158500 678399 158600 678639
rect 158860 678399 186713 678639
rect 157440 678299 186713 678399
rect 157440 678059 157520 678299
rect 157780 678059 157880 678299
rect 158140 678059 158240 678299
rect 158500 678059 158600 678299
rect 158860 678059 186713 678299
rect 157440 677959 186713 678059
rect 157440 677719 157520 677959
rect 157780 677719 157880 677959
rect 158140 677719 158240 677959
rect 158500 677719 158600 677959
rect 158860 677719 186713 677959
rect 157440 677619 186713 677719
rect 157440 677379 157520 677619
rect 157780 677379 157880 677619
rect 158140 677379 158240 677619
rect 158500 677379 158600 677619
rect 158860 677379 186713 677619
rect 157440 677279 186713 677379
rect 157440 677039 157520 677279
rect 157780 677039 157880 677279
rect 158140 677039 158240 677279
rect 158500 677039 158600 677279
rect 158860 677039 186713 677279
rect 157440 676939 186713 677039
rect 157440 676699 157520 676939
rect 157780 676699 157880 676939
rect 158140 676699 158240 676939
rect 158500 676699 158600 676939
rect 158860 676699 186713 676939
rect 157440 676599 186713 676699
rect 157440 676359 157520 676599
rect 157780 676359 157880 676599
rect 158140 676359 158240 676599
rect 158500 676359 158600 676599
rect 158860 676359 186713 676599
rect 157440 676259 186713 676359
rect 157440 676019 157520 676259
rect 157780 676019 157880 676259
rect 158140 676019 158240 676259
rect 158500 676019 158600 676259
rect 158860 676019 186713 676259
rect 157440 675919 186713 676019
rect 157440 675679 157520 675919
rect 157780 675679 157880 675919
rect 158140 675679 158240 675919
rect 158500 675679 158600 675919
rect 158860 675679 186713 675919
rect 157440 675579 186713 675679
rect 157440 675339 157520 675579
rect 157780 675339 157880 675579
rect 158140 675339 158240 675579
rect 158500 675339 158600 675579
rect 158860 675339 186713 675579
rect 157440 675239 186713 675339
rect 157440 674999 157520 675239
rect 157780 674999 157880 675239
rect 158140 674999 158240 675239
rect 158500 674999 158600 675239
rect 158860 674999 186713 675239
rect 157440 674899 186713 674999
rect 157440 674659 157520 674899
rect 157780 674659 157880 674899
rect 158140 674659 158240 674899
rect 158500 674659 158600 674899
rect 158860 674659 186713 674899
rect 157440 674559 186713 674659
rect 157440 674319 157520 674559
rect 157780 674319 157880 674559
rect 158140 674319 158240 674559
rect 158500 674319 158600 674559
rect 158860 674319 186713 674559
rect 157440 674152 186713 674319
rect 110760 673900 155960 674010
rect 110760 673660 110810 673900
rect 111050 673660 111160 673900
rect 111400 673660 111490 673900
rect 111730 673660 111820 673900
rect 112060 673660 112150 673900
rect 112390 673660 112500 673900
rect 112740 673660 112830 673900
rect 113070 673660 113160 673900
rect 113400 673660 113490 673900
rect 113730 673660 113840 673900
rect 114080 673660 114170 673900
rect 114410 673660 114500 673900
rect 114740 673660 114830 673900
rect 115070 673660 115180 673900
rect 115420 673660 115510 673900
rect 115750 673660 115840 673900
rect 116080 673660 116170 673900
rect 116410 673660 116520 673900
rect 116760 673660 116850 673900
rect 117090 673660 117180 673900
rect 117420 673660 117510 673900
rect 117750 673660 117860 673900
rect 118100 673660 118190 673900
rect 118430 673660 118520 673900
rect 118760 673660 118850 673900
rect 119090 673660 119200 673900
rect 119440 673660 119530 673900
rect 119770 673660 119860 673900
rect 120100 673660 120190 673900
rect 120430 673660 120540 673900
rect 120780 673660 120870 673900
rect 121110 673660 121200 673900
rect 121440 673660 121530 673900
rect 121770 673660 122190 673900
rect 122430 673660 122540 673900
rect 122780 673660 122870 673900
rect 123110 673660 123200 673900
rect 123440 673660 123530 673900
rect 123770 673660 123880 673900
rect 124120 673660 124210 673900
rect 124450 673660 124540 673900
rect 124780 673660 124870 673900
rect 125110 673660 125220 673900
rect 125460 673660 125550 673900
rect 125790 673660 125880 673900
rect 126120 673660 126210 673900
rect 126450 673660 126560 673900
rect 126800 673660 126890 673900
rect 127130 673660 127220 673900
rect 127460 673660 127550 673900
rect 127790 673660 127900 673900
rect 128140 673660 128230 673900
rect 128470 673660 128560 673900
rect 128800 673660 128890 673900
rect 129130 673660 129240 673900
rect 129480 673660 129570 673900
rect 129810 673660 129900 673900
rect 130140 673660 130230 673900
rect 130470 673660 130580 673900
rect 130820 673660 130910 673900
rect 131150 673660 131240 673900
rect 131480 673660 131570 673900
rect 131810 673660 131920 673900
rect 132160 673660 132250 673900
rect 132490 673660 132580 673900
rect 132820 673660 132910 673900
rect 133150 673660 133570 673900
rect 133810 673660 133920 673900
rect 134160 673660 134250 673900
rect 134490 673660 134580 673900
rect 134820 673660 134910 673900
rect 135150 673660 135260 673900
rect 135500 673660 135590 673900
rect 135830 673660 135920 673900
rect 136160 673660 136250 673900
rect 136490 673660 136600 673900
rect 136840 673660 136930 673900
rect 137170 673660 137260 673900
rect 137500 673660 137590 673900
rect 137830 673660 137940 673900
rect 138180 673660 138270 673900
rect 138510 673660 138600 673900
rect 138840 673660 138930 673900
rect 139170 673660 139280 673900
rect 139520 673660 139610 673900
rect 139850 673660 139940 673900
rect 140180 673660 140270 673900
rect 140510 673660 140620 673900
rect 140860 673660 140950 673900
rect 141190 673660 141280 673900
rect 141520 673660 141610 673900
rect 141850 673660 141960 673900
rect 142200 673660 142290 673900
rect 142530 673660 142620 673900
rect 142860 673660 142950 673900
rect 143190 673660 143300 673900
rect 143540 673660 143630 673900
rect 143870 673660 143960 673900
rect 144200 673660 144290 673900
rect 144530 673660 144950 673900
rect 145190 673660 145300 673900
rect 145540 673660 145630 673900
rect 145870 673660 145960 673900
rect 146200 673660 146290 673900
rect 146530 673660 146640 673900
rect 146880 673660 146970 673900
rect 147210 673660 147300 673900
rect 147540 673660 147630 673900
rect 147870 673660 147980 673900
rect 148220 673660 148310 673900
rect 148550 673660 148640 673900
rect 148880 673660 148970 673900
rect 149210 673660 149320 673900
rect 149560 673660 149650 673900
rect 149890 673660 149980 673900
rect 150220 673660 150310 673900
rect 150550 673660 150660 673900
rect 150900 673660 150990 673900
rect 151230 673660 151320 673900
rect 151560 673660 151650 673900
rect 151890 673660 152000 673900
rect 152240 673660 152330 673900
rect 152570 673660 152660 673900
rect 152900 673660 152990 673900
rect 153230 673660 153340 673900
rect 153580 673660 153670 673900
rect 153910 673660 154000 673900
rect 154240 673660 154330 673900
rect 154570 673660 154680 673900
rect 154920 673660 155010 673900
rect 155250 673660 155340 673900
rect 155580 673660 155670 673900
rect 155910 673660 155960 673900
rect 110760 673570 155960 673660
rect 110760 673330 110810 673570
rect 111050 673330 111160 673570
rect 111400 673330 111490 673570
rect 111730 673330 111820 673570
rect 112060 673330 112150 673570
rect 112390 673330 112500 673570
rect 112740 673330 112830 673570
rect 113070 673330 113160 673570
rect 113400 673330 113490 673570
rect 113730 673330 113840 673570
rect 114080 673330 114170 673570
rect 114410 673330 114500 673570
rect 114740 673330 114830 673570
rect 115070 673330 115180 673570
rect 115420 673330 115510 673570
rect 115750 673330 115840 673570
rect 116080 673330 116170 673570
rect 116410 673330 116520 673570
rect 116760 673330 116850 673570
rect 117090 673330 117180 673570
rect 117420 673330 117510 673570
rect 117750 673330 117860 673570
rect 118100 673330 118190 673570
rect 118430 673330 118520 673570
rect 118760 673330 118850 673570
rect 119090 673330 119200 673570
rect 119440 673330 119530 673570
rect 119770 673330 119860 673570
rect 120100 673330 120190 673570
rect 120430 673330 120540 673570
rect 120780 673330 120870 673570
rect 121110 673330 121200 673570
rect 121440 673330 121530 673570
rect 121770 673330 122190 673570
rect 122430 673330 122540 673570
rect 122780 673330 122870 673570
rect 123110 673330 123200 673570
rect 123440 673330 123530 673570
rect 123770 673330 123880 673570
rect 124120 673330 124210 673570
rect 124450 673330 124540 673570
rect 124780 673330 124870 673570
rect 125110 673330 125220 673570
rect 125460 673330 125550 673570
rect 125790 673330 125880 673570
rect 126120 673330 126210 673570
rect 126450 673330 126560 673570
rect 126800 673330 126890 673570
rect 127130 673330 127220 673570
rect 127460 673330 127550 673570
rect 127790 673330 127900 673570
rect 128140 673330 128230 673570
rect 128470 673330 128560 673570
rect 128800 673330 128890 673570
rect 129130 673330 129240 673570
rect 129480 673330 129570 673570
rect 129810 673330 129900 673570
rect 130140 673330 130230 673570
rect 130470 673330 130580 673570
rect 130820 673330 130910 673570
rect 131150 673330 131240 673570
rect 131480 673330 131570 673570
rect 131810 673330 131920 673570
rect 132160 673330 132250 673570
rect 132490 673330 132580 673570
rect 132820 673330 132910 673570
rect 133150 673330 133570 673570
rect 133810 673330 133920 673570
rect 134160 673330 134250 673570
rect 134490 673330 134580 673570
rect 134820 673330 134910 673570
rect 135150 673330 135260 673570
rect 135500 673330 135590 673570
rect 135830 673330 135920 673570
rect 136160 673330 136250 673570
rect 136490 673330 136600 673570
rect 136840 673330 136930 673570
rect 137170 673330 137260 673570
rect 137500 673330 137590 673570
rect 137830 673330 137940 673570
rect 138180 673330 138270 673570
rect 138510 673330 138600 673570
rect 138840 673330 138930 673570
rect 139170 673330 139280 673570
rect 139520 673330 139610 673570
rect 139850 673330 139940 673570
rect 140180 673330 140270 673570
rect 140510 673330 140620 673570
rect 140860 673330 140950 673570
rect 141190 673330 141280 673570
rect 141520 673330 141610 673570
rect 141850 673330 141960 673570
rect 142200 673330 142290 673570
rect 142530 673330 142620 673570
rect 142860 673330 142950 673570
rect 143190 673330 143300 673570
rect 143540 673330 143630 673570
rect 143870 673330 143960 673570
rect 144200 673330 144290 673570
rect 144530 673330 144950 673570
rect 145190 673330 145300 673570
rect 145540 673330 145630 673570
rect 145870 673330 145960 673570
rect 146200 673330 146290 673570
rect 146530 673330 146640 673570
rect 146880 673330 146970 673570
rect 147210 673330 147300 673570
rect 147540 673330 147630 673570
rect 147870 673330 147980 673570
rect 148220 673330 148310 673570
rect 148550 673330 148640 673570
rect 148880 673330 148970 673570
rect 149210 673330 149320 673570
rect 149560 673330 149650 673570
rect 149890 673330 149980 673570
rect 150220 673330 150310 673570
rect 150550 673330 150660 673570
rect 150900 673330 150990 673570
rect 151230 673330 151320 673570
rect 151560 673330 151650 673570
rect 151890 673330 152000 673570
rect 152240 673330 152330 673570
rect 152570 673330 152660 673570
rect 152900 673330 152990 673570
rect 153230 673330 153340 673570
rect 153580 673330 153670 673570
rect 153910 673330 154000 673570
rect 154240 673330 154330 673570
rect 154570 673330 154680 673570
rect 154920 673330 155010 673570
rect 155250 673330 155340 673570
rect 155580 673330 155670 673570
rect 155910 673330 155960 673570
rect 110760 673240 155960 673330
rect 110760 673000 110810 673240
rect 111050 673000 111160 673240
rect 111400 673000 111490 673240
rect 111730 673000 111820 673240
rect 112060 673000 112150 673240
rect 112390 673000 112500 673240
rect 112740 673000 112830 673240
rect 113070 673000 113160 673240
rect 113400 673000 113490 673240
rect 113730 673000 113840 673240
rect 114080 673000 114170 673240
rect 114410 673000 114500 673240
rect 114740 673000 114830 673240
rect 115070 673000 115180 673240
rect 115420 673000 115510 673240
rect 115750 673000 115840 673240
rect 116080 673000 116170 673240
rect 116410 673000 116520 673240
rect 116760 673000 116850 673240
rect 117090 673000 117180 673240
rect 117420 673000 117510 673240
rect 117750 673000 117860 673240
rect 118100 673000 118190 673240
rect 118430 673000 118520 673240
rect 118760 673000 118850 673240
rect 119090 673000 119200 673240
rect 119440 673000 119530 673240
rect 119770 673000 119860 673240
rect 120100 673000 120190 673240
rect 120430 673000 120540 673240
rect 120780 673000 120870 673240
rect 121110 673000 121200 673240
rect 121440 673000 121530 673240
rect 121770 673000 122190 673240
rect 122430 673000 122540 673240
rect 122780 673000 122870 673240
rect 123110 673000 123200 673240
rect 123440 673000 123530 673240
rect 123770 673000 123880 673240
rect 124120 673000 124210 673240
rect 124450 673000 124540 673240
rect 124780 673000 124870 673240
rect 125110 673000 125220 673240
rect 125460 673000 125550 673240
rect 125790 673000 125880 673240
rect 126120 673000 126210 673240
rect 126450 673000 126560 673240
rect 126800 673000 126890 673240
rect 127130 673000 127220 673240
rect 127460 673000 127550 673240
rect 127790 673000 127900 673240
rect 128140 673000 128230 673240
rect 128470 673000 128560 673240
rect 128800 673000 128890 673240
rect 129130 673000 129240 673240
rect 129480 673000 129570 673240
rect 129810 673000 129900 673240
rect 130140 673000 130230 673240
rect 130470 673000 130580 673240
rect 130820 673000 130910 673240
rect 131150 673000 131240 673240
rect 131480 673000 131570 673240
rect 131810 673000 131920 673240
rect 132160 673000 132250 673240
rect 132490 673000 132580 673240
rect 132820 673000 132910 673240
rect 133150 673000 133570 673240
rect 133810 673000 133920 673240
rect 134160 673000 134250 673240
rect 134490 673000 134580 673240
rect 134820 673000 134910 673240
rect 135150 673000 135260 673240
rect 135500 673000 135590 673240
rect 135830 673000 135920 673240
rect 136160 673000 136250 673240
rect 136490 673000 136600 673240
rect 136840 673000 136930 673240
rect 137170 673000 137260 673240
rect 137500 673000 137590 673240
rect 137830 673000 137940 673240
rect 138180 673000 138270 673240
rect 138510 673000 138600 673240
rect 138840 673000 138930 673240
rect 139170 673000 139280 673240
rect 139520 673000 139610 673240
rect 139850 673000 139940 673240
rect 140180 673000 140270 673240
rect 140510 673000 140620 673240
rect 140860 673000 140950 673240
rect 141190 673000 141280 673240
rect 141520 673000 141610 673240
rect 141850 673000 141960 673240
rect 142200 673000 142290 673240
rect 142530 673000 142620 673240
rect 142860 673000 142950 673240
rect 143190 673000 143300 673240
rect 143540 673000 143630 673240
rect 143870 673000 143960 673240
rect 144200 673000 144290 673240
rect 144530 673000 144950 673240
rect 145190 673000 145300 673240
rect 145540 673000 145630 673240
rect 145870 673000 145960 673240
rect 146200 673000 146290 673240
rect 146530 673000 146640 673240
rect 146880 673000 146970 673240
rect 147210 673000 147300 673240
rect 147540 673000 147630 673240
rect 147870 673000 147980 673240
rect 148220 673000 148310 673240
rect 148550 673000 148640 673240
rect 148880 673000 148970 673240
rect 149210 673000 149320 673240
rect 149560 673000 149650 673240
rect 149890 673000 149980 673240
rect 150220 673000 150310 673240
rect 150550 673000 150660 673240
rect 150900 673000 150990 673240
rect 151230 673000 151320 673240
rect 151560 673000 151650 673240
rect 151890 673000 152000 673240
rect 152240 673000 152330 673240
rect 152570 673000 152660 673240
rect 152900 673000 152990 673240
rect 153230 673000 153340 673240
rect 153580 673000 153670 673240
rect 153910 673000 154000 673240
rect 154240 673000 154330 673240
rect 154570 673000 154680 673240
rect 154920 673000 155010 673240
rect 155250 673000 155340 673240
rect 155580 673000 155670 673240
rect 155910 673000 155960 673240
rect 110760 672910 155960 673000
rect 110760 672670 110810 672910
rect 111050 672670 111160 672910
rect 111400 672670 111490 672910
rect 111730 672670 111820 672910
rect 112060 672670 112150 672910
rect 112390 672670 112500 672910
rect 112740 672670 112830 672910
rect 113070 672670 113160 672910
rect 113400 672670 113490 672910
rect 113730 672670 113840 672910
rect 114080 672670 114170 672910
rect 114410 672670 114500 672910
rect 114740 672670 114830 672910
rect 115070 672670 115180 672910
rect 115420 672670 115510 672910
rect 115750 672670 115840 672910
rect 116080 672670 116170 672910
rect 116410 672670 116520 672910
rect 116760 672670 116850 672910
rect 117090 672670 117180 672910
rect 117420 672670 117510 672910
rect 117750 672670 117860 672910
rect 118100 672670 118190 672910
rect 118430 672670 118520 672910
rect 118760 672670 118850 672910
rect 119090 672670 119200 672910
rect 119440 672670 119530 672910
rect 119770 672670 119860 672910
rect 120100 672670 120190 672910
rect 120430 672670 120540 672910
rect 120780 672670 120870 672910
rect 121110 672670 121200 672910
rect 121440 672670 121530 672910
rect 121770 672670 122190 672910
rect 122430 672670 122540 672910
rect 122780 672670 122870 672910
rect 123110 672670 123200 672910
rect 123440 672670 123530 672910
rect 123770 672670 123880 672910
rect 124120 672670 124210 672910
rect 124450 672670 124540 672910
rect 124780 672670 124870 672910
rect 125110 672670 125220 672910
rect 125460 672670 125550 672910
rect 125790 672670 125880 672910
rect 126120 672670 126210 672910
rect 126450 672670 126560 672910
rect 126800 672670 126890 672910
rect 127130 672670 127220 672910
rect 127460 672670 127550 672910
rect 127790 672670 127900 672910
rect 128140 672670 128230 672910
rect 128470 672670 128560 672910
rect 128800 672670 128890 672910
rect 129130 672670 129240 672910
rect 129480 672670 129570 672910
rect 129810 672670 129900 672910
rect 130140 672670 130230 672910
rect 130470 672670 130580 672910
rect 130820 672670 130910 672910
rect 131150 672670 131240 672910
rect 131480 672670 131570 672910
rect 131810 672670 131920 672910
rect 132160 672670 132250 672910
rect 132490 672670 132580 672910
rect 132820 672670 132910 672910
rect 133150 672670 133570 672910
rect 133810 672670 133920 672910
rect 134160 672670 134250 672910
rect 134490 672670 134580 672910
rect 134820 672670 134910 672910
rect 135150 672670 135260 672910
rect 135500 672670 135590 672910
rect 135830 672670 135920 672910
rect 136160 672670 136250 672910
rect 136490 672670 136600 672910
rect 136840 672670 136930 672910
rect 137170 672670 137260 672910
rect 137500 672670 137590 672910
rect 137830 672670 137940 672910
rect 138180 672670 138270 672910
rect 138510 672670 138600 672910
rect 138840 672670 138930 672910
rect 139170 672670 139280 672910
rect 139520 672670 139610 672910
rect 139850 672670 139940 672910
rect 140180 672670 140270 672910
rect 140510 672670 140620 672910
rect 140860 672670 140950 672910
rect 141190 672670 141280 672910
rect 141520 672670 141610 672910
rect 141850 672670 141960 672910
rect 142200 672670 142290 672910
rect 142530 672670 142620 672910
rect 142860 672670 142950 672910
rect 143190 672670 143300 672910
rect 143540 672670 143630 672910
rect 143870 672670 143960 672910
rect 144200 672670 144290 672910
rect 144530 672670 144950 672910
rect 145190 672670 145300 672910
rect 145540 672670 145630 672910
rect 145870 672670 145960 672910
rect 146200 672670 146290 672910
rect 146530 672670 146640 672910
rect 146880 672670 146970 672910
rect 147210 672670 147300 672910
rect 147540 672670 147630 672910
rect 147870 672670 147980 672910
rect 148220 672670 148310 672910
rect 148550 672670 148640 672910
rect 148880 672670 148970 672910
rect 149210 672670 149320 672910
rect 149560 672670 149650 672910
rect 149890 672670 149980 672910
rect 150220 672670 150310 672910
rect 150550 672670 150660 672910
rect 150900 672670 150990 672910
rect 151230 672670 151320 672910
rect 151560 672670 151650 672910
rect 151890 672670 152000 672910
rect 152240 672670 152330 672910
rect 152570 672670 152660 672910
rect 152900 672670 152990 672910
rect 153230 672670 153340 672910
rect 153580 672670 153670 672910
rect 153910 672670 154000 672910
rect 154240 672670 154330 672910
rect 154570 672670 154680 672910
rect 154920 672670 155010 672910
rect 155250 672670 155340 672910
rect 155580 672670 155670 672910
rect 155910 672670 155960 672910
rect 110760 672560 155960 672670
rect 110760 672320 110810 672560
rect 111050 672320 111160 672560
rect 111400 672320 111490 672560
rect 111730 672320 111820 672560
rect 112060 672320 112150 672560
rect 112390 672320 112500 672560
rect 112740 672320 112830 672560
rect 113070 672320 113160 672560
rect 113400 672320 113490 672560
rect 113730 672320 113840 672560
rect 114080 672320 114170 672560
rect 114410 672320 114500 672560
rect 114740 672320 114830 672560
rect 115070 672320 115180 672560
rect 115420 672320 115510 672560
rect 115750 672320 115840 672560
rect 116080 672320 116170 672560
rect 116410 672320 116520 672560
rect 116760 672320 116850 672560
rect 117090 672320 117180 672560
rect 117420 672320 117510 672560
rect 117750 672320 117860 672560
rect 118100 672320 118190 672560
rect 118430 672320 118520 672560
rect 118760 672320 118850 672560
rect 119090 672320 119200 672560
rect 119440 672320 119530 672560
rect 119770 672320 119860 672560
rect 120100 672320 120190 672560
rect 120430 672320 120540 672560
rect 120780 672320 120870 672560
rect 121110 672320 121200 672560
rect 121440 672320 121530 672560
rect 121770 672320 122190 672560
rect 122430 672320 122540 672560
rect 122780 672320 122870 672560
rect 123110 672320 123200 672560
rect 123440 672320 123530 672560
rect 123770 672320 123880 672560
rect 124120 672320 124210 672560
rect 124450 672320 124540 672560
rect 124780 672320 124870 672560
rect 125110 672320 125220 672560
rect 125460 672320 125550 672560
rect 125790 672320 125880 672560
rect 126120 672320 126210 672560
rect 126450 672320 126560 672560
rect 126800 672320 126890 672560
rect 127130 672320 127220 672560
rect 127460 672320 127550 672560
rect 127790 672320 127900 672560
rect 128140 672320 128230 672560
rect 128470 672320 128560 672560
rect 128800 672320 128890 672560
rect 129130 672320 129240 672560
rect 129480 672320 129570 672560
rect 129810 672320 129900 672560
rect 130140 672320 130230 672560
rect 130470 672320 130580 672560
rect 130820 672320 130910 672560
rect 131150 672320 131240 672560
rect 131480 672320 131570 672560
rect 131810 672320 131920 672560
rect 132160 672320 132250 672560
rect 132490 672320 132580 672560
rect 132820 672320 132910 672560
rect 133150 672320 133570 672560
rect 133810 672320 133920 672560
rect 134160 672320 134250 672560
rect 134490 672320 134580 672560
rect 134820 672320 134910 672560
rect 135150 672320 135260 672560
rect 135500 672320 135590 672560
rect 135830 672320 135920 672560
rect 136160 672320 136250 672560
rect 136490 672320 136600 672560
rect 136840 672320 136930 672560
rect 137170 672320 137260 672560
rect 137500 672320 137590 672560
rect 137830 672320 137940 672560
rect 138180 672320 138270 672560
rect 138510 672320 138600 672560
rect 138840 672320 138930 672560
rect 139170 672320 139280 672560
rect 139520 672320 139610 672560
rect 139850 672320 139940 672560
rect 140180 672320 140270 672560
rect 140510 672320 140620 672560
rect 140860 672320 140950 672560
rect 141190 672320 141280 672560
rect 141520 672320 141610 672560
rect 141850 672320 141960 672560
rect 142200 672320 142290 672560
rect 142530 672320 142620 672560
rect 142860 672320 142950 672560
rect 143190 672320 143300 672560
rect 143540 672320 143630 672560
rect 143870 672320 143960 672560
rect 144200 672320 144290 672560
rect 144530 672320 144950 672560
rect 145190 672320 145300 672560
rect 145540 672320 145630 672560
rect 145870 672320 145960 672560
rect 146200 672320 146290 672560
rect 146530 672320 146640 672560
rect 146880 672320 146970 672560
rect 147210 672320 147300 672560
rect 147540 672320 147630 672560
rect 147870 672320 147980 672560
rect 148220 672320 148310 672560
rect 148550 672320 148640 672560
rect 148880 672320 148970 672560
rect 149210 672320 149320 672560
rect 149560 672320 149650 672560
rect 149890 672320 149980 672560
rect 150220 672320 150310 672560
rect 150550 672320 150660 672560
rect 150900 672320 150990 672560
rect 151230 672320 151320 672560
rect 151560 672320 151650 672560
rect 151890 672320 152000 672560
rect 152240 672320 152330 672560
rect 152570 672320 152660 672560
rect 152900 672320 152990 672560
rect 153230 672320 153340 672560
rect 153580 672320 153670 672560
rect 153910 672320 154000 672560
rect 154240 672320 154330 672560
rect 154570 672320 154680 672560
rect 154920 672320 155010 672560
rect 155250 672320 155340 672560
rect 155580 672320 155670 672560
rect 155910 672320 155960 672560
rect 110760 671900 155960 672320
rect 110760 671660 110810 671900
rect 111050 671660 111140 671900
rect 111380 671660 111470 671900
rect 111710 671660 111800 671900
rect 112040 671660 112150 671900
rect 112390 671660 112480 671900
rect 112720 671660 112810 671900
rect 113050 671660 113140 671900
rect 113380 671660 113490 671900
rect 113730 671660 113820 671900
rect 114060 671660 114150 671900
rect 114390 671660 114480 671900
rect 114720 671660 114830 671900
rect 115070 671660 115160 671900
rect 115400 671660 115490 671900
rect 115730 671660 115820 671900
rect 116060 671660 116170 671900
rect 116410 671660 116500 671900
rect 116740 671660 116830 671900
rect 117070 671660 117160 671900
rect 117400 671660 117510 671900
rect 117750 671660 117840 671900
rect 118080 671660 118170 671900
rect 118410 671660 118500 671900
rect 118740 671660 118850 671900
rect 119090 671660 119180 671900
rect 119420 671660 119510 671900
rect 119750 671660 119840 671900
rect 120080 671660 120190 671900
rect 120430 671660 120520 671900
rect 120760 671660 120850 671900
rect 121090 671660 121180 671900
rect 121420 671660 121530 671900
rect 121770 671660 122190 671900
rect 122430 671660 122520 671900
rect 122760 671660 122850 671900
rect 123090 671660 123180 671900
rect 123420 671660 123530 671900
rect 123770 671660 123860 671900
rect 124100 671660 124190 671900
rect 124430 671660 124520 671900
rect 124760 671660 124870 671900
rect 125110 671660 125200 671900
rect 125440 671660 125530 671900
rect 125770 671660 125860 671900
rect 126100 671660 126210 671900
rect 126450 671660 126540 671900
rect 126780 671660 126870 671900
rect 127110 671660 127200 671900
rect 127440 671660 127550 671900
rect 127790 671660 127880 671900
rect 128120 671660 128210 671900
rect 128450 671660 128540 671900
rect 128780 671660 128890 671900
rect 129130 671660 129220 671900
rect 129460 671660 129550 671900
rect 129790 671660 129880 671900
rect 130120 671660 130230 671900
rect 130470 671660 130560 671900
rect 130800 671660 130890 671900
rect 131130 671660 131220 671900
rect 131460 671660 131570 671900
rect 131810 671660 131900 671900
rect 132140 671660 132230 671900
rect 132470 671660 132560 671900
rect 132800 671660 132910 671900
rect 133150 671660 133570 671900
rect 133810 671660 133900 671900
rect 134140 671660 134230 671900
rect 134470 671660 134560 671900
rect 134800 671660 134910 671900
rect 135150 671660 135240 671900
rect 135480 671660 135570 671900
rect 135810 671660 135900 671900
rect 136140 671660 136250 671900
rect 136490 671660 136580 671900
rect 136820 671660 136910 671900
rect 137150 671660 137240 671900
rect 137480 671660 137590 671900
rect 137830 671660 137920 671900
rect 138160 671660 138250 671900
rect 138490 671660 138580 671900
rect 138820 671660 138930 671900
rect 139170 671660 139260 671900
rect 139500 671660 139590 671900
rect 139830 671660 139920 671900
rect 140160 671660 140270 671900
rect 140510 671660 140600 671900
rect 140840 671660 140930 671900
rect 141170 671660 141260 671900
rect 141500 671660 141610 671900
rect 141850 671660 141940 671900
rect 142180 671660 142270 671900
rect 142510 671660 142600 671900
rect 142840 671660 142950 671900
rect 143190 671660 143280 671900
rect 143520 671660 143610 671900
rect 143850 671660 143940 671900
rect 144180 671660 144290 671900
rect 144530 671660 144950 671900
rect 145190 671660 145280 671900
rect 145520 671660 145610 671900
rect 145850 671660 145940 671900
rect 146180 671660 146290 671900
rect 146530 671660 146620 671900
rect 146860 671660 146950 671900
rect 147190 671660 147280 671900
rect 147520 671660 147630 671900
rect 147870 671660 147960 671900
rect 148200 671660 148290 671900
rect 148530 671660 148620 671900
rect 148860 671660 148970 671900
rect 149210 671660 149300 671900
rect 149540 671660 149630 671900
rect 149870 671660 149960 671900
rect 150200 671660 150310 671900
rect 150550 671660 150640 671900
rect 150880 671660 150970 671900
rect 151210 671660 151300 671900
rect 151540 671660 151650 671900
rect 151890 671660 151980 671900
rect 152220 671660 152310 671900
rect 152550 671660 152640 671900
rect 152880 671660 152990 671900
rect 153230 671660 153320 671900
rect 153560 671660 153650 671900
rect 153890 671660 153980 671900
rect 154220 671660 154330 671900
rect 154570 671660 154660 671900
rect 154900 671660 154990 671900
rect 155230 671660 155320 671900
rect 155560 671660 155670 671900
rect 155910 671660 155960 671900
rect 110760 671550 155960 671660
rect 110760 671310 110810 671550
rect 111050 671310 111140 671550
rect 111380 671310 111470 671550
rect 111710 671310 111800 671550
rect 112040 671310 112150 671550
rect 112390 671310 112480 671550
rect 112720 671310 112810 671550
rect 113050 671310 113140 671550
rect 113380 671310 113490 671550
rect 113730 671310 113820 671550
rect 114060 671310 114150 671550
rect 114390 671310 114480 671550
rect 114720 671310 114830 671550
rect 115070 671310 115160 671550
rect 115400 671310 115490 671550
rect 115730 671310 115820 671550
rect 116060 671310 116170 671550
rect 116410 671310 116500 671550
rect 116740 671310 116830 671550
rect 117070 671310 117160 671550
rect 117400 671310 117510 671550
rect 117750 671310 117840 671550
rect 118080 671310 118170 671550
rect 118410 671310 118500 671550
rect 118740 671310 118850 671550
rect 119090 671310 119180 671550
rect 119420 671310 119510 671550
rect 119750 671310 119840 671550
rect 120080 671310 120190 671550
rect 120430 671310 120520 671550
rect 120760 671310 120850 671550
rect 121090 671310 121180 671550
rect 121420 671310 121530 671550
rect 121770 671310 122190 671550
rect 122430 671310 122520 671550
rect 122760 671310 122850 671550
rect 123090 671310 123180 671550
rect 123420 671310 123530 671550
rect 123770 671310 123860 671550
rect 124100 671310 124190 671550
rect 124430 671310 124520 671550
rect 124760 671310 124870 671550
rect 125110 671310 125200 671550
rect 125440 671310 125530 671550
rect 125770 671310 125860 671550
rect 126100 671310 126210 671550
rect 126450 671310 126540 671550
rect 126780 671310 126870 671550
rect 127110 671310 127200 671550
rect 127440 671310 127550 671550
rect 127790 671310 127880 671550
rect 128120 671310 128210 671550
rect 128450 671310 128540 671550
rect 128780 671310 128890 671550
rect 129130 671310 129220 671550
rect 129460 671310 129550 671550
rect 129790 671310 129880 671550
rect 130120 671310 130230 671550
rect 130470 671310 130560 671550
rect 130800 671310 130890 671550
rect 131130 671310 131220 671550
rect 131460 671310 131570 671550
rect 131810 671310 131900 671550
rect 132140 671310 132230 671550
rect 132470 671310 132560 671550
rect 132800 671310 132910 671550
rect 133150 671310 133570 671550
rect 133810 671310 133900 671550
rect 134140 671310 134230 671550
rect 134470 671310 134560 671550
rect 134800 671310 134910 671550
rect 135150 671310 135240 671550
rect 135480 671310 135570 671550
rect 135810 671310 135900 671550
rect 136140 671310 136250 671550
rect 136490 671310 136580 671550
rect 136820 671310 136910 671550
rect 137150 671310 137240 671550
rect 137480 671310 137590 671550
rect 137830 671310 137920 671550
rect 138160 671310 138250 671550
rect 138490 671310 138580 671550
rect 138820 671310 138930 671550
rect 139170 671310 139260 671550
rect 139500 671310 139590 671550
rect 139830 671310 139920 671550
rect 140160 671310 140270 671550
rect 140510 671310 140600 671550
rect 140840 671310 140930 671550
rect 141170 671310 141260 671550
rect 141500 671310 141610 671550
rect 141850 671310 141940 671550
rect 142180 671310 142270 671550
rect 142510 671310 142600 671550
rect 142840 671310 142950 671550
rect 143190 671310 143280 671550
rect 143520 671310 143610 671550
rect 143850 671310 143940 671550
rect 144180 671310 144290 671550
rect 144530 671310 144950 671550
rect 145190 671310 145280 671550
rect 145520 671310 145610 671550
rect 145850 671310 145940 671550
rect 146180 671310 146290 671550
rect 146530 671310 146620 671550
rect 146860 671310 146950 671550
rect 147190 671310 147280 671550
rect 147520 671310 147630 671550
rect 147870 671310 147960 671550
rect 148200 671310 148290 671550
rect 148530 671310 148620 671550
rect 148860 671310 148970 671550
rect 149210 671310 149300 671550
rect 149540 671310 149630 671550
rect 149870 671310 149960 671550
rect 150200 671310 150310 671550
rect 150550 671310 150640 671550
rect 150880 671310 150970 671550
rect 151210 671310 151300 671550
rect 151540 671310 151650 671550
rect 151890 671310 151980 671550
rect 152220 671310 152310 671550
rect 152550 671310 152640 671550
rect 152880 671310 152990 671550
rect 153230 671310 153320 671550
rect 153560 671310 153650 671550
rect 153890 671310 153980 671550
rect 154220 671310 154330 671550
rect 154570 671310 154660 671550
rect 154900 671310 154990 671550
rect 155230 671310 155320 671550
rect 155560 671310 155670 671550
rect 155910 671310 155960 671550
rect 110760 671220 155960 671310
rect 110760 670980 110810 671220
rect 111050 670980 111140 671220
rect 111380 670980 111470 671220
rect 111710 670980 111800 671220
rect 112040 670980 112150 671220
rect 112390 670980 112480 671220
rect 112720 670980 112810 671220
rect 113050 670980 113140 671220
rect 113380 670980 113490 671220
rect 113730 670980 113820 671220
rect 114060 670980 114150 671220
rect 114390 670980 114480 671220
rect 114720 670980 114830 671220
rect 115070 670980 115160 671220
rect 115400 670980 115490 671220
rect 115730 670980 115820 671220
rect 116060 670980 116170 671220
rect 116410 670980 116500 671220
rect 116740 670980 116830 671220
rect 117070 670980 117160 671220
rect 117400 670980 117510 671220
rect 117750 670980 117840 671220
rect 118080 670980 118170 671220
rect 118410 670980 118500 671220
rect 118740 670980 118850 671220
rect 119090 670980 119180 671220
rect 119420 670980 119510 671220
rect 119750 670980 119840 671220
rect 120080 670980 120190 671220
rect 120430 670980 120520 671220
rect 120760 670980 120850 671220
rect 121090 670980 121180 671220
rect 121420 670980 121530 671220
rect 121770 670980 122190 671220
rect 122430 670980 122520 671220
rect 122760 670980 122850 671220
rect 123090 670980 123180 671220
rect 123420 670980 123530 671220
rect 123770 670980 123860 671220
rect 124100 670980 124190 671220
rect 124430 670980 124520 671220
rect 124760 670980 124870 671220
rect 125110 670980 125200 671220
rect 125440 670980 125530 671220
rect 125770 670980 125860 671220
rect 126100 670980 126210 671220
rect 126450 670980 126540 671220
rect 126780 670980 126870 671220
rect 127110 670980 127200 671220
rect 127440 670980 127550 671220
rect 127790 670980 127880 671220
rect 128120 670980 128210 671220
rect 128450 670980 128540 671220
rect 128780 670980 128890 671220
rect 129130 670980 129220 671220
rect 129460 670980 129550 671220
rect 129790 670980 129880 671220
rect 130120 670980 130230 671220
rect 130470 670980 130560 671220
rect 130800 670980 130890 671220
rect 131130 670980 131220 671220
rect 131460 670980 131570 671220
rect 131810 670980 131900 671220
rect 132140 670980 132230 671220
rect 132470 670980 132560 671220
rect 132800 670980 132910 671220
rect 133150 670980 133570 671220
rect 133810 670980 133900 671220
rect 134140 670980 134230 671220
rect 134470 670980 134560 671220
rect 134800 670980 134910 671220
rect 135150 670980 135240 671220
rect 135480 670980 135570 671220
rect 135810 670980 135900 671220
rect 136140 670980 136250 671220
rect 136490 670980 136580 671220
rect 136820 670980 136910 671220
rect 137150 670980 137240 671220
rect 137480 670980 137590 671220
rect 137830 670980 137920 671220
rect 138160 670980 138250 671220
rect 138490 670980 138580 671220
rect 138820 670980 138930 671220
rect 139170 670980 139260 671220
rect 139500 670980 139590 671220
rect 139830 670980 139920 671220
rect 140160 670980 140270 671220
rect 140510 670980 140600 671220
rect 140840 670980 140930 671220
rect 141170 670980 141260 671220
rect 141500 670980 141610 671220
rect 141850 670980 141940 671220
rect 142180 670980 142270 671220
rect 142510 670980 142600 671220
rect 142840 670980 142950 671220
rect 143190 670980 143280 671220
rect 143520 670980 143610 671220
rect 143850 670980 143940 671220
rect 144180 670980 144290 671220
rect 144530 670980 144950 671220
rect 145190 670980 145280 671220
rect 145520 670980 145610 671220
rect 145850 670980 145940 671220
rect 146180 670980 146290 671220
rect 146530 670980 146620 671220
rect 146860 670980 146950 671220
rect 147190 670980 147280 671220
rect 147520 670980 147630 671220
rect 147870 670980 147960 671220
rect 148200 670980 148290 671220
rect 148530 670980 148620 671220
rect 148860 670980 148970 671220
rect 149210 670980 149300 671220
rect 149540 670980 149630 671220
rect 149870 670980 149960 671220
rect 150200 670980 150310 671220
rect 150550 670980 150640 671220
rect 150880 670980 150970 671220
rect 151210 670980 151300 671220
rect 151540 670980 151650 671220
rect 151890 670980 151980 671220
rect 152220 670980 152310 671220
rect 152550 670980 152640 671220
rect 152880 670980 152990 671220
rect 153230 670980 153320 671220
rect 153560 670980 153650 671220
rect 153890 670980 153980 671220
rect 154220 670980 154330 671220
rect 154570 670980 154660 671220
rect 154900 670980 154990 671220
rect 155230 670980 155320 671220
rect 155560 670980 155670 671220
rect 155910 670980 155960 671220
rect 110760 670890 155960 670980
rect 110760 670650 110810 670890
rect 111050 670650 111140 670890
rect 111380 670650 111470 670890
rect 111710 670650 111800 670890
rect 112040 670650 112150 670890
rect 112390 670650 112480 670890
rect 112720 670650 112810 670890
rect 113050 670650 113140 670890
rect 113380 670650 113490 670890
rect 113730 670650 113820 670890
rect 114060 670650 114150 670890
rect 114390 670650 114480 670890
rect 114720 670650 114830 670890
rect 115070 670650 115160 670890
rect 115400 670650 115490 670890
rect 115730 670650 115820 670890
rect 116060 670650 116170 670890
rect 116410 670650 116500 670890
rect 116740 670650 116830 670890
rect 117070 670650 117160 670890
rect 117400 670650 117510 670890
rect 117750 670650 117840 670890
rect 118080 670650 118170 670890
rect 118410 670650 118500 670890
rect 118740 670650 118850 670890
rect 119090 670650 119180 670890
rect 119420 670650 119510 670890
rect 119750 670650 119840 670890
rect 120080 670650 120190 670890
rect 120430 670650 120520 670890
rect 120760 670650 120850 670890
rect 121090 670650 121180 670890
rect 121420 670650 121530 670890
rect 121770 670650 122190 670890
rect 122430 670650 122520 670890
rect 122760 670650 122850 670890
rect 123090 670650 123180 670890
rect 123420 670650 123530 670890
rect 123770 670650 123860 670890
rect 124100 670650 124190 670890
rect 124430 670650 124520 670890
rect 124760 670650 124870 670890
rect 125110 670650 125200 670890
rect 125440 670650 125530 670890
rect 125770 670650 125860 670890
rect 126100 670650 126210 670890
rect 126450 670650 126540 670890
rect 126780 670650 126870 670890
rect 127110 670650 127200 670890
rect 127440 670650 127550 670890
rect 127790 670650 127880 670890
rect 128120 670650 128210 670890
rect 128450 670650 128540 670890
rect 128780 670650 128890 670890
rect 129130 670650 129220 670890
rect 129460 670650 129550 670890
rect 129790 670650 129880 670890
rect 130120 670650 130230 670890
rect 130470 670650 130560 670890
rect 130800 670650 130890 670890
rect 131130 670650 131220 670890
rect 131460 670650 131570 670890
rect 131810 670650 131900 670890
rect 132140 670650 132230 670890
rect 132470 670650 132560 670890
rect 132800 670650 132910 670890
rect 133150 670650 133570 670890
rect 133810 670650 133900 670890
rect 134140 670650 134230 670890
rect 134470 670650 134560 670890
rect 134800 670650 134910 670890
rect 135150 670650 135240 670890
rect 135480 670650 135570 670890
rect 135810 670650 135900 670890
rect 136140 670650 136250 670890
rect 136490 670650 136580 670890
rect 136820 670650 136910 670890
rect 137150 670650 137240 670890
rect 137480 670650 137590 670890
rect 137830 670650 137920 670890
rect 138160 670650 138250 670890
rect 138490 670650 138580 670890
rect 138820 670650 138930 670890
rect 139170 670650 139260 670890
rect 139500 670650 139590 670890
rect 139830 670650 139920 670890
rect 140160 670650 140270 670890
rect 140510 670650 140600 670890
rect 140840 670650 140930 670890
rect 141170 670650 141260 670890
rect 141500 670650 141610 670890
rect 141850 670650 141940 670890
rect 142180 670650 142270 670890
rect 142510 670650 142600 670890
rect 142840 670650 142950 670890
rect 143190 670650 143280 670890
rect 143520 670650 143610 670890
rect 143850 670650 143940 670890
rect 144180 670650 144290 670890
rect 144530 670650 144950 670890
rect 145190 670650 145280 670890
rect 145520 670650 145610 670890
rect 145850 670650 145940 670890
rect 146180 670650 146290 670890
rect 146530 670650 146620 670890
rect 146860 670650 146950 670890
rect 147190 670650 147280 670890
rect 147520 670650 147630 670890
rect 147870 670650 147960 670890
rect 148200 670650 148290 670890
rect 148530 670650 148620 670890
rect 148860 670650 148970 670890
rect 149210 670650 149300 670890
rect 149540 670650 149630 670890
rect 149870 670650 149960 670890
rect 150200 670650 150310 670890
rect 150550 670650 150640 670890
rect 150880 670650 150970 670890
rect 151210 670650 151300 670890
rect 151540 670650 151650 670890
rect 151890 670650 151980 670890
rect 152220 670650 152310 670890
rect 152550 670650 152640 670890
rect 152880 670650 152990 670890
rect 153230 670650 153320 670890
rect 153560 670650 153650 670890
rect 153890 670650 153980 670890
rect 154220 670650 154330 670890
rect 154570 670650 154660 670890
rect 154900 670650 154990 670890
rect 155230 670650 155320 670890
rect 155560 670650 155670 670890
rect 155910 670650 155960 670890
rect 110760 670560 155960 670650
rect 110760 670320 110810 670560
rect 111050 670320 111140 670560
rect 111380 670320 111470 670560
rect 111710 670320 111800 670560
rect 112040 670320 112150 670560
rect 112390 670320 112480 670560
rect 112720 670320 112810 670560
rect 113050 670320 113140 670560
rect 113380 670320 113490 670560
rect 113730 670320 113820 670560
rect 114060 670320 114150 670560
rect 114390 670320 114480 670560
rect 114720 670320 114830 670560
rect 115070 670320 115160 670560
rect 115400 670320 115490 670560
rect 115730 670320 115820 670560
rect 116060 670320 116170 670560
rect 116410 670320 116500 670560
rect 116740 670320 116830 670560
rect 117070 670320 117160 670560
rect 117400 670320 117510 670560
rect 117750 670320 117840 670560
rect 118080 670320 118170 670560
rect 118410 670320 118500 670560
rect 118740 670320 118850 670560
rect 119090 670320 119180 670560
rect 119420 670320 119510 670560
rect 119750 670320 119840 670560
rect 120080 670320 120190 670560
rect 120430 670320 120520 670560
rect 120760 670320 120850 670560
rect 121090 670320 121180 670560
rect 121420 670320 121530 670560
rect 121770 670320 122190 670560
rect 122430 670320 122520 670560
rect 122760 670320 122850 670560
rect 123090 670320 123180 670560
rect 123420 670320 123530 670560
rect 123770 670320 123860 670560
rect 124100 670320 124190 670560
rect 124430 670320 124520 670560
rect 124760 670320 124870 670560
rect 125110 670320 125200 670560
rect 125440 670320 125530 670560
rect 125770 670320 125860 670560
rect 126100 670320 126210 670560
rect 126450 670320 126540 670560
rect 126780 670320 126870 670560
rect 127110 670320 127200 670560
rect 127440 670320 127550 670560
rect 127790 670320 127880 670560
rect 128120 670320 128210 670560
rect 128450 670320 128540 670560
rect 128780 670320 128890 670560
rect 129130 670320 129220 670560
rect 129460 670320 129550 670560
rect 129790 670320 129880 670560
rect 130120 670320 130230 670560
rect 130470 670320 130560 670560
rect 130800 670320 130890 670560
rect 131130 670320 131220 670560
rect 131460 670320 131570 670560
rect 131810 670320 131900 670560
rect 132140 670320 132230 670560
rect 132470 670320 132560 670560
rect 132800 670320 132910 670560
rect 133150 670320 133570 670560
rect 133810 670320 133900 670560
rect 134140 670320 134230 670560
rect 134470 670320 134560 670560
rect 134800 670320 134910 670560
rect 135150 670320 135240 670560
rect 135480 670320 135570 670560
rect 135810 670320 135900 670560
rect 136140 670320 136250 670560
rect 136490 670320 136580 670560
rect 136820 670320 136910 670560
rect 137150 670320 137240 670560
rect 137480 670320 137590 670560
rect 137830 670320 137920 670560
rect 138160 670320 138250 670560
rect 138490 670320 138580 670560
rect 138820 670320 138930 670560
rect 139170 670320 139260 670560
rect 139500 670320 139590 670560
rect 139830 670320 139920 670560
rect 140160 670320 140270 670560
rect 140510 670320 140600 670560
rect 140840 670320 140930 670560
rect 141170 670320 141260 670560
rect 141500 670320 141610 670560
rect 141850 670320 141940 670560
rect 142180 670320 142270 670560
rect 142510 670320 142600 670560
rect 142840 670320 142950 670560
rect 143190 670320 143280 670560
rect 143520 670320 143610 670560
rect 143850 670320 143940 670560
rect 144180 670320 144290 670560
rect 144530 670320 144950 670560
rect 145190 670320 145280 670560
rect 145520 670320 145610 670560
rect 145850 670320 145940 670560
rect 146180 670320 146290 670560
rect 146530 670320 146620 670560
rect 146860 670320 146950 670560
rect 147190 670320 147280 670560
rect 147520 670320 147630 670560
rect 147870 670320 147960 670560
rect 148200 670320 148290 670560
rect 148530 670320 148620 670560
rect 148860 670320 148970 670560
rect 149210 670320 149300 670560
rect 149540 670320 149630 670560
rect 149870 670320 149960 670560
rect 150200 670320 150310 670560
rect 150550 670320 150640 670560
rect 150880 670320 150970 670560
rect 151210 670320 151300 670560
rect 151540 670320 151650 670560
rect 151890 670320 151980 670560
rect 152220 670320 152310 670560
rect 152550 670320 152640 670560
rect 152880 670320 152990 670560
rect 153230 670320 153320 670560
rect 153560 670320 153650 670560
rect 153890 670320 153980 670560
rect 154220 670320 154330 670560
rect 154570 670320 154660 670560
rect 154900 670320 154990 670560
rect 155230 670320 155320 670560
rect 155560 670320 155670 670560
rect 155910 670320 155960 670560
rect 110760 670210 155960 670320
rect 110760 669970 110810 670210
rect 111050 669970 111140 670210
rect 111380 669970 111470 670210
rect 111710 669970 111800 670210
rect 112040 669970 112150 670210
rect 112390 669970 112480 670210
rect 112720 669970 112810 670210
rect 113050 669970 113140 670210
rect 113380 669970 113490 670210
rect 113730 669970 113820 670210
rect 114060 669970 114150 670210
rect 114390 669970 114480 670210
rect 114720 669970 114830 670210
rect 115070 669970 115160 670210
rect 115400 669970 115490 670210
rect 115730 669970 115820 670210
rect 116060 669970 116170 670210
rect 116410 669970 116500 670210
rect 116740 669970 116830 670210
rect 117070 669970 117160 670210
rect 117400 669970 117510 670210
rect 117750 669970 117840 670210
rect 118080 669970 118170 670210
rect 118410 669970 118500 670210
rect 118740 669970 118850 670210
rect 119090 669970 119180 670210
rect 119420 669970 119510 670210
rect 119750 669970 119840 670210
rect 120080 669970 120190 670210
rect 120430 669970 120520 670210
rect 120760 669970 120850 670210
rect 121090 669970 121180 670210
rect 121420 669970 121530 670210
rect 121770 669970 122190 670210
rect 122430 669970 122520 670210
rect 122760 669970 122850 670210
rect 123090 669970 123180 670210
rect 123420 669970 123530 670210
rect 123770 669970 123860 670210
rect 124100 669970 124190 670210
rect 124430 669970 124520 670210
rect 124760 669970 124870 670210
rect 125110 669970 125200 670210
rect 125440 669970 125530 670210
rect 125770 669970 125860 670210
rect 126100 669970 126210 670210
rect 126450 669970 126540 670210
rect 126780 669970 126870 670210
rect 127110 669970 127200 670210
rect 127440 669970 127550 670210
rect 127790 669970 127880 670210
rect 128120 669970 128210 670210
rect 128450 669970 128540 670210
rect 128780 669970 128890 670210
rect 129130 669970 129220 670210
rect 129460 669970 129550 670210
rect 129790 669970 129880 670210
rect 130120 669970 130230 670210
rect 130470 669970 130560 670210
rect 130800 669970 130890 670210
rect 131130 669970 131220 670210
rect 131460 669970 131570 670210
rect 131810 669970 131900 670210
rect 132140 669970 132230 670210
rect 132470 669970 132560 670210
rect 132800 669970 132910 670210
rect 133150 669970 133570 670210
rect 133810 669970 133900 670210
rect 134140 669970 134230 670210
rect 134470 669970 134560 670210
rect 134800 669970 134910 670210
rect 135150 669970 135240 670210
rect 135480 669970 135570 670210
rect 135810 669970 135900 670210
rect 136140 669970 136250 670210
rect 136490 669970 136580 670210
rect 136820 669970 136910 670210
rect 137150 669970 137240 670210
rect 137480 669970 137590 670210
rect 137830 669970 137920 670210
rect 138160 669970 138250 670210
rect 138490 669970 138580 670210
rect 138820 669970 138930 670210
rect 139170 669970 139260 670210
rect 139500 669970 139590 670210
rect 139830 669970 139920 670210
rect 140160 669970 140270 670210
rect 140510 669970 140600 670210
rect 140840 669970 140930 670210
rect 141170 669970 141260 670210
rect 141500 669970 141610 670210
rect 141850 669970 141940 670210
rect 142180 669970 142270 670210
rect 142510 669970 142600 670210
rect 142840 669970 142950 670210
rect 143190 669970 143280 670210
rect 143520 669970 143610 670210
rect 143850 669970 143940 670210
rect 144180 669970 144290 670210
rect 144530 669970 144950 670210
rect 145190 669970 145280 670210
rect 145520 669970 145610 670210
rect 145850 669970 145940 670210
rect 146180 669970 146290 670210
rect 146530 669970 146620 670210
rect 146860 669970 146950 670210
rect 147190 669970 147280 670210
rect 147520 669970 147630 670210
rect 147870 669970 147960 670210
rect 148200 669970 148290 670210
rect 148530 669970 148620 670210
rect 148860 669970 148970 670210
rect 149210 669970 149300 670210
rect 149540 669970 149630 670210
rect 149870 669970 149960 670210
rect 150200 669970 150310 670210
rect 150550 669970 150640 670210
rect 150880 669970 150970 670210
rect 151210 669970 151300 670210
rect 151540 669970 151650 670210
rect 151890 669970 151980 670210
rect 152220 669970 152310 670210
rect 152550 669970 152640 670210
rect 152880 669970 152990 670210
rect 153230 669970 153320 670210
rect 153560 669970 153650 670210
rect 153890 669970 153980 670210
rect 154220 669970 154330 670210
rect 154570 669970 154660 670210
rect 154900 669970 154990 670210
rect 155230 669970 155320 670210
rect 155560 669970 155670 670210
rect 155910 669970 155960 670210
rect 110760 669880 155960 669970
rect 110760 669640 110810 669880
rect 111050 669640 111140 669880
rect 111380 669640 111470 669880
rect 111710 669640 111800 669880
rect 112040 669640 112150 669880
rect 112390 669640 112480 669880
rect 112720 669640 112810 669880
rect 113050 669640 113140 669880
rect 113380 669640 113490 669880
rect 113730 669640 113820 669880
rect 114060 669640 114150 669880
rect 114390 669640 114480 669880
rect 114720 669640 114830 669880
rect 115070 669640 115160 669880
rect 115400 669640 115490 669880
rect 115730 669640 115820 669880
rect 116060 669640 116170 669880
rect 116410 669640 116500 669880
rect 116740 669640 116830 669880
rect 117070 669640 117160 669880
rect 117400 669640 117510 669880
rect 117750 669640 117840 669880
rect 118080 669640 118170 669880
rect 118410 669640 118500 669880
rect 118740 669640 118850 669880
rect 119090 669640 119180 669880
rect 119420 669640 119510 669880
rect 119750 669640 119840 669880
rect 120080 669640 120190 669880
rect 120430 669640 120520 669880
rect 120760 669640 120850 669880
rect 121090 669640 121180 669880
rect 121420 669640 121530 669880
rect 121770 669640 122190 669880
rect 122430 669640 122520 669880
rect 122760 669640 122850 669880
rect 123090 669640 123180 669880
rect 123420 669640 123530 669880
rect 123770 669640 123860 669880
rect 124100 669640 124190 669880
rect 124430 669640 124520 669880
rect 124760 669640 124870 669880
rect 125110 669640 125200 669880
rect 125440 669640 125530 669880
rect 125770 669640 125860 669880
rect 126100 669640 126210 669880
rect 126450 669640 126540 669880
rect 126780 669640 126870 669880
rect 127110 669640 127200 669880
rect 127440 669640 127550 669880
rect 127790 669640 127880 669880
rect 128120 669640 128210 669880
rect 128450 669640 128540 669880
rect 128780 669640 128890 669880
rect 129130 669640 129220 669880
rect 129460 669640 129550 669880
rect 129790 669640 129880 669880
rect 130120 669640 130230 669880
rect 130470 669640 130560 669880
rect 130800 669640 130890 669880
rect 131130 669640 131220 669880
rect 131460 669640 131570 669880
rect 131810 669640 131900 669880
rect 132140 669640 132230 669880
rect 132470 669640 132560 669880
rect 132800 669640 132910 669880
rect 133150 669640 133570 669880
rect 133810 669640 133900 669880
rect 134140 669640 134230 669880
rect 134470 669640 134560 669880
rect 134800 669640 134910 669880
rect 135150 669640 135240 669880
rect 135480 669640 135570 669880
rect 135810 669640 135900 669880
rect 136140 669640 136250 669880
rect 136490 669640 136580 669880
rect 136820 669640 136910 669880
rect 137150 669640 137240 669880
rect 137480 669640 137590 669880
rect 137830 669640 137920 669880
rect 138160 669640 138250 669880
rect 138490 669640 138580 669880
rect 138820 669640 138930 669880
rect 139170 669640 139260 669880
rect 139500 669640 139590 669880
rect 139830 669640 139920 669880
rect 140160 669640 140270 669880
rect 140510 669640 140600 669880
rect 140840 669640 140930 669880
rect 141170 669640 141260 669880
rect 141500 669640 141610 669880
rect 141850 669640 141940 669880
rect 142180 669640 142270 669880
rect 142510 669640 142600 669880
rect 142840 669640 142950 669880
rect 143190 669640 143280 669880
rect 143520 669640 143610 669880
rect 143850 669640 143940 669880
rect 144180 669640 144290 669880
rect 144530 669640 144950 669880
rect 145190 669640 145280 669880
rect 145520 669640 145610 669880
rect 145850 669640 145940 669880
rect 146180 669640 146290 669880
rect 146530 669640 146620 669880
rect 146860 669640 146950 669880
rect 147190 669640 147280 669880
rect 147520 669640 147630 669880
rect 147870 669640 147960 669880
rect 148200 669640 148290 669880
rect 148530 669640 148620 669880
rect 148860 669640 148970 669880
rect 149210 669640 149300 669880
rect 149540 669640 149630 669880
rect 149870 669640 149960 669880
rect 150200 669640 150310 669880
rect 150550 669640 150640 669880
rect 150880 669640 150970 669880
rect 151210 669640 151300 669880
rect 151540 669640 151650 669880
rect 151890 669640 151980 669880
rect 152220 669640 152310 669880
rect 152550 669640 152640 669880
rect 152880 669640 152990 669880
rect 153230 669640 153320 669880
rect 153560 669640 153650 669880
rect 153890 669640 153980 669880
rect 154220 669640 154330 669880
rect 154570 669640 154660 669880
rect 154900 669640 154990 669880
rect 155230 669640 155320 669880
rect 155560 669640 155670 669880
rect 155910 669640 155960 669880
rect 110760 669550 155960 669640
rect 110760 669310 110810 669550
rect 111050 669310 111140 669550
rect 111380 669310 111470 669550
rect 111710 669310 111800 669550
rect 112040 669310 112150 669550
rect 112390 669310 112480 669550
rect 112720 669310 112810 669550
rect 113050 669310 113140 669550
rect 113380 669310 113490 669550
rect 113730 669310 113820 669550
rect 114060 669310 114150 669550
rect 114390 669310 114480 669550
rect 114720 669310 114830 669550
rect 115070 669310 115160 669550
rect 115400 669310 115490 669550
rect 115730 669310 115820 669550
rect 116060 669310 116170 669550
rect 116410 669310 116500 669550
rect 116740 669310 116830 669550
rect 117070 669310 117160 669550
rect 117400 669310 117510 669550
rect 117750 669310 117840 669550
rect 118080 669310 118170 669550
rect 118410 669310 118500 669550
rect 118740 669310 118850 669550
rect 119090 669310 119180 669550
rect 119420 669310 119510 669550
rect 119750 669310 119840 669550
rect 120080 669310 120190 669550
rect 120430 669310 120520 669550
rect 120760 669310 120850 669550
rect 121090 669310 121180 669550
rect 121420 669310 121530 669550
rect 121770 669310 122190 669550
rect 122430 669310 122520 669550
rect 122760 669310 122850 669550
rect 123090 669310 123180 669550
rect 123420 669310 123530 669550
rect 123770 669310 123860 669550
rect 124100 669310 124190 669550
rect 124430 669310 124520 669550
rect 124760 669310 124870 669550
rect 125110 669310 125200 669550
rect 125440 669310 125530 669550
rect 125770 669310 125860 669550
rect 126100 669310 126210 669550
rect 126450 669310 126540 669550
rect 126780 669310 126870 669550
rect 127110 669310 127200 669550
rect 127440 669310 127550 669550
rect 127790 669310 127880 669550
rect 128120 669310 128210 669550
rect 128450 669310 128540 669550
rect 128780 669310 128890 669550
rect 129130 669310 129220 669550
rect 129460 669310 129550 669550
rect 129790 669310 129880 669550
rect 130120 669310 130230 669550
rect 130470 669310 130560 669550
rect 130800 669310 130890 669550
rect 131130 669310 131220 669550
rect 131460 669310 131570 669550
rect 131810 669310 131900 669550
rect 132140 669310 132230 669550
rect 132470 669310 132560 669550
rect 132800 669310 132910 669550
rect 133150 669310 133570 669550
rect 133810 669310 133900 669550
rect 134140 669310 134230 669550
rect 134470 669310 134560 669550
rect 134800 669310 134910 669550
rect 135150 669310 135240 669550
rect 135480 669310 135570 669550
rect 135810 669310 135900 669550
rect 136140 669310 136250 669550
rect 136490 669310 136580 669550
rect 136820 669310 136910 669550
rect 137150 669310 137240 669550
rect 137480 669310 137590 669550
rect 137830 669310 137920 669550
rect 138160 669310 138250 669550
rect 138490 669310 138580 669550
rect 138820 669310 138930 669550
rect 139170 669310 139260 669550
rect 139500 669310 139590 669550
rect 139830 669310 139920 669550
rect 140160 669310 140270 669550
rect 140510 669310 140600 669550
rect 140840 669310 140930 669550
rect 141170 669310 141260 669550
rect 141500 669310 141610 669550
rect 141850 669310 141940 669550
rect 142180 669310 142270 669550
rect 142510 669310 142600 669550
rect 142840 669310 142950 669550
rect 143190 669310 143280 669550
rect 143520 669310 143610 669550
rect 143850 669310 143940 669550
rect 144180 669310 144290 669550
rect 144530 669310 144950 669550
rect 145190 669310 145280 669550
rect 145520 669310 145610 669550
rect 145850 669310 145940 669550
rect 146180 669310 146290 669550
rect 146530 669310 146620 669550
rect 146860 669310 146950 669550
rect 147190 669310 147280 669550
rect 147520 669310 147630 669550
rect 147870 669310 147960 669550
rect 148200 669310 148290 669550
rect 148530 669310 148620 669550
rect 148860 669310 148970 669550
rect 149210 669310 149300 669550
rect 149540 669310 149630 669550
rect 149870 669310 149960 669550
rect 150200 669310 150310 669550
rect 150550 669310 150640 669550
rect 150880 669310 150970 669550
rect 151210 669310 151300 669550
rect 151540 669310 151650 669550
rect 151890 669310 151980 669550
rect 152220 669310 152310 669550
rect 152550 669310 152640 669550
rect 152880 669310 152990 669550
rect 153230 669310 153320 669550
rect 153560 669310 153650 669550
rect 153890 669310 153980 669550
rect 154220 669310 154330 669550
rect 154570 669310 154660 669550
rect 154900 669310 154990 669550
rect 155230 669310 155320 669550
rect 155560 669310 155670 669550
rect 155910 669310 155960 669550
rect 110760 669220 155960 669310
rect 110760 668980 110810 669220
rect 111050 668980 111140 669220
rect 111380 668980 111470 669220
rect 111710 668980 111800 669220
rect 112040 668980 112150 669220
rect 112390 668980 112480 669220
rect 112720 668980 112810 669220
rect 113050 668980 113140 669220
rect 113380 668980 113490 669220
rect 113730 668980 113820 669220
rect 114060 668980 114150 669220
rect 114390 668980 114480 669220
rect 114720 668980 114830 669220
rect 115070 668980 115160 669220
rect 115400 668980 115490 669220
rect 115730 668980 115820 669220
rect 116060 668980 116170 669220
rect 116410 668980 116500 669220
rect 116740 668980 116830 669220
rect 117070 668980 117160 669220
rect 117400 668980 117510 669220
rect 117750 668980 117840 669220
rect 118080 668980 118170 669220
rect 118410 668980 118500 669220
rect 118740 668980 118850 669220
rect 119090 668980 119180 669220
rect 119420 668980 119510 669220
rect 119750 668980 119840 669220
rect 120080 668980 120190 669220
rect 120430 668980 120520 669220
rect 120760 668980 120850 669220
rect 121090 668980 121180 669220
rect 121420 668980 121530 669220
rect 121770 668980 122190 669220
rect 122430 668980 122520 669220
rect 122760 668980 122850 669220
rect 123090 668980 123180 669220
rect 123420 668980 123530 669220
rect 123770 668980 123860 669220
rect 124100 668980 124190 669220
rect 124430 668980 124520 669220
rect 124760 668980 124870 669220
rect 125110 668980 125200 669220
rect 125440 668980 125530 669220
rect 125770 668980 125860 669220
rect 126100 668980 126210 669220
rect 126450 668980 126540 669220
rect 126780 668980 126870 669220
rect 127110 668980 127200 669220
rect 127440 668980 127550 669220
rect 127790 668980 127880 669220
rect 128120 668980 128210 669220
rect 128450 668980 128540 669220
rect 128780 668980 128890 669220
rect 129130 668980 129220 669220
rect 129460 668980 129550 669220
rect 129790 668980 129880 669220
rect 130120 668980 130230 669220
rect 130470 668980 130560 669220
rect 130800 668980 130890 669220
rect 131130 668980 131220 669220
rect 131460 668980 131570 669220
rect 131810 668980 131900 669220
rect 132140 668980 132230 669220
rect 132470 668980 132560 669220
rect 132800 668980 132910 669220
rect 133150 668980 133570 669220
rect 133810 668980 133900 669220
rect 134140 668980 134230 669220
rect 134470 668980 134560 669220
rect 134800 668980 134910 669220
rect 135150 668980 135240 669220
rect 135480 668980 135570 669220
rect 135810 668980 135900 669220
rect 136140 668980 136250 669220
rect 136490 668980 136580 669220
rect 136820 668980 136910 669220
rect 137150 668980 137240 669220
rect 137480 668980 137590 669220
rect 137830 668980 137920 669220
rect 138160 668980 138250 669220
rect 138490 668980 138580 669220
rect 138820 668980 138930 669220
rect 139170 668980 139260 669220
rect 139500 668980 139590 669220
rect 139830 668980 139920 669220
rect 140160 668980 140270 669220
rect 140510 668980 140600 669220
rect 140840 668980 140930 669220
rect 141170 668980 141260 669220
rect 141500 668980 141610 669220
rect 141850 668980 141940 669220
rect 142180 668980 142270 669220
rect 142510 668980 142600 669220
rect 142840 668980 142950 669220
rect 143190 668980 143280 669220
rect 143520 668980 143610 669220
rect 143850 668980 143940 669220
rect 144180 668980 144290 669220
rect 144530 668980 144950 669220
rect 145190 668980 145280 669220
rect 145520 668980 145610 669220
rect 145850 668980 145940 669220
rect 146180 668980 146290 669220
rect 146530 668980 146620 669220
rect 146860 668980 146950 669220
rect 147190 668980 147280 669220
rect 147520 668980 147630 669220
rect 147870 668980 147960 669220
rect 148200 668980 148290 669220
rect 148530 668980 148620 669220
rect 148860 668980 148970 669220
rect 149210 668980 149300 669220
rect 149540 668980 149630 669220
rect 149870 668980 149960 669220
rect 150200 668980 150310 669220
rect 150550 668980 150640 669220
rect 150880 668980 150970 669220
rect 151210 668980 151300 669220
rect 151540 668980 151650 669220
rect 151890 668980 151980 669220
rect 152220 668980 152310 669220
rect 152550 668980 152640 669220
rect 152880 668980 152990 669220
rect 153230 668980 153320 669220
rect 153560 668980 153650 669220
rect 153890 668980 153980 669220
rect 154220 668980 154330 669220
rect 154570 668980 154660 669220
rect 154900 668980 154990 669220
rect 155230 668980 155320 669220
rect 155560 668980 155670 669220
rect 155910 668980 155960 669220
rect 110760 668870 155960 668980
rect 110760 668630 110810 668870
rect 111050 668630 111140 668870
rect 111380 668630 111470 668870
rect 111710 668630 111800 668870
rect 112040 668630 112150 668870
rect 112390 668630 112480 668870
rect 112720 668630 112810 668870
rect 113050 668630 113140 668870
rect 113380 668630 113490 668870
rect 113730 668630 113820 668870
rect 114060 668630 114150 668870
rect 114390 668630 114480 668870
rect 114720 668630 114830 668870
rect 115070 668630 115160 668870
rect 115400 668630 115490 668870
rect 115730 668630 115820 668870
rect 116060 668630 116170 668870
rect 116410 668630 116500 668870
rect 116740 668630 116830 668870
rect 117070 668630 117160 668870
rect 117400 668630 117510 668870
rect 117750 668630 117840 668870
rect 118080 668630 118170 668870
rect 118410 668630 118500 668870
rect 118740 668630 118850 668870
rect 119090 668630 119180 668870
rect 119420 668630 119510 668870
rect 119750 668630 119840 668870
rect 120080 668630 120190 668870
rect 120430 668630 120520 668870
rect 120760 668630 120850 668870
rect 121090 668630 121180 668870
rect 121420 668630 121530 668870
rect 121770 668630 122190 668870
rect 122430 668630 122520 668870
rect 122760 668630 122850 668870
rect 123090 668630 123180 668870
rect 123420 668630 123530 668870
rect 123770 668630 123860 668870
rect 124100 668630 124190 668870
rect 124430 668630 124520 668870
rect 124760 668630 124870 668870
rect 125110 668630 125200 668870
rect 125440 668630 125530 668870
rect 125770 668630 125860 668870
rect 126100 668630 126210 668870
rect 126450 668630 126540 668870
rect 126780 668630 126870 668870
rect 127110 668630 127200 668870
rect 127440 668630 127550 668870
rect 127790 668630 127880 668870
rect 128120 668630 128210 668870
rect 128450 668630 128540 668870
rect 128780 668630 128890 668870
rect 129130 668630 129220 668870
rect 129460 668630 129550 668870
rect 129790 668630 129880 668870
rect 130120 668630 130230 668870
rect 130470 668630 130560 668870
rect 130800 668630 130890 668870
rect 131130 668630 131220 668870
rect 131460 668630 131570 668870
rect 131810 668630 131900 668870
rect 132140 668630 132230 668870
rect 132470 668630 132560 668870
rect 132800 668630 132910 668870
rect 133150 668630 133570 668870
rect 133810 668630 133900 668870
rect 134140 668630 134230 668870
rect 134470 668630 134560 668870
rect 134800 668630 134910 668870
rect 135150 668630 135240 668870
rect 135480 668630 135570 668870
rect 135810 668630 135900 668870
rect 136140 668630 136250 668870
rect 136490 668630 136580 668870
rect 136820 668630 136910 668870
rect 137150 668630 137240 668870
rect 137480 668630 137590 668870
rect 137830 668630 137920 668870
rect 138160 668630 138250 668870
rect 138490 668630 138580 668870
rect 138820 668630 138930 668870
rect 139170 668630 139260 668870
rect 139500 668630 139590 668870
rect 139830 668630 139920 668870
rect 140160 668630 140270 668870
rect 140510 668630 140600 668870
rect 140840 668630 140930 668870
rect 141170 668630 141260 668870
rect 141500 668630 141610 668870
rect 141850 668630 141940 668870
rect 142180 668630 142270 668870
rect 142510 668630 142600 668870
rect 142840 668630 142950 668870
rect 143190 668630 143280 668870
rect 143520 668630 143610 668870
rect 143850 668630 143940 668870
rect 144180 668630 144290 668870
rect 144530 668630 144950 668870
rect 145190 668630 145280 668870
rect 145520 668630 145610 668870
rect 145850 668630 145940 668870
rect 146180 668630 146290 668870
rect 146530 668630 146620 668870
rect 146860 668630 146950 668870
rect 147190 668630 147280 668870
rect 147520 668630 147630 668870
rect 147870 668630 147960 668870
rect 148200 668630 148290 668870
rect 148530 668630 148620 668870
rect 148860 668630 148970 668870
rect 149210 668630 149300 668870
rect 149540 668630 149630 668870
rect 149870 668630 149960 668870
rect 150200 668630 150310 668870
rect 150550 668630 150640 668870
rect 150880 668630 150970 668870
rect 151210 668630 151300 668870
rect 151540 668630 151650 668870
rect 151890 668630 151980 668870
rect 152220 668630 152310 668870
rect 152550 668630 152640 668870
rect 152880 668630 152990 668870
rect 153230 668630 153320 668870
rect 153560 668630 153650 668870
rect 153890 668630 153980 668870
rect 154220 668630 154330 668870
rect 154570 668630 154660 668870
rect 154900 668630 154990 668870
rect 155230 668630 155320 668870
rect 155560 668630 155670 668870
rect 155910 668630 155960 668870
rect 110760 668540 155960 668630
rect 110760 668300 110810 668540
rect 111050 668300 111140 668540
rect 111380 668300 111470 668540
rect 111710 668300 111800 668540
rect 112040 668300 112150 668540
rect 112390 668300 112480 668540
rect 112720 668300 112810 668540
rect 113050 668300 113140 668540
rect 113380 668300 113490 668540
rect 113730 668300 113820 668540
rect 114060 668300 114150 668540
rect 114390 668300 114480 668540
rect 114720 668300 114830 668540
rect 115070 668300 115160 668540
rect 115400 668300 115490 668540
rect 115730 668300 115820 668540
rect 116060 668300 116170 668540
rect 116410 668300 116500 668540
rect 116740 668300 116830 668540
rect 117070 668300 117160 668540
rect 117400 668300 117510 668540
rect 117750 668300 117840 668540
rect 118080 668300 118170 668540
rect 118410 668300 118500 668540
rect 118740 668300 118850 668540
rect 119090 668300 119180 668540
rect 119420 668300 119510 668540
rect 119750 668300 119840 668540
rect 120080 668300 120190 668540
rect 120430 668300 120520 668540
rect 120760 668300 120850 668540
rect 121090 668300 121180 668540
rect 121420 668300 121530 668540
rect 121770 668300 122190 668540
rect 122430 668300 122520 668540
rect 122760 668300 122850 668540
rect 123090 668300 123180 668540
rect 123420 668300 123530 668540
rect 123770 668300 123860 668540
rect 124100 668300 124190 668540
rect 124430 668300 124520 668540
rect 124760 668300 124870 668540
rect 125110 668300 125200 668540
rect 125440 668300 125530 668540
rect 125770 668300 125860 668540
rect 126100 668300 126210 668540
rect 126450 668300 126540 668540
rect 126780 668300 126870 668540
rect 127110 668300 127200 668540
rect 127440 668300 127550 668540
rect 127790 668300 127880 668540
rect 128120 668300 128210 668540
rect 128450 668300 128540 668540
rect 128780 668300 128890 668540
rect 129130 668300 129220 668540
rect 129460 668300 129550 668540
rect 129790 668300 129880 668540
rect 130120 668300 130230 668540
rect 130470 668300 130560 668540
rect 130800 668300 130890 668540
rect 131130 668300 131220 668540
rect 131460 668300 131570 668540
rect 131810 668300 131900 668540
rect 132140 668300 132230 668540
rect 132470 668300 132560 668540
rect 132800 668300 132910 668540
rect 133150 668300 133570 668540
rect 133810 668300 133900 668540
rect 134140 668300 134230 668540
rect 134470 668300 134560 668540
rect 134800 668300 134910 668540
rect 135150 668300 135240 668540
rect 135480 668300 135570 668540
rect 135810 668300 135900 668540
rect 136140 668300 136250 668540
rect 136490 668300 136580 668540
rect 136820 668300 136910 668540
rect 137150 668300 137240 668540
rect 137480 668300 137590 668540
rect 137830 668300 137920 668540
rect 138160 668300 138250 668540
rect 138490 668300 138580 668540
rect 138820 668300 138930 668540
rect 139170 668300 139260 668540
rect 139500 668300 139590 668540
rect 139830 668300 139920 668540
rect 140160 668300 140270 668540
rect 140510 668300 140600 668540
rect 140840 668300 140930 668540
rect 141170 668300 141260 668540
rect 141500 668300 141610 668540
rect 141850 668300 141940 668540
rect 142180 668300 142270 668540
rect 142510 668300 142600 668540
rect 142840 668300 142950 668540
rect 143190 668300 143280 668540
rect 143520 668300 143610 668540
rect 143850 668300 143940 668540
rect 144180 668300 144290 668540
rect 144530 668300 144950 668540
rect 145190 668300 145280 668540
rect 145520 668300 145610 668540
rect 145850 668300 145940 668540
rect 146180 668300 146290 668540
rect 146530 668300 146620 668540
rect 146860 668300 146950 668540
rect 147190 668300 147280 668540
rect 147520 668300 147630 668540
rect 147870 668300 147960 668540
rect 148200 668300 148290 668540
rect 148530 668300 148620 668540
rect 148860 668300 148970 668540
rect 149210 668300 149300 668540
rect 149540 668300 149630 668540
rect 149870 668300 149960 668540
rect 150200 668300 150310 668540
rect 150550 668300 150640 668540
rect 150880 668300 150970 668540
rect 151210 668300 151300 668540
rect 151540 668300 151650 668540
rect 151890 668300 151980 668540
rect 152220 668300 152310 668540
rect 152550 668300 152640 668540
rect 152880 668300 152990 668540
rect 153230 668300 153320 668540
rect 153560 668300 153650 668540
rect 153890 668300 153980 668540
rect 154220 668300 154330 668540
rect 154570 668300 154660 668540
rect 154900 668300 154990 668540
rect 155230 668300 155320 668540
rect 155560 668300 155670 668540
rect 155910 668300 155960 668540
rect 110760 668210 155960 668300
rect 110760 667970 110810 668210
rect 111050 667970 111140 668210
rect 111380 667970 111470 668210
rect 111710 667970 111800 668210
rect 112040 667970 112150 668210
rect 112390 667970 112480 668210
rect 112720 667970 112810 668210
rect 113050 667970 113140 668210
rect 113380 667970 113490 668210
rect 113730 667970 113820 668210
rect 114060 667970 114150 668210
rect 114390 667970 114480 668210
rect 114720 667970 114830 668210
rect 115070 667970 115160 668210
rect 115400 667970 115490 668210
rect 115730 667970 115820 668210
rect 116060 667970 116170 668210
rect 116410 667970 116500 668210
rect 116740 667970 116830 668210
rect 117070 667970 117160 668210
rect 117400 667970 117510 668210
rect 117750 667970 117840 668210
rect 118080 667970 118170 668210
rect 118410 667970 118500 668210
rect 118740 667970 118850 668210
rect 119090 667970 119180 668210
rect 119420 667970 119510 668210
rect 119750 667970 119840 668210
rect 120080 667970 120190 668210
rect 120430 667970 120520 668210
rect 120760 667970 120850 668210
rect 121090 667970 121180 668210
rect 121420 667970 121530 668210
rect 121770 667970 122190 668210
rect 122430 667970 122520 668210
rect 122760 667970 122850 668210
rect 123090 667970 123180 668210
rect 123420 667970 123530 668210
rect 123770 667970 123860 668210
rect 124100 667970 124190 668210
rect 124430 667970 124520 668210
rect 124760 667970 124870 668210
rect 125110 667970 125200 668210
rect 125440 667970 125530 668210
rect 125770 667970 125860 668210
rect 126100 667970 126210 668210
rect 126450 667970 126540 668210
rect 126780 667970 126870 668210
rect 127110 667970 127200 668210
rect 127440 667970 127550 668210
rect 127790 667970 127880 668210
rect 128120 667970 128210 668210
rect 128450 667970 128540 668210
rect 128780 667970 128890 668210
rect 129130 667970 129220 668210
rect 129460 667970 129550 668210
rect 129790 667970 129880 668210
rect 130120 667970 130230 668210
rect 130470 667970 130560 668210
rect 130800 667970 130890 668210
rect 131130 667970 131220 668210
rect 131460 667970 131570 668210
rect 131810 667970 131900 668210
rect 132140 667970 132230 668210
rect 132470 667970 132560 668210
rect 132800 667970 132910 668210
rect 133150 667970 133570 668210
rect 133810 667970 133900 668210
rect 134140 667970 134230 668210
rect 134470 667970 134560 668210
rect 134800 667970 134910 668210
rect 135150 667970 135240 668210
rect 135480 667970 135570 668210
rect 135810 667970 135900 668210
rect 136140 667970 136250 668210
rect 136490 667970 136580 668210
rect 136820 667970 136910 668210
rect 137150 667970 137240 668210
rect 137480 667970 137590 668210
rect 137830 667970 137920 668210
rect 138160 667970 138250 668210
rect 138490 667970 138580 668210
rect 138820 667970 138930 668210
rect 139170 667970 139260 668210
rect 139500 667970 139590 668210
rect 139830 667970 139920 668210
rect 140160 667970 140270 668210
rect 140510 667970 140600 668210
rect 140840 667970 140930 668210
rect 141170 667970 141260 668210
rect 141500 667970 141610 668210
rect 141850 667970 141940 668210
rect 142180 667970 142270 668210
rect 142510 667970 142600 668210
rect 142840 667970 142950 668210
rect 143190 667970 143280 668210
rect 143520 667970 143610 668210
rect 143850 667970 143940 668210
rect 144180 667970 144290 668210
rect 144530 667970 144950 668210
rect 145190 667970 145280 668210
rect 145520 667970 145610 668210
rect 145850 667970 145940 668210
rect 146180 667970 146290 668210
rect 146530 667970 146620 668210
rect 146860 667970 146950 668210
rect 147190 667970 147280 668210
rect 147520 667970 147630 668210
rect 147870 667970 147960 668210
rect 148200 667970 148290 668210
rect 148530 667970 148620 668210
rect 148860 667970 148970 668210
rect 149210 667970 149300 668210
rect 149540 667970 149630 668210
rect 149870 667970 149960 668210
rect 150200 667970 150310 668210
rect 150550 667970 150640 668210
rect 150880 667970 150970 668210
rect 151210 667970 151300 668210
rect 151540 667970 151650 668210
rect 151890 667970 151980 668210
rect 152220 667970 152310 668210
rect 152550 667970 152640 668210
rect 152880 667970 152990 668210
rect 153230 667970 153320 668210
rect 153560 667970 153650 668210
rect 153890 667970 153980 668210
rect 154220 667970 154330 668210
rect 154570 667970 154660 668210
rect 154900 667970 154990 668210
rect 155230 667970 155320 668210
rect 155560 667970 155670 668210
rect 155910 667970 155960 668210
rect 110760 667880 155960 667970
rect 110760 667640 110810 667880
rect 111050 667640 111140 667880
rect 111380 667640 111470 667880
rect 111710 667640 111800 667880
rect 112040 667640 112150 667880
rect 112390 667640 112480 667880
rect 112720 667640 112810 667880
rect 113050 667640 113140 667880
rect 113380 667640 113490 667880
rect 113730 667640 113820 667880
rect 114060 667640 114150 667880
rect 114390 667640 114480 667880
rect 114720 667640 114830 667880
rect 115070 667640 115160 667880
rect 115400 667640 115490 667880
rect 115730 667640 115820 667880
rect 116060 667640 116170 667880
rect 116410 667640 116500 667880
rect 116740 667640 116830 667880
rect 117070 667640 117160 667880
rect 117400 667640 117510 667880
rect 117750 667640 117840 667880
rect 118080 667640 118170 667880
rect 118410 667640 118500 667880
rect 118740 667640 118850 667880
rect 119090 667640 119180 667880
rect 119420 667640 119510 667880
rect 119750 667640 119840 667880
rect 120080 667640 120190 667880
rect 120430 667640 120520 667880
rect 120760 667640 120850 667880
rect 121090 667640 121180 667880
rect 121420 667640 121530 667880
rect 121770 667640 122190 667880
rect 122430 667640 122520 667880
rect 122760 667640 122850 667880
rect 123090 667640 123180 667880
rect 123420 667640 123530 667880
rect 123770 667640 123860 667880
rect 124100 667640 124190 667880
rect 124430 667640 124520 667880
rect 124760 667640 124870 667880
rect 125110 667640 125200 667880
rect 125440 667640 125530 667880
rect 125770 667640 125860 667880
rect 126100 667640 126210 667880
rect 126450 667640 126540 667880
rect 126780 667640 126870 667880
rect 127110 667640 127200 667880
rect 127440 667640 127550 667880
rect 127790 667640 127880 667880
rect 128120 667640 128210 667880
rect 128450 667640 128540 667880
rect 128780 667640 128890 667880
rect 129130 667640 129220 667880
rect 129460 667640 129550 667880
rect 129790 667640 129880 667880
rect 130120 667640 130230 667880
rect 130470 667640 130560 667880
rect 130800 667640 130890 667880
rect 131130 667640 131220 667880
rect 131460 667640 131570 667880
rect 131810 667640 131900 667880
rect 132140 667640 132230 667880
rect 132470 667640 132560 667880
rect 132800 667640 132910 667880
rect 133150 667640 133570 667880
rect 133810 667640 133900 667880
rect 134140 667640 134230 667880
rect 134470 667640 134560 667880
rect 134800 667640 134910 667880
rect 135150 667640 135240 667880
rect 135480 667640 135570 667880
rect 135810 667640 135900 667880
rect 136140 667640 136250 667880
rect 136490 667640 136580 667880
rect 136820 667640 136910 667880
rect 137150 667640 137240 667880
rect 137480 667640 137590 667880
rect 137830 667640 137920 667880
rect 138160 667640 138250 667880
rect 138490 667640 138580 667880
rect 138820 667640 138930 667880
rect 139170 667640 139260 667880
rect 139500 667640 139590 667880
rect 139830 667640 139920 667880
rect 140160 667640 140270 667880
rect 140510 667640 140600 667880
rect 140840 667640 140930 667880
rect 141170 667640 141260 667880
rect 141500 667640 141610 667880
rect 141850 667640 141940 667880
rect 142180 667640 142270 667880
rect 142510 667640 142600 667880
rect 142840 667640 142950 667880
rect 143190 667640 143280 667880
rect 143520 667640 143610 667880
rect 143850 667640 143940 667880
rect 144180 667640 144290 667880
rect 144530 667640 144950 667880
rect 145190 667640 145280 667880
rect 145520 667640 145610 667880
rect 145850 667640 145940 667880
rect 146180 667640 146290 667880
rect 146530 667640 146620 667880
rect 146860 667640 146950 667880
rect 147190 667640 147280 667880
rect 147520 667640 147630 667880
rect 147870 667640 147960 667880
rect 148200 667640 148290 667880
rect 148530 667640 148620 667880
rect 148860 667640 148970 667880
rect 149210 667640 149300 667880
rect 149540 667640 149630 667880
rect 149870 667640 149960 667880
rect 150200 667640 150310 667880
rect 150550 667640 150640 667880
rect 150880 667640 150970 667880
rect 151210 667640 151300 667880
rect 151540 667640 151650 667880
rect 151890 667640 151980 667880
rect 152220 667640 152310 667880
rect 152550 667640 152640 667880
rect 152880 667640 152990 667880
rect 153230 667640 153320 667880
rect 153560 667640 153650 667880
rect 153890 667640 153980 667880
rect 154220 667640 154330 667880
rect 154570 667640 154660 667880
rect 154900 667640 154990 667880
rect 155230 667640 155320 667880
rect 155560 667640 155670 667880
rect 155910 667640 155960 667880
rect 110760 667530 155960 667640
rect 110760 667290 110810 667530
rect 111050 667290 111140 667530
rect 111380 667290 111470 667530
rect 111710 667290 111800 667530
rect 112040 667290 112150 667530
rect 112390 667290 112480 667530
rect 112720 667290 112810 667530
rect 113050 667290 113140 667530
rect 113380 667290 113490 667530
rect 113730 667290 113820 667530
rect 114060 667290 114150 667530
rect 114390 667290 114480 667530
rect 114720 667290 114830 667530
rect 115070 667290 115160 667530
rect 115400 667290 115490 667530
rect 115730 667290 115820 667530
rect 116060 667290 116170 667530
rect 116410 667290 116500 667530
rect 116740 667290 116830 667530
rect 117070 667290 117160 667530
rect 117400 667290 117510 667530
rect 117750 667290 117840 667530
rect 118080 667290 118170 667530
rect 118410 667290 118500 667530
rect 118740 667290 118850 667530
rect 119090 667290 119180 667530
rect 119420 667290 119510 667530
rect 119750 667290 119840 667530
rect 120080 667290 120190 667530
rect 120430 667290 120520 667530
rect 120760 667290 120850 667530
rect 121090 667290 121180 667530
rect 121420 667290 121530 667530
rect 121770 667290 122190 667530
rect 122430 667290 122520 667530
rect 122760 667290 122850 667530
rect 123090 667290 123180 667530
rect 123420 667290 123530 667530
rect 123770 667290 123860 667530
rect 124100 667290 124190 667530
rect 124430 667290 124520 667530
rect 124760 667290 124870 667530
rect 125110 667290 125200 667530
rect 125440 667290 125530 667530
rect 125770 667290 125860 667530
rect 126100 667290 126210 667530
rect 126450 667290 126540 667530
rect 126780 667290 126870 667530
rect 127110 667290 127200 667530
rect 127440 667290 127550 667530
rect 127790 667290 127880 667530
rect 128120 667290 128210 667530
rect 128450 667290 128540 667530
rect 128780 667290 128890 667530
rect 129130 667290 129220 667530
rect 129460 667290 129550 667530
rect 129790 667290 129880 667530
rect 130120 667290 130230 667530
rect 130470 667290 130560 667530
rect 130800 667290 130890 667530
rect 131130 667290 131220 667530
rect 131460 667290 131570 667530
rect 131810 667290 131900 667530
rect 132140 667290 132230 667530
rect 132470 667290 132560 667530
rect 132800 667290 132910 667530
rect 133150 667290 133570 667530
rect 133810 667290 133900 667530
rect 134140 667290 134230 667530
rect 134470 667290 134560 667530
rect 134800 667290 134910 667530
rect 135150 667290 135240 667530
rect 135480 667290 135570 667530
rect 135810 667290 135900 667530
rect 136140 667290 136250 667530
rect 136490 667290 136580 667530
rect 136820 667290 136910 667530
rect 137150 667290 137240 667530
rect 137480 667290 137590 667530
rect 137830 667290 137920 667530
rect 138160 667290 138250 667530
rect 138490 667290 138580 667530
rect 138820 667290 138930 667530
rect 139170 667290 139260 667530
rect 139500 667290 139590 667530
rect 139830 667290 139920 667530
rect 140160 667290 140270 667530
rect 140510 667290 140600 667530
rect 140840 667290 140930 667530
rect 141170 667290 141260 667530
rect 141500 667290 141610 667530
rect 141850 667290 141940 667530
rect 142180 667290 142270 667530
rect 142510 667290 142600 667530
rect 142840 667290 142950 667530
rect 143190 667290 143280 667530
rect 143520 667290 143610 667530
rect 143850 667290 143940 667530
rect 144180 667290 144290 667530
rect 144530 667290 144950 667530
rect 145190 667290 145280 667530
rect 145520 667290 145610 667530
rect 145850 667290 145940 667530
rect 146180 667290 146290 667530
rect 146530 667290 146620 667530
rect 146860 667290 146950 667530
rect 147190 667290 147280 667530
rect 147520 667290 147630 667530
rect 147870 667290 147960 667530
rect 148200 667290 148290 667530
rect 148530 667290 148620 667530
rect 148860 667290 148970 667530
rect 149210 667290 149300 667530
rect 149540 667290 149630 667530
rect 149870 667290 149960 667530
rect 150200 667290 150310 667530
rect 150550 667290 150640 667530
rect 150880 667290 150970 667530
rect 151210 667290 151300 667530
rect 151540 667290 151650 667530
rect 151890 667290 151980 667530
rect 152220 667290 152310 667530
rect 152550 667290 152640 667530
rect 152880 667290 152990 667530
rect 153230 667290 153320 667530
rect 153560 667290 153650 667530
rect 153890 667290 153980 667530
rect 154220 667290 154330 667530
rect 154570 667290 154660 667530
rect 154900 667290 154990 667530
rect 155230 667290 155320 667530
rect 155560 667290 155670 667530
rect 155910 667290 155960 667530
rect 110760 667200 155960 667290
rect 110760 666960 110810 667200
rect 111050 666960 111140 667200
rect 111380 666960 111470 667200
rect 111710 666960 111800 667200
rect 112040 666960 112150 667200
rect 112390 666960 112480 667200
rect 112720 666960 112810 667200
rect 113050 666960 113140 667200
rect 113380 666960 113490 667200
rect 113730 666960 113820 667200
rect 114060 666960 114150 667200
rect 114390 666960 114480 667200
rect 114720 666960 114830 667200
rect 115070 666960 115160 667200
rect 115400 666960 115490 667200
rect 115730 666960 115820 667200
rect 116060 666960 116170 667200
rect 116410 666960 116500 667200
rect 116740 666960 116830 667200
rect 117070 666960 117160 667200
rect 117400 666960 117510 667200
rect 117750 666960 117840 667200
rect 118080 666960 118170 667200
rect 118410 666960 118500 667200
rect 118740 666960 118850 667200
rect 119090 666960 119180 667200
rect 119420 666960 119510 667200
rect 119750 666960 119840 667200
rect 120080 666960 120190 667200
rect 120430 666960 120520 667200
rect 120760 666960 120850 667200
rect 121090 666960 121180 667200
rect 121420 666960 121530 667200
rect 121770 666960 122190 667200
rect 122430 666960 122520 667200
rect 122760 666960 122850 667200
rect 123090 666960 123180 667200
rect 123420 666960 123530 667200
rect 123770 666960 123860 667200
rect 124100 666960 124190 667200
rect 124430 666960 124520 667200
rect 124760 666960 124870 667200
rect 125110 666960 125200 667200
rect 125440 666960 125530 667200
rect 125770 666960 125860 667200
rect 126100 666960 126210 667200
rect 126450 666960 126540 667200
rect 126780 666960 126870 667200
rect 127110 666960 127200 667200
rect 127440 666960 127550 667200
rect 127790 666960 127880 667200
rect 128120 666960 128210 667200
rect 128450 666960 128540 667200
rect 128780 666960 128890 667200
rect 129130 666960 129220 667200
rect 129460 666960 129550 667200
rect 129790 666960 129880 667200
rect 130120 666960 130230 667200
rect 130470 666960 130560 667200
rect 130800 666960 130890 667200
rect 131130 666960 131220 667200
rect 131460 666960 131570 667200
rect 131810 666960 131900 667200
rect 132140 666960 132230 667200
rect 132470 666960 132560 667200
rect 132800 666960 132910 667200
rect 133150 666960 133570 667200
rect 133810 666960 133900 667200
rect 134140 666960 134230 667200
rect 134470 666960 134560 667200
rect 134800 666960 134910 667200
rect 135150 666960 135240 667200
rect 135480 666960 135570 667200
rect 135810 666960 135900 667200
rect 136140 666960 136250 667200
rect 136490 666960 136580 667200
rect 136820 666960 136910 667200
rect 137150 666960 137240 667200
rect 137480 666960 137590 667200
rect 137830 666960 137920 667200
rect 138160 666960 138250 667200
rect 138490 666960 138580 667200
rect 138820 666960 138930 667200
rect 139170 666960 139260 667200
rect 139500 666960 139590 667200
rect 139830 666960 139920 667200
rect 140160 666960 140270 667200
rect 140510 666960 140600 667200
rect 140840 666960 140930 667200
rect 141170 666960 141260 667200
rect 141500 666960 141610 667200
rect 141850 666960 141940 667200
rect 142180 666960 142270 667200
rect 142510 666960 142600 667200
rect 142840 666960 142950 667200
rect 143190 666960 143280 667200
rect 143520 666960 143610 667200
rect 143850 666960 143940 667200
rect 144180 666960 144290 667200
rect 144530 666960 144950 667200
rect 145190 666960 145280 667200
rect 145520 666960 145610 667200
rect 145850 666960 145940 667200
rect 146180 666960 146290 667200
rect 146530 666960 146620 667200
rect 146860 666960 146950 667200
rect 147190 666960 147280 667200
rect 147520 666960 147630 667200
rect 147870 666960 147960 667200
rect 148200 666960 148290 667200
rect 148530 666960 148620 667200
rect 148860 666960 148970 667200
rect 149210 666960 149300 667200
rect 149540 666960 149630 667200
rect 149870 666960 149960 667200
rect 150200 666960 150310 667200
rect 150550 666960 150640 667200
rect 150880 666960 150970 667200
rect 151210 666960 151300 667200
rect 151540 666960 151650 667200
rect 151890 666960 151980 667200
rect 152220 666960 152310 667200
rect 152550 666960 152640 667200
rect 152880 666960 152990 667200
rect 153230 666960 153320 667200
rect 153560 666960 153650 667200
rect 153890 666960 153980 667200
rect 154220 666960 154330 667200
rect 154570 666960 154660 667200
rect 154900 666960 154990 667200
rect 155230 666960 155320 667200
rect 155560 666960 155670 667200
rect 155910 666960 155960 667200
rect 110760 666870 155960 666960
rect 110760 666630 110810 666870
rect 111050 666630 111140 666870
rect 111380 666630 111470 666870
rect 111710 666630 111800 666870
rect 112040 666630 112150 666870
rect 112390 666630 112480 666870
rect 112720 666630 112810 666870
rect 113050 666630 113140 666870
rect 113380 666630 113490 666870
rect 113730 666630 113820 666870
rect 114060 666630 114150 666870
rect 114390 666630 114480 666870
rect 114720 666630 114830 666870
rect 115070 666630 115160 666870
rect 115400 666630 115490 666870
rect 115730 666630 115820 666870
rect 116060 666630 116170 666870
rect 116410 666630 116500 666870
rect 116740 666630 116830 666870
rect 117070 666630 117160 666870
rect 117400 666630 117510 666870
rect 117750 666630 117840 666870
rect 118080 666630 118170 666870
rect 118410 666630 118500 666870
rect 118740 666630 118850 666870
rect 119090 666630 119180 666870
rect 119420 666630 119510 666870
rect 119750 666630 119840 666870
rect 120080 666630 120190 666870
rect 120430 666630 120520 666870
rect 120760 666630 120850 666870
rect 121090 666630 121180 666870
rect 121420 666630 121530 666870
rect 121770 666630 122190 666870
rect 122430 666630 122520 666870
rect 122760 666630 122850 666870
rect 123090 666630 123180 666870
rect 123420 666630 123530 666870
rect 123770 666630 123860 666870
rect 124100 666630 124190 666870
rect 124430 666630 124520 666870
rect 124760 666630 124870 666870
rect 125110 666630 125200 666870
rect 125440 666630 125530 666870
rect 125770 666630 125860 666870
rect 126100 666630 126210 666870
rect 126450 666630 126540 666870
rect 126780 666630 126870 666870
rect 127110 666630 127200 666870
rect 127440 666630 127550 666870
rect 127790 666630 127880 666870
rect 128120 666630 128210 666870
rect 128450 666630 128540 666870
rect 128780 666630 128890 666870
rect 129130 666630 129220 666870
rect 129460 666630 129550 666870
rect 129790 666630 129880 666870
rect 130120 666630 130230 666870
rect 130470 666630 130560 666870
rect 130800 666630 130890 666870
rect 131130 666630 131220 666870
rect 131460 666630 131570 666870
rect 131810 666630 131900 666870
rect 132140 666630 132230 666870
rect 132470 666630 132560 666870
rect 132800 666630 132910 666870
rect 133150 666630 133570 666870
rect 133810 666630 133900 666870
rect 134140 666630 134230 666870
rect 134470 666630 134560 666870
rect 134800 666630 134910 666870
rect 135150 666630 135240 666870
rect 135480 666630 135570 666870
rect 135810 666630 135900 666870
rect 136140 666630 136250 666870
rect 136490 666630 136580 666870
rect 136820 666630 136910 666870
rect 137150 666630 137240 666870
rect 137480 666630 137590 666870
rect 137830 666630 137920 666870
rect 138160 666630 138250 666870
rect 138490 666630 138580 666870
rect 138820 666630 138930 666870
rect 139170 666630 139260 666870
rect 139500 666630 139590 666870
rect 139830 666630 139920 666870
rect 140160 666630 140270 666870
rect 140510 666630 140600 666870
rect 140840 666630 140930 666870
rect 141170 666630 141260 666870
rect 141500 666630 141610 666870
rect 141850 666630 141940 666870
rect 142180 666630 142270 666870
rect 142510 666630 142600 666870
rect 142840 666630 142950 666870
rect 143190 666630 143280 666870
rect 143520 666630 143610 666870
rect 143850 666630 143940 666870
rect 144180 666630 144290 666870
rect 144530 666630 144950 666870
rect 145190 666630 145280 666870
rect 145520 666630 145610 666870
rect 145850 666630 145940 666870
rect 146180 666630 146290 666870
rect 146530 666630 146620 666870
rect 146860 666630 146950 666870
rect 147190 666630 147280 666870
rect 147520 666630 147630 666870
rect 147870 666630 147960 666870
rect 148200 666630 148290 666870
rect 148530 666630 148620 666870
rect 148860 666630 148970 666870
rect 149210 666630 149300 666870
rect 149540 666630 149630 666870
rect 149870 666630 149960 666870
rect 150200 666630 150310 666870
rect 150550 666630 150640 666870
rect 150880 666630 150970 666870
rect 151210 666630 151300 666870
rect 151540 666630 151650 666870
rect 151890 666630 151980 666870
rect 152220 666630 152310 666870
rect 152550 666630 152640 666870
rect 152880 666630 152990 666870
rect 153230 666630 153320 666870
rect 153560 666630 153650 666870
rect 153890 666630 153980 666870
rect 154220 666630 154330 666870
rect 154570 666630 154660 666870
rect 154900 666630 154990 666870
rect 155230 666630 155320 666870
rect 155560 666630 155670 666870
rect 155910 666630 155960 666870
rect 110760 666540 155960 666630
rect 110760 666300 110810 666540
rect 111050 666300 111140 666540
rect 111380 666300 111470 666540
rect 111710 666300 111800 666540
rect 112040 666300 112150 666540
rect 112390 666300 112480 666540
rect 112720 666300 112810 666540
rect 113050 666300 113140 666540
rect 113380 666300 113490 666540
rect 113730 666300 113820 666540
rect 114060 666300 114150 666540
rect 114390 666300 114480 666540
rect 114720 666300 114830 666540
rect 115070 666300 115160 666540
rect 115400 666300 115490 666540
rect 115730 666300 115820 666540
rect 116060 666300 116170 666540
rect 116410 666300 116500 666540
rect 116740 666300 116830 666540
rect 117070 666300 117160 666540
rect 117400 666300 117510 666540
rect 117750 666300 117840 666540
rect 118080 666300 118170 666540
rect 118410 666300 118500 666540
rect 118740 666300 118850 666540
rect 119090 666300 119180 666540
rect 119420 666300 119510 666540
rect 119750 666300 119840 666540
rect 120080 666300 120190 666540
rect 120430 666300 120520 666540
rect 120760 666300 120850 666540
rect 121090 666300 121180 666540
rect 121420 666300 121530 666540
rect 121770 666300 122190 666540
rect 122430 666300 122520 666540
rect 122760 666300 122850 666540
rect 123090 666300 123180 666540
rect 123420 666300 123530 666540
rect 123770 666300 123860 666540
rect 124100 666300 124190 666540
rect 124430 666300 124520 666540
rect 124760 666300 124870 666540
rect 125110 666300 125200 666540
rect 125440 666300 125530 666540
rect 125770 666300 125860 666540
rect 126100 666300 126210 666540
rect 126450 666300 126540 666540
rect 126780 666300 126870 666540
rect 127110 666300 127200 666540
rect 127440 666300 127550 666540
rect 127790 666300 127880 666540
rect 128120 666300 128210 666540
rect 128450 666300 128540 666540
rect 128780 666300 128890 666540
rect 129130 666300 129220 666540
rect 129460 666300 129550 666540
rect 129790 666300 129880 666540
rect 130120 666300 130230 666540
rect 130470 666300 130560 666540
rect 130800 666300 130890 666540
rect 131130 666300 131220 666540
rect 131460 666300 131570 666540
rect 131810 666300 131900 666540
rect 132140 666300 132230 666540
rect 132470 666300 132560 666540
rect 132800 666300 132910 666540
rect 133150 666300 133570 666540
rect 133810 666300 133900 666540
rect 134140 666300 134230 666540
rect 134470 666300 134560 666540
rect 134800 666300 134910 666540
rect 135150 666300 135240 666540
rect 135480 666300 135570 666540
rect 135810 666300 135900 666540
rect 136140 666300 136250 666540
rect 136490 666300 136580 666540
rect 136820 666300 136910 666540
rect 137150 666300 137240 666540
rect 137480 666300 137590 666540
rect 137830 666300 137920 666540
rect 138160 666300 138250 666540
rect 138490 666300 138580 666540
rect 138820 666300 138930 666540
rect 139170 666300 139260 666540
rect 139500 666300 139590 666540
rect 139830 666300 139920 666540
rect 140160 666300 140270 666540
rect 140510 666300 140600 666540
rect 140840 666300 140930 666540
rect 141170 666300 141260 666540
rect 141500 666300 141610 666540
rect 141850 666300 141940 666540
rect 142180 666300 142270 666540
rect 142510 666300 142600 666540
rect 142840 666300 142950 666540
rect 143190 666300 143280 666540
rect 143520 666300 143610 666540
rect 143850 666300 143940 666540
rect 144180 666300 144290 666540
rect 144530 666300 144950 666540
rect 145190 666300 145280 666540
rect 145520 666300 145610 666540
rect 145850 666300 145940 666540
rect 146180 666300 146290 666540
rect 146530 666300 146620 666540
rect 146860 666300 146950 666540
rect 147190 666300 147280 666540
rect 147520 666300 147630 666540
rect 147870 666300 147960 666540
rect 148200 666300 148290 666540
rect 148530 666300 148620 666540
rect 148860 666300 148970 666540
rect 149210 666300 149300 666540
rect 149540 666300 149630 666540
rect 149870 666300 149960 666540
rect 150200 666300 150310 666540
rect 150550 666300 150640 666540
rect 150880 666300 150970 666540
rect 151210 666300 151300 666540
rect 151540 666300 151650 666540
rect 151890 666300 151980 666540
rect 152220 666300 152310 666540
rect 152550 666300 152640 666540
rect 152880 666300 152990 666540
rect 153230 666300 153320 666540
rect 153560 666300 153650 666540
rect 153890 666300 153980 666540
rect 154220 666300 154330 666540
rect 154570 666300 154660 666540
rect 154900 666300 154990 666540
rect 155230 666300 155320 666540
rect 155560 666300 155670 666540
rect 155910 666300 155960 666540
rect 110760 666190 155960 666300
rect 110760 665950 110810 666190
rect 111050 665950 111140 666190
rect 111380 665950 111470 666190
rect 111710 665950 111800 666190
rect 112040 665950 112150 666190
rect 112390 665950 112480 666190
rect 112720 665950 112810 666190
rect 113050 665950 113140 666190
rect 113380 665950 113490 666190
rect 113730 665950 113820 666190
rect 114060 665950 114150 666190
rect 114390 665950 114480 666190
rect 114720 665950 114830 666190
rect 115070 665950 115160 666190
rect 115400 665950 115490 666190
rect 115730 665950 115820 666190
rect 116060 665950 116170 666190
rect 116410 665950 116500 666190
rect 116740 665950 116830 666190
rect 117070 665950 117160 666190
rect 117400 665950 117510 666190
rect 117750 665950 117840 666190
rect 118080 665950 118170 666190
rect 118410 665950 118500 666190
rect 118740 665950 118850 666190
rect 119090 665950 119180 666190
rect 119420 665950 119510 666190
rect 119750 665950 119840 666190
rect 120080 665950 120190 666190
rect 120430 665950 120520 666190
rect 120760 665950 120850 666190
rect 121090 665950 121180 666190
rect 121420 665950 121530 666190
rect 121770 665950 122190 666190
rect 122430 665950 122520 666190
rect 122760 665950 122850 666190
rect 123090 665950 123180 666190
rect 123420 665950 123530 666190
rect 123770 665950 123860 666190
rect 124100 665950 124190 666190
rect 124430 665950 124520 666190
rect 124760 665950 124870 666190
rect 125110 665950 125200 666190
rect 125440 665950 125530 666190
rect 125770 665950 125860 666190
rect 126100 665950 126210 666190
rect 126450 665950 126540 666190
rect 126780 665950 126870 666190
rect 127110 665950 127200 666190
rect 127440 665950 127550 666190
rect 127790 665950 127880 666190
rect 128120 665950 128210 666190
rect 128450 665950 128540 666190
rect 128780 665950 128890 666190
rect 129130 665950 129220 666190
rect 129460 665950 129550 666190
rect 129790 665950 129880 666190
rect 130120 665950 130230 666190
rect 130470 665950 130560 666190
rect 130800 665950 130890 666190
rect 131130 665950 131220 666190
rect 131460 665950 131570 666190
rect 131810 665950 131900 666190
rect 132140 665950 132230 666190
rect 132470 665950 132560 666190
rect 132800 665950 132910 666190
rect 133150 665950 133570 666190
rect 133810 665950 133900 666190
rect 134140 665950 134230 666190
rect 134470 665950 134560 666190
rect 134800 665950 134910 666190
rect 135150 665950 135240 666190
rect 135480 665950 135570 666190
rect 135810 665950 135900 666190
rect 136140 665950 136250 666190
rect 136490 665950 136580 666190
rect 136820 665950 136910 666190
rect 137150 665950 137240 666190
rect 137480 665950 137590 666190
rect 137830 665950 137920 666190
rect 138160 665950 138250 666190
rect 138490 665950 138580 666190
rect 138820 665950 138930 666190
rect 139170 665950 139260 666190
rect 139500 665950 139590 666190
rect 139830 665950 139920 666190
rect 140160 665950 140270 666190
rect 140510 665950 140600 666190
rect 140840 665950 140930 666190
rect 141170 665950 141260 666190
rect 141500 665950 141610 666190
rect 141850 665950 141940 666190
rect 142180 665950 142270 666190
rect 142510 665950 142600 666190
rect 142840 665950 142950 666190
rect 143190 665950 143280 666190
rect 143520 665950 143610 666190
rect 143850 665950 143940 666190
rect 144180 665950 144290 666190
rect 144530 665950 144950 666190
rect 145190 665950 145280 666190
rect 145520 665950 145610 666190
rect 145850 665950 145940 666190
rect 146180 665950 146290 666190
rect 146530 665950 146620 666190
rect 146860 665950 146950 666190
rect 147190 665950 147280 666190
rect 147520 665950 147630 666190
rect 147870 665950 147960 666190
rect 148200 665950 148290 666190
rect 148530 665950 148620 666190
rect 148860 665950 148970 666190
rect 149210 665950 149300 666190
rect 149540 665950 149630 666190
rect 149870 665950 149960 666190
rect 150200 665950 150310 666190
rect 150550 665950 150640 666190
rect 150880 665950 150970 666190
rect 151210 665950 151300 666190
rect 151540 665950 151650 666190
rect 151890 665950 151980 666190
rect 152220 665950 152310 666190
rect 152550 665950 152640 666190
rect 152880 665950 152990 666190
rect 153230 665950 153320 666190
rect 153560 665950 153650 666190
rect 153890 665950 153980 666190
rect 154220 665950 154330 666190
rect 154570 665950 154660 666190
rect 154900 665950 154990 666190
rect 155230 665950 155320 666190
rect 155560 665950 155670 666190
rect 155910 665950 155960 666190
rect 110760 665860 155960 665950
rect 110760 665620 110810 665860
rect 111050 665620 111140 665860
rect 111380 665620 111470 665860
rect 111710 665620 111800 665860
rect 112040 665620 112150 665860
rect 112390 665620 112480 665860
rect 112720 665620 112810 665860
rect 113050 665620 113140 665860
rect 113380 665620 113490 665860
rect 113730 665620 113820 665860
rect 114060 665620 114150 665860
rect 114390 665620 114480 665860
rect 114720 665620 114830 665860
rect 115070 665620 115160 665860
rect 115400 665620 115490 665860
rect 115730 665620 115820 665860
rect 116060 665620 116170 665860
rect 116410 665620 116500 665860
rect 116740 665620 116830 665860
rect 117070 665620 117160 665860
rect 117400 665620 117510 665860
rect 117750 665620 117840 665860
rect 118080 665620 118170 665860
rect 118410 665620 118500 665860
rect 118740 665620 118850 665860
rect 119090 665620 119180 665860
rect 119420 665620 119510 665860
rect 119750 665620 119840 665860
rect 120080 665620 120190 665860
rect 120430 665620 120520 665860
rect 120760 665620 120850 665860
rect 121090 665620 121180 665860
rect 121420 665620 121530 665860
rect 121770 665620 122190 665860
rect 122430 665620 122520 665860
rect 122760 665620 122850 665860
rect 123090 665620 123180 665860
rect 123420 665620 123530 665860
rect 123770 665620 123860 665860
rect 124100 665620 124190 665860
rect 124430 665620 124520 665860
rect 124760 665620 124870 665860
rect 125110 665620 125200 665860
rect 125440 665620 125530 665860
rect 125770 665620 125860 665860
rect 126100 665620 126210 665860
rect 126450 665620 126540 665860
rect 126780 665620 126870 665860
rect 127110 665620 127200 665860
rect 127440 665620 127550 665860
rect 127790 665620 127880 665860
rect 128120 665620 128210 665860
rect 128450 665620 128540 665860
rect 128780 665620 128890 665860
rect 129130 665620 129220 665860
rect 129460 665620 129550 665860
rect 129790 665620 129880 665860
rect 130120 665620 130230 665860
rect 130470 665620 130560 665860
rect 130800 665620 130890 665860
rect 131130 665620 131220 665860
rect 131460 665620 131570 665860
rect 131810 665620 131900 665860
rect 132140 665620 132230 665860
rect 132470 665620 132560 665860
rect 132800 665620 132910 665860
rect 133150 665620 133570 665860
rect 133810 665620 133900 665860
rect 134140 665620 134230 665860
rect 134470 665620 134560 665860
rect 134800 665620 134910 665860
rect 135150 665620 135240 665860
rect 135480 665620 135570 665860
rect 135810 665620 135900 665860
rect 136140 665620 136250 665860
rect 136490 665620 136580 665860
rect 136820 665620 136910 665860
rect 137150 665620 137240 665860
rect 137480 665620 137590 665860
rect 137830 665620 137920 665860
rect 138160 665620 138250 665860
rect 138490 665620 138580 665860
rect 138820 665620 138930 665860
rect 139170 665620 139260 665860
rect 139500 665620 139590 665860
rect 139830 665620 139920 665860
rect 140160 665620 140270 665860
rect 140510 665620 140600 665860
rect 140840 665620 140930 665860
rect 141170 665620 141260 665860
rect 141500 665620 141610 665860
rect 141850 665620 141940 665860
rect 142180 665620 142270 665860
rect 142510 665620 142600 665860
rect 142840 665620 142950 665860
rect 143190 665620 143280 665860
rect 143520 665620 143610 665860
rect 143850 665620 143940 665860
rect 144180 665620 144290 665860
rect 144530 665620 144950 665860
rect 145190 665620 145280 665860
rect 145520 665620 145610 665860
rect 145850 665620 145940 665860
rect 146180 665620 146290 665860
rect 146530 665620 146620 665860
rect 146860 665620 146950 665860
rect 147190 665620 147280 665860
rect 147520 665620 147630 665860
rect 147870 665620 147960 665860
rect 148200 665620 148290 665860
rect 148530 665620 148620 665860
rect 148860 665620 148970 665860
rect 149210 665620 149300 665860
rect 149540 665620 149630 665860
rect 149870 665620 149960 665860
rect 150200 665620 150310 665860
rect 150550 665620 150640 665860
rect 150880 665620 150970 665860
rect 151210 665620 151300 665860
rect 151540 665620 151650 665860
rect 151890 665620 151980 665860
rect 152220 665620 152310 665860
rect 152550 665620 152640 665860
rect 152880 665620 152990 665860
rect 153230 665620 153320 665860
rect 153560 665620 153650 665860
rect 153890 665620 153980 665860
rect 154220 665620 154330 665860
rect 154570 665620 154660 665860
rect 154900 665620 154990 665860
rect 155230 665620 155320 665860
rect 155560 665620 155670 665860
rect 155910 665620 155960 665860
rect 110760 665530 155960 665620
rect 110760 665500 110810 665530
rect 2500 665290 110810 665500
rect 111050 665290 111140 665530
rect 111380 665290 111470 665530
rect 111710 665290 111800 665530
rect 112040 665290 112150 665530
rect 112390 665290 112480 665530
rect 112720 665290 112810 665530
rect 113050 665290 113140 665530
rect 113380 665290 113490 665530
rect 113730 665290 113820 665530
rect 114060 665290 114150 665530
rect 114390 665290 114480 665530
rect 114720 665290 114830 665530
rect 115070 665290 115160 665530
rect 115400 665290 115490 665530
rect 115730 665290 115820 665530
rect 116060 665290 116170 665530
rect 116410 665290 116500 665530
rect 116740 665290 116830 665530
rect 117070 665290 117160 665530
rect 117400 665290 117510 665530
rect 117750 665290 117840 665530
rect 118080 665290 118170 665530
rect 118410 665290 118500 665530
rect 118740 665290 118850 665530
rect 119090 665290 119180 665530
rect 119420 665290 119510 665530
rect 119750 665290 119840 665530
rect 120080 665290 120190 665530
rect 120430 665290 120520 665530
rect 120760 665290 120850 665530
rect 121090 665290 121180 665530
rect 121420 665290 121530 665530
rect 121770 665290 122190 665530
rect 122430 665290 122520 665530
rect 122760 665290 122850 665530
rect 123090 665290 123180 665530
rect 123420 665290 123530 665530
rect 123770 665290 123860 665530
rect 124100 665290 124190 665530
rect 124430 665290 124520 665530
rect 124760 665290 124870 665530
rect 125110 665290 125200 665530
rect 125440 665290 125530 665530
rect 125770 665290 125860 665530
rect 126100 665290 126210 665530
rect 126450 665290 126540 665530
rect 126780 665290 126870 665530
rect 127110 665290 127200 665530
rect 127440 665290 127550 665530
rect 127790 665290 127880 665530
rect 128120 665290 128210 665530
rect 128450 665290 128540 665530
rect 128780 665290 128890 665530
rect 129130 665290 129220 665530
rect 129460 665290 129550 665530
rect 129790 665290 129880 665530
rect 130120 665290 130230 665530
rect 130470 665290 130560 665530
rect 130800 665290 130890 665530
rect 131130 665290 131220 665530
rect 131460 665290 131570 665530
rect 131810 665290 131900 665530
rect 132140 665290 132230 665530
rect 132470 665290 132560 665530
rect 132800 665290 132910 665530
rect 133150 665290 133570 665530
rect 133810 665290 133900 665530
rect 134140 665290 134230 665530
rect 134470 665290 134560 665530
rect 134800 665290 134910 665530
rect 135150 665290 135240 665530
rect 135480 665290 135570 665530
rect 135810 665290 135900 665530
rect 136140 665290 136250 665530
rect 136490 665290 136580 665530
rect 136820 665290 136910 665530
rect 137150 665290 137240 665530
rect 137480 665290 137590 665530
rect 137830 665290 137920 665530
rect 138160 665290 138250 665530
rect 138490 665290 138580 665530
rect 138820 665290 138930 665530
rect 139170 665290 139260 665530
rect 139500 665290 139590 665530
rect 139830 665290 139920 665530
rect 140160 665290 140270 665530
rect 140510 665290 140600 665530
rect 140840 665290 140930 665530
rect 141170 665290 141260 665530
rect 141500 665290 141610 665530
rect 141850 665290 141940 665530
rect 142180 665290 142270 665530
rect 142510 665290 142600 665530
rect 142840 665290 142950 665530
rect 143190 665290 143280 665530
rect 143520 665290 143610 665530
rect 143850 665290 143940 665530
rect 144180 665290 144290 665530
rect 144530 665290 144950 665530
rect 145190 665290 145280 665530
rect 145520 665290 145610 665530
rect 145850 665290 145940 665530
rect 146180 665290 146290 665530
rect 146530 665290 146620 665530
rect 146860 665290 146950 665530
rect 147190 665290 147280 665530
rect 147520 665290 147630 665530
rect 147870 665290 147960 665530
rect 148200 665290 148290 665530
rect 148530 665290 148620 665530
rect 148860 665290 148970 665530
rect 149210 665290 149300 665530
rect 149540 665290 149630 665530
rect 149870 665290 149960 665530
rect 150200 665290 150310 665530
rect 150550 665290 150640 665530
rect 150880 665290 150970 665530
rect 151210 665290 151300 665530
rect 151540 665290 151650 665530
rect 151890 665290 151980 665530
rect 152220 665290 152310 665530
rect 152550 665290 152640 665530
rect 152880 665290 152990 665530
rect 153230 665290 153320 665530
rect 153560 665290 153650 665530
rect 153890 665290 153980 665530
rect 154220 665290 154330 665530
rect 154570 665290 154660 665530
rect 154900 665290 154990 665530
rect 155230 665290 155320 665530
rect 155560 665290 155670 665530
rect 155910 665500 155960 665530
rect 155910 665290 164457 665500
rect 2500 665200 164457 665290
rect 2500 664960 110810 665200
rect 111050 664960 111140 665200
rect 111380 664960 111470 665200
rect 111710 664960 111800 665200
rect 112040 664960 112150 665200
rect 112390 664960 112480 665200
rect 112720 664960 112810 665200
rect 113050 664960 113140 665200
rect 113380 664960 113490 665200
rect 113730 664960 113820 665200
rect 114060 664960 114150 665200
rect 114390 664960 114480 665200
rect 114720 664960 114830 665200
rect 115070 664960 115160 665200
rect 115400 664960 115490 665200
rect 115730 664960 115820 665200
rect 116060 664960 116170 665200
rect 116410 664960 116500 665200
rect 116740 664960 116830 665200
rect 117070 664960 117160 665200
rect 117400 664960 117510 665200
rect 117750 664960 117840 665200
rect 118080 664960 118170 665200
rect 118410 664960 118500 665200
rect 118740 664960 118850 665200
rect 119090 664960 119180 665200
rect 119420 664960 119510 665200
rect 119750 664960 119840 665200
rect 120080 664960 120190 665200
rect 120430 664960 120520 665200
rect 120760 664960 120850 665200
rect 121090 664960 121180 665200
rect 121420 664960 121530 665200
rect 121770 664960 122190 665200
rect 122430 664960 122520 665200
rect 122760 664960 122850 665200
rect 123090 664960 123180 665200
rect 123420 664960 123530 665200
rect 123770 664960 123860 665200
rect 124100 664960 124190 665200
rect 124430 664960 124520 665200
rect 124760 664960 124870 665200
rect 125110 664960 125200 665200
rect 125440 664960 125530 665200
rect 125770 664960 125860 665200
rect 126100 664960 126210 665200
rect 126450 664960 126540 665200
rect 126780 664960 126870 665200
rect 127110 664960 127200 665200
rect 127440 664960 127550 665200
rect 127790 664960 127880 665200
rect 128120 664960 128210 665200
rect 128450 664960 128540 665200
rect 128780 664960 128890 665200
rect 129130 664960 129220 665200
rect 129460 664960 129550 665200
rect 129790 664960 129880 665200
rect 130120 664960 130230 665200
rect 130470 664960 130560 665200
rect 130800 664960 130890 665200
rect 131130 664960 131220 665200
rect 131460 664960 131570 665200
rect 131810 664960 131900 665200
rect 132140 664960 132230 665200
rect 132470 664960 132560 665200
rect 132800 664960 132910 665200
rect 133150 664960 133570 665200
rect 133810 664960 133900 665200
rect 134140 664960 134230 665200
rect 134470 664960 134560 665200
rect 134800 664960 134910 665200
rect 135150 664960 135240 665200
rect 135480 664960 135570 665200
rect 135810 664960 135900 665200
rect 136140 664960 136250 665200
rect 136490 664960 136580 665200
rect 136820 664960 136910 665200
rect 137150 664960 137240 665200
rect 137480 664960 137590 665200
rect 137830 664960 137920 665200
rect 138160 664960 138250 665200
rect 138490 664960 138580 665200
rect 138820 664960 138930 665200
rect 139170 664960 139260 665200
rect 139500 664960 139590 665200
rect 139830 664960 139920 665200
rect 140160 664960 140270 665200
rect 140510 664960 140600 665200
rect 140840 664960 140930 665200
rect 141170 664960 141260 665200
rect 141500 664960 141610 665200
rect 141850 664960 141940 665200
rect 142180 664960 142270 665200
rect 142510 664960 142600 665200
rect 142840 664960 142950 665200
rect 143190 664960 143280 665200
rect 143520 664960 143610 665200
rect 143850 664960 143940 665200
rect 144180 664960 144290 665200
rect 144530 664960 144950 665200
rect 145190 664960 145280 665200
rect 145520 664960 145610 665200
rect 145850 664960 145940 665200
rect 146180 664960 146290 665200
rect 146530 664960 146620 665200
rect 146860 664960 146950 665200
rect 147190 664960 147280 665200
rect 147520 664960 147630 665200
rect 147870 664960 147960 665200
rect 148200 664960 148290 665200
rect 148530 664960 148620 665200
rect 148860 664960 148970 665200
rect 149210 664960 149300 665200
rect 149540 664960 149630 665200
rect 149870 664960 149960 665200
rect 150200 664960 150310 665200
rect 150550 664960 150640 665200
rect 150880 664960 150970 665200
rect 151210 664960 151300 665200
rect 151540 664960 151650 665200
rect 151890 664960 151980 665200
rect 152220 664960 152310 665200
rect 152550 664960 152640 665200
rect 152880 664960 152990 665200
rect 153230 664960 153320 665200
rect 153560 664960 153650 665200
rect 153890 664960 153980 665200
rect 154220 664960 154330 665200
rect 154570 664960 154660 665200
rect 154900 664960 154990 665200
rect 155230 664960 155320 665200
rect 155560 664960 155670 665200
rect 155910 664960 164457 665200
rect 2500 664850 164457 664960
rect 2500 664610 110810 664850
rect 111050 664610 111140 664850
rect 111380 664610 111470 664850
rect 111710 664610 111800 664850
rect 112040 664610 112150 664850
rect 112390 664610 112480 664850
rect 112720 664610 112810 664850
rect 113050 664610 113140 664850
rect 113380 664610 113490 664850
rect 113730 664610 113820 664850
rect 114060 664610 114150 664850
rect 114390 664610 114480 664850
rect 114720 664610 114830 664850
rect 115070 664610 115160 664850
rect 115400 664610 115490 664850
rect 115730 664610 115820 664850
rect 116060 664610 116170 664850
rect 116410 664610 116500 664850
rect 116740 664610 116830 664850
rect 117070 664610 117160 664850
rect 117400 664610 117510 664850
rect 117750 664610 117840 664850
rect 118080 664610 118170 664850
rect 118410 664610 118500 664850
rect 118740 664610 118850 664850
rect 119090 664610 119180 664850
rect 119420 664610 119510 664850
rect 119750 664610 119840 664850
rect 120080 664610 120190 664850
rect 120430 664610 120520 664850
rect 120760 664610 120850 664850
rect 121090 664610 121180 664850
rect 121420 664610 121530 664850
rect 121770 664610 122190 664850
rect 122430 664610 122520 664850
rect 122760 664610 122850 664850
rect 123090 664610 123180 664850
rect 123420 664610 123530 664850
rect 123770 664610 123860 664850
rect 124100 664610 124190 664850
rect 124430 664610 124520 664850
rect 124760 664610 124870 664850
rect 125110 664610 125200 664850
rect 125440 664610 125530 664850
rect 125770 664610 125860 664850
rect 126100 664610 126210 664850
rect 126450 664610 126540 664850
rect 126780 664610 126870 664850
rect 127110 664610 127200 664850
rect 127440 664610 127550 664850
rect 127790 664610 127880 664850
rect 128120 664610 128210 664850
rect 128450 664610 128540 664850
rect 128780 664610 128890 664850
rect 129130 664610 129220 664850
rect 129460 664610 129550 664850
rect 129790 664610 129880 664850
rect 130120 664610 130230 664850
rect 130470 664610 130560 664850
rect 130800 664610 130890 664850
rect 131130 664610 131220 664850
rect 131460 664610 131570 664850
rect 131810 664610 131900 664850
rect 132140 664610 132230 664850
rect 132470 664610 132560 664850
rect 132800 664610 132910 664850
rect 133150 664610 133570 664850
rect 133810 664610 133900 664850
rect 134140 664610 134230 664850
rect 134470 664610 134560 664850
rect 134800 664610 134910 664850
rect 135150 664610 135240 664850
rect 135480 664610 135570 664850
rect 135810 664610 135900 664850
rect 136140 664610 136250 664850
rect 136490 664610 136580 664850
rect 136820 664610 136910 664850
rect 137150 664610 137240 664850
rect 137480 664610 137590 664850
rect 137830 664610 137920 664850
rect 138160 664610 138250 664850
rect 138490 664610 138580 664850
rect 138820 664610 138930 664850
rect 139170 664610 139260 664850
rect 139500 664610 139590 664850
rect 139830 664610 139920 664850
rect 140160 664610 140270 664850
rect 140510 664610 140600 664850
rect 140840 664610 140930 664850
rect 141170 664610 141260 664850
rect 141500 664610 141610 664850
rect 141850 664610 141940 664850
rect 142180 664610 142270 664850
rect 142510 664610 142600 664850
rect 142840 664610 142950 664850
rect 143190 664610 143280 664850
rect 143520 664610 143610 664850
rect 143850 664610 143940 664850
rect 144180 664610 144290 664850
rect 144530 664610 144950 664850
rect 145190 664610 145280 664850
rect 145520 664610 145610 664850
rect 145850 664610 145940 664850
rect 146180 664610 146290 664850
rect 146530 664610 146620 664850
rect 146860 664610 146950 664850
rect 147190 664610 147280 664850
rect 147520 664610 147630 664850
rect 147870 664610 147960 664850
rect 148200 664610 148290 664850
rect 148530 664610 148620 664850
rect 148860 664610 148970 664850
rect 149210 664610 149300 664850
rect 149540 664610 149630 664850
rect 149870 664610 149960 664850
rect 150200 664610 150310 664850
rect 150550 664610 150640 664850
rect 150880 664610 150970 664850
rect 151210 664610 151300 664850
rect 151540 664610 151650 664850
rect 151890 664610 151980 664850
rect 152220 664610 152310 664850
rect 152550 664610 152640 664850
rect 152880 664610 152990 664850
rect 153230 664610 153320 664850
rect 153560 664610 153650 664850
rect 153890 664610 153980 664850
rect 154220 664610 154330 664850
rect 154570 664610 154660 664850
rect 154900 664610 154990 664850
rect 155230 664610 155320 664850
rect 155560 664610 155670 664850
rect 155910 664610 164457 664850
rect 2500 664520 164457 664610
rect 2500 664280 110810 664520
rect 111050 664280 111140 664520
rect 111380 664280 111470 664520
rect 111710 664280 111800 664520
rect 112040 664280 112150 664520
rect 112390 664280 112480 664520
rect 112720 664280 112810 664520
rect 113050 664280 113140 664520
rect 113380 664280 113490 664520
rect 113730 664280 113820 664520
rect 114060 664280 114150 664520
rect 114390 664280 114480 664520
rect 114720 664280 114830 664520
rect 115070 664280 115160 664520
rect 115400 664280 115490 664520
rect 115730 664280 115820 664520
rect 116060 664280 116170 664520
rect 116410 664280 116500 664520
rect 116740 664280 116830 664520
rect 117070 664280 117160 664520
rect 117400 664280 117510 664520
rect 117750 664280 117840 664520
rect 118080 664280 118170 664520
rect 118410 664280 118500 664520
rect 118740 664280 118850 664520
rect 119090 664280 119180 664520
rect 119420 664280 119510 664520
rect 119750 664280 119840 664520
rect 120080 664280 120190 664520
rect 120430 664280 120520 664520
rect 120760 664280 120850 664520
rect 121090 664280 121180 664520
rect 121420 664280 121530 664520
rect 121770 664280 122190 664520
rect 122430 664280 122520 664520
rect 122760 664280 122850 664520
rect 123090 664280 123180 664520
rect 123420 664280 123530 664520
rect 123770 664280 123860 664520
rect 124100 664280 124190 664520
rect 124430 664280 124520 664520
rect 124760 664280 124870 664520
rect 125110 664280 125200 664520
rect 125440 664280 125530 664520
rect 125770 664280 125860 664520
rect 126100 664280 126210 664520
rect 126450 664280 126540 664520
rect 126780 664280 126870 664520
rect 127110 664280 127200 664520
rect 127440 664280 127550 664520
rect 127790 664280 127880 664520
rect 128120 664280 128210 664520
rect 128450 664280 128540 664520
rect 128780 664280 128890 664520
rect 129130 664280 129220 664520
rect 129460 664280 129550 664520
rect 129790 664280 129880 664520
rect 130120 664280 130230 664520
rect 130470 664280 130560 664520
rect 130800 664280 130890 664520
rect 131130 664280 131220 664520
rect 131460 664280 131570 664520
rect 131810 664280 131900 664520
rect 132140 664280 132230 664520
rect 132470 664280 132560 664520
rect 132800 664280 132910 664520
rect 133150 664280 133570 664520
rect 133810 664280 133900 664520
rect 134140 664280 134230 664520
rect 134470 664280 134560 664520
rect 134800 664280 134910 664520
rect 135150 664280 135240 664520
rect 135480 664280 135570 664520
rect 135810 664280 135900 664520
rect 136140 664280 136250 664520
rect 136490 664280 136580 664520
rect 136820 664280 136910 664520
rect 137150 664280 137240 664520
rect 137480 664280 137590 664520
rect 137830 664280 137920 664520
rect 138160 664280 138250 664520
rect 138490 664280 138580 664520
rect 138820 664280 138930 664520
rect 139170 664280 139260 664520
rect 139500 664280 139590 664520
rect 139830 664280 139920 664520
rect 140160 664280 140270 664520
rect 140510 664280 140600 664520
rect 140840 664280 140930 664520
rect 141170 664280 141260 664520
rect 141500 664280 141610 664520
rect 141850 664280 141940 664520
rect 142180 664280 142270 664520
rect 142510 664280 142600 664520
rect 142840 664280 142950 664520
rect 143190 664280 143280 664520
rect 143520 664280 143610 664520
rect 143850 664280 143940 664520
rect 144180 664280 144290 664520
rect 144530 664280 144950 664520
rect 145190 664280 145280 664520
rect 145520 664280 145610 664520
rect 145850 664280 145940 664520
rect 146180 664280 146290 664520
rect 146530 664280 146620 664520
rect 146860 664280 146950 664520
rect 147190 664280 147280 664520
rect 147520 664280 147630 664520
rect 147870 664280 147960 664520
rect 148200 664280 148290 664520
rect 148530 664280 148620 664520
rect 148860 664280 148970 664520
rect 149210 664280 149300 664520
rect 149540 664280 149630 664520
rect 149870 664280 149960 664520
rect 150200 664280 150310 664520
rect 150550 664280 150640 664520
rect 150880 664280 150970 664520
rect 151210 664280 151300 664520
rect 151540 664280 151650 664520
rect 151890 664280 151980 664520
rect 152220 664280 152310 664520
rect 152550 664280 152640 664520
rect 152880 664280 152990 664520
rect 153230 664280 153320 664520
rect 153560 664280 153650 664520
rect 153890 664280 153980 664520
rect 154220 664280 154330 664520
rect 154570 664280 154660 664520
rect 154900 664280 154990 664520
rect 155230 664280 155320 664520
rect 155560 664280 155670 664520
rect 155910 664280 164457 664520
rect 2500 664190 164457 664280
rect 2500 663950 110810 664190
rect 111050 663950 111140 664190
rect 111380 663950 111470 664190
rect 111710 663950 111800 664190
rect 112040 663950 112150 664190
rect 112390 663950 112480 664190
rect 112720 663950 112810 664190
rect 113050 663950 113140 664190
rect 113380 663950 113490 664190
rect 113730 663950 113820 664190
rect 114060 663950 114150 664190
rect 114390 663950 114480 664190
rect 114720 663950 114830 664190
rect 115070 663950 115160 664190
rect 115400 663950 115490 664190
rect 115730 663950 115820 664190
rect 116060 663950 116170 664190
rect 116410 663950 116500 664190
rect 116740 663950 116830 664190
rect 117070 663950 117160 664190
rect 117400 663950 117510 664190
rect 117750 663950 117840 664190
rect 118080 663950 118170 664190
rect 118410 663950 118500 664190
rect 118740 663950 118850 664190
rect 119090 663950 119180 664190
rect 119420 663950 119510 664190
rect 119750 663950 119840 664190
rect 120080 663950 120190 664190
rect 120430 663950 120520 664190
rect 120760 663950 120850 664190
rect 121090 663950 121180 664190
rect 121420 663950 121530 664190
rect 121770 663950 122190 664190
rect 122430 663950 122520 664190
rect 122760 663950 122850 664190
rect 123090 663950 123180 664190
rect 123420 663950 123530 664190
rect 123770 663950 123860 664190
rect 124100 663950 124190 664190
rect 124430 663950 124520 664190
rect 124760 663950 124870 664190
rect 125110 663950 125200 664190
rect 125440 663950 125530 664190
rect 125770 663950 125860 664190
rect 126100 663950 126210 664190
rect 126450 663950 126540 664190
rect 126780 663950 126870 664190
rect 127110 663950 127200 664190
rect 127440 663950 127550 664190
rect 127790 663950 127880 664190
rect 128120 663950 128210 664190
rect 128450 663950 128540 664190
rect 128780 663950 128890 664190
rect 129130 663950 129220 664190
rect 129460 663950 129550 664190
rect 129790 663950 129880 664190
rect 130120 663950 130230 664190
rect 130470 663950 130560 664190
rect 130800 663950 130890 664190
rect 131130 663950 131220 664190
rect 131460 663950 131570 664190
rect 131810 663950 131900 664190
rect 132140 663950 132230 664190
rect 132470 663950 132560 664190
rect 132800 663950 132910 664190
rect 133150 663950 133570 664190
rect 133810 663950 133900 664190
rect 134140 663950 134230 664190
rect 134470 663950 134560 664190
rect 134800 663950 134910 664190
rect 135150 663950 135240 664190
rect 135480 663950 135570 664190
rect 135810 663950 135900 664190
rect 136140 663950 136250 664190
rect 136490 663950 136580 664190
rect 136820 663950 136910 664190
rect 137150 663950 137240 664190
rect 137480 663950 137590 664190
rect 137830 663950 137920 664190
rect 138160 663950 138250 664190
rect 138490 663950 138580 664190
rect 138820 663950 138930 664190
rect 139170 663950 139260 664190
rect 139500 663950 139590 664190
rect 139830 663950 139920 664190
rect 140160 663950 140270 664190
rect 140510 663950 140600 664190
rect 140840 663950 140930 664190
rect 141170 663950 141260 664190
rect 141500 663950 141610 664190
rect 141850 663950 141940 664190
rect 142180 663950 142270 664190
rect 142510 663950 142600 664190
rect 142840 663950 142950 664190
rect 143190 663950 143280 664190
rect 143520 663950 143610 664190
rect 143850 663950 143940 664190
rect 144180 663950 144290 664190
rect 144530 663950 144950 664190
rect 145190 663950 145280 664190
rect 145520 663950 145610 664190
rect 145850 663950 145940 664190
rect 146180 663950 146290 664190
rect 146530 663950 146620 664190
rect 146860 663950 146950 664190
rect 147190 663950 147280 664190
rect 147520 663950 147630 664190
rect 147870 663950 147960 664190
rect 148200 663950 148290 664190
rect 148530 663950 148620 664190
rect 148860 663950 148970 664190
rect 149210 663950 149300 664190
rect 149540 663950 149630 664190
rect 149870 663950 149960 664190
rect 150200 663950 150310 664190
rect 150550 663950 150640 664190
rect 150880 663950 150970 664190
rect 151210 663950 151300 664190
rect 151540 663950 151650 664190
rect 151890 663950 151980 664190
rect 152220 663950 152310 664190
rect 152550 663950 152640 664190
rect 152880 663950 152990 664190
rect 153230 663950 153320 664190
rect 153560 663950 153650 664190
rect 153890 663950 153980 664190
rect 154220 663950 154330 664190
rect 154570 663950 154660 664190
rect 154900 663950 154990 664190
rect 155230 663950 155320 664190
rect 155560 663950 155670 664190
rect 155910 663950 164457 664190
rect 2500 663860 164457 663950
rect 2500 663620 110810 663860
rect 111050 663620 111140 663860
rect 111380 663620 111470 663860
rect 111710 663620 111800 663860
rect 112040 663620 112150 663860
rect 112390 663620 112480 663860
rect 112720 663620 112810 663860
rect 113050 663620 113140 663860
rect 113380 663620 113490 663860
rect 113730 663620 113820 663860
rect 114060 663620 114150 663860
rect 114390 663620 114480 663860
rect 114720 663620 114830 663860
rect 115070 663620 115160 663860
rect 115400 663620 115490 663860
rect 115730 663620 115820 663860
rect 116060 663620 116170 663860
rect 116410 663620 116500 663860
rect 116740 663620 116830 663860
rect 117070 663620 117160 663860
rect 117400 663620 117510 663860
rect 117750 663620 117840 663860
rect 118080 663620 118170 663860
rect 118410 663620 118500 663860
rect 118740 663620 118850 663860
rect 119090 663620 119180 663860
rect 119420 663620 119510 663860
rect 119750 663620 119840 663860
rect 120080 663620 120190 663860
rect 120430 663620 120520 663860
rect 120760 663620 120850 663860
rect 121090 663620 121180 663860
rect 121420 663620 121530 663860
rect 121770 663620 122190 663860
rect 122430 663620 122520 663860
rect 122760 663620 122850 663860
rect 123090 663620 123180 663860
rect 123420 663620 123530 663860
rect 123770 663620 123860 663860
rect 124100 663620 124190 663860
rect 124430 663620 124520 663860
rect 124760 663620 124870 663860
rect 125110 663620 125200 663860
rect 125440 663620 125530 663860
rect 125770 663620 125860 663860
rect 126100 663620 126210 663860
rect 126450 663620 126540 663860
rect 126780 663620 126870 663860
rect 127110 663620 127200 663860
rect 127440 663620 127550 663860
rect 127790 663620 127880 663860
rect 128120 663620 128210 663860
rect 128450 663620 128540 663860
rect 128780 663620 128890 663860
rect 129130 663620 129220 663860
rect 129460 663620 129550 663860
rect 129790 663620 129880 663860
rect 130120 663620 130230 663860
rect 130470 663620 130560 663860
rect 130800 663620 130890 663860
rect 131130 663620 131220 663860
rect 131460 663620 131570 663860
rect 131810 663620 131900 663860
rect 132140 663620 132230 663860
rect 132470 663620 132560 663860
rect 132800 663620 132910 663860
rect 133150 663620 133570 663860
rect 133810 663620 133900 663860
rect 134140 663620 134230 663860
rect 134470 663620 134560 663860
rect 134800 663620 134910 663860
rect 135150 663620 135240 663860
rect 135480 663620 135570 663860
rect 135810 663620 135900 663860
rect 136140 663620 136250 663860
rect 136490 663620 136580 663860
rect 136820 663620 136910 663860
rect 137150 663620 137240 663860
rect 137480 663620 137590 663860
rect 137830 663620 137920 663860
rect 138160 663620 138250 663860
rect 138490 663620 138580 663860
rect 138820 663620 138930 663860
rect 139170 663620 139260 663860
rect 139500 663620 139590 663860
rect 139830 663620 139920 663860
rect 140160 663620 140270 663860
rect 140510 663620 140600 663860
rect 140840 663620 140930 663860
rect 141170 663620 141260 663860
rect 141500 663620 141610 663860
rect 141850 663620 141940 663860
rect 142180 663620 142270 663860
rect 142510 663620 142600 663860
rect 142840 663620 142950 663860
rect 143190 663620 143280 663860
rect 143520 663620 143610 663860
rect 143850 663620 143940 663860
rect 144180 663620 144290 663860
rect 144530 663620 144950 663860
rect 145190 663620 145280 663860
rect 145520 663620 145610 663860
rect 145850 663620 145940 663860
rect 146180 663620 146290 663860
rect 146530 663620 146620 663860
rect 146860 663620 146950 663860
rect 147190 663620 147280 663860
rect 147520 663620 147630 663860
rect 147870 663620 147960 663860
rect 148200 663620 148290 663860
rect 148530 663620 148620 663860
rect 148860 663620 148970 663860
rect 149210 663620 149300 663860
rect 149540 663620 149630 663860
rect 149870 663620 149960 663860
rect 150200 663620 150310 663860
rect 150550 663620 150640 663860
rect 150880 663620 150970 663860
rect 151210 663620 151300 663860
rect 151540 663620 151650 663860
rect 151890 663620 151980 663860
rect 152220 663620 152310 663860
rect 152550 663620 152640 663860
rect 152880 663620 152990 663860
rect 153230 663620 153320 663860
rect 153560 663620 153650 663860
rect 153890 663620 153980 663860
rect 154220 663620 154330 663860
rect 154570 663620 154660 663860
rect 154900 663620 154990 663860
rect 155230 663620 155320 663860
rect 155560 663620 155670 663860
rect 155910 663620 164457 663860
rect 2500 663510 164457 663620
rect 2500 663270 110810 663510
rect 111050 663270 111140 663510
rect 111380 663270 111470 663510
rect 111710 663270 111800 663510
rect 112040 663270 112150 663510
rect 112390 663270 112480 663510
rect 112720 663270 112810 663510
rect 113050 663270 113140 663510
rect 113380 663270 113490 663510
rect 113730 663270 113820 663510
rect 114060 663270 114150 663510
rect 114390 663270 114480 663510
rect 114720 663270 114830 663510
rect 115070 663270 115160 663510
rect 115400 663270 115490 663510
rect 115730 663270 115820 663510
rect 116060 663270 116170 663510
rect 116410 663270 116500 663510
rect 116740 663270 116830 663510
rect 117070 663270 117160 663510
rect 117400 663270 117510 663510
rect 117750 663270 117840 663510
rect 118080 663270 118170 663510
rect 118410 663270 118500 663510
rect 118740 663270 118850 663510
rect 119090 663270 119180 663510
rect 119420 663270 119510 663510
rect 119750 663270 119840 663510
rect 120080 663270 120190 663510
rect 120430 663270 120520 663510
rect 120760 663270 120850 663510
rect 121090 663270 121180 663510
rect 121420 663270 121530 663510
rect 121770 663270 122190 663510
rect 122430 663270 122520 663510
rect 122760 663270 122850 663510
rect 123090 663270 123180 663510
rect 123420 663270 123530 663510
rect 123770 663270 123860 663510
rect 124100 663270 124190 663510
rect 124430 663270 124520 663510
rect 124760 663270 124870 663510
rect 125110 663270 125200 663510
rect 125440 663270 125530 663510
rect 125770 663270 125860 663510
rect 126100 663270 126210 663510
rect 126450 663270 126540 663510
rect 126780 663270 126870 663510
rect 127110 663270 127200 663510
rect 127440 663270 127550 663510
rect 127790 663270 127880 663510
rect 128120 663270 128210 663510
rect 128450 663270 128540 663510
rect 128780 663270 128890 663510
rect 129130 663270 129220 663510
rect 129460 663270 129550 663510
rect 129790 663270 129880 663510
rect 130120 663270 130230 663510
rect 130470 663270 130560 663510
rect 130800 663270 130890 663510
rect 131130 663270 131220 663510
rect 131460 663270 131570 663510
rect 131810 663270 131900 663510
rect 132140 663270 132230 663510
rect 132470 663270 132560 663510
rect 132800 663270 132910 663510
rect 133150 663270 133570 663510
rect 133810 663270 133900 663510
rect 134140 663270 134230 663510
rect 134470 663270 134560 663510
rect 134800 663270 134910 663510
rect 135150 663270 135240 663510
rect 135480 663270 135570 663510
rect 135810 663270 135900 663510
rect 136140 663270 136250 663510
rect 136490 663270 136580 663510
rect 136820 663270 136910 663510
rect 137150 663270 137240 663510
rect 137480 663270 137590 663510
rect 137830 663270 137920 663510
rect 138160 663270 138250 663510
rect 138490 663270 138580 663510
rect 138820 663270 138930 663510
rect 139170 663270 139260 663510
rect 139500 663270 139590 663510
rect 139830 663270 139920 663510
rect 140160 663270 140270 663510
rect 140510 663270 140600 663510
rect 140840 663270 140930 663510
rect 141170 663270 141260 663510
rect 141500 663270 141610 663510
rect 141850 663270 141940 663510
rect 142180 663270 142270 663510
rect 142510 663270 142600 663510
rect 142840 663270 142950 663510
rect 143190 663270 143280 663510
rect 143520 663270 143610 663510
rect 143850 663270 143940 663510
rect 144180 663270 144290 663510
rect 144530 663270 144950 663510
rect 145190 663270 145280 663510
rect 145520 663270 145610 663510
rect 145850 663270 145940 663510
rect 146180 663270 146290 663510
rect 146530 663270 146620 663510
rect 146860 663270 146950 663510
rect 147190 663270 147280 663510
rect 147520 663270 147630 663510
rect 147870 663270 147960 663510
rect 148200 663270 148290 663510
rect 148530 663270 148620 663510
rect 148860 663270 148970 663510
rect 149210 663270 149300 663510
rect 149540 663270 149630 663510
rect 149870 663270 149960 663510
rect 150200 663270 150310 663510
rect 150550 663270 150640 663510
rect 150880 663270 150970 663510
rect 151210 663270 151300 663510
rect 151540 663270 151650 663510
rect 151890 663270 151980 663510
rect 152220 663270 152310 663510
rect 152550 663270 152640 663510
rect 152880 663270 152990 663510
rect 153230 663270 153320 663510
rect 153560 663270 153650 663510
rect 153890 663270 153980 663510
rect 154220 663270 154330 663510
rect 154570 663270 154660 663510
rect 154900 663270 154990 663510
rect 155230 663270 155320 663510
rect 155560 663270 155670 663510
rect 155910 663270 164457 663510
rect 2500 663180 164457 663270
rect 2500 662940 110810 663180
rect 111050 662940 111140 663180
rect 111380 662940 111470 663180
rect 111710 662940 111800 663180
rect 112040 662940 112150 663180
rect 112390 662940 112480 663180
rect 112720 662940 112810 663180
rect 113050 662940 113140 663180
rect 113380 662940 113490 663180
rect 113730 662940 113820 663180
rect 114060 662940 114150 663180
rect 114390 662940 114480 663180
rect 114720 662940 114830 663180
rect 115070 662940 115160 663180
rect 115400 662940 115490 663180
rect 115730 662940 115820 663180
rect 116060 662940 116170 663180
rect 116410 662940 116500 663180
rect 116740 662940 116830 663180
rect 117070 662940 117160 663180
rect 117400 662940 117510 663180
rect 117750 662940 117840 663180
rect 118080 662940 118170 663180
rect 118410 662940 118500 663180
rect 118740 662940 118850 663180
rect 119090 662940 119180 663180
rect 119420 662940 119510 663180
rect 119750 662940 119840 663180
rect 120080 662940 120190 663180
rect 120430 662940 120520 663180
rect 120760 662940 120850 663180
rect 121090 662940 121180 663180
rect 121420 662940 121530 663180
rect 121770 662940 122190 663180
rect 122430 662940 122520 663180
rect 122760 662940 122850 663180
rect 123090 662940 123180 663180
rect 123420 662940 123530 663180
rect 123770 662940 123860 663180
rect 124100 662940 124190 663180
rect 124430 662940 124520 663180
rect 124760 662940 124870 663180
rect 125110 662940 125200 663180
rect 125440 662940 125530 663180
rect 125770 662940 125860 663180
rect 126100 662940 126210 663180
rect 126450 662940 126540 663180
rect 126780 662940 126870 663180
rect 127110 662940 127200 663180
rect 127440 662940 127550 663180
rect 127790 662940 127880 663180
rect 128120 662940 128210 663180
rect 128450 662940 128540 663180
rect 128780 662940 128890 663180
rect 129130 662940 129220 663180
rect 129460 662940 129550 663180
rect 129790 662940 129880 663180
rect 130120 662940 130230 663180
rect 130470 662940 130560 663180
rect 130800 662940 130890 663180
rect 131130 662940 131220 663180
rect 131460 662940 131570 663180
rect 131810 662940 131900 663180
rect 132140 662940 132230 663180
rect 132470 662940 132560 663180
rect 132800 662940 132910 663180
rect 133150 662940 133570 663180
rect 133810 662940 133900 663180
rect 134140 662940 134230 663180
rect 134470 662940 134560 663180
rect 134800 662940 134910 663180
rect 135150 662940 135240 663180
rect 135480 662940 135570 663180
rect 135810 662940 135900 663180
rect 136140 662940 136250 663180
rect 136490 662940 136580 663180
rect 136820 662940 136910 663180
rect 137150 662940 137240 663180
rect 137480 662940 137590 663180
rect 137830 662940 137920 663180
rect 138160 662940 138250 663180
rect 138490 662940 138580 663180
rect 138820 662940 138930 663180
rect 139170 662940 139260 663180
rect 139500 662940 139590 663180
rect 139830 662940 139920 663180
rect 140160 662940 140270 663180
rect 140510 662940 140600 663180
rect 140840 662940 140930 663180
rect 141170 662940 141260 663180
rect 141500 662940 141610 663180
rect 141850 662940 141940 663180
rect 142180 662940 142270 663180
rect 142510 662940 142600 663180
rect 142840 662940 142950 663180
rect 143190 662940 143280 663180
rect 143520 662940 143610 663180
rect 143850 662940 143940 663180
rect 144180 662940 144290 663180
rect 144530 662940 144950 663180
rect 145190 662940 145280 663180
rect 145520 662940 145610 663180
rect 145850 662940 145940 663180
rect 146180 662940 146290 663180
rect 146530 662940 146620 663180
rect 146860 662940 146950 663180
rect 147190 662940 147280 663180
rect 147520 662940 147630 663180
rect 147870 662940 147960 663180
rect 148200 662940 148290 663180
rect 148530 662940 148620 663180
rect 148860 662940 148970 663180
rect 149210 662940 149300 663180
rect 149540 662940 149630 663180
rect 149870 662940 149960 663180
rect 150200 662940 150310 663180
rect 150550 662940 150640 663180
rect 150880 662940 150970 663180
rect 151210 662940 151300 663180
rect 151540 662940 151650 663180
rect 151890 662940 151980 663180
rect 152220 662940 152310 663180
rect 152550 662940 152640 663180
rect 152880 662940 152990 663180
rect 153230 662940 153320 663180
rect 153560 662940 153650 663180
rect 153890 662940 153980 663180
rect 154220 662940 154330 663180
rect 154570 662940 154660 663180
rect 154900 662940 154990 663180
rect 155230 662940 155320 663180
rect 155560 662940 155670 663180
rect 155910 662940 164457 663180
rect 2500 662850 164457 662940
rect 2500 662610 110810 662850
rect 111050 662610 111140 662850
rect 111380 662610 111470 662850
rect 111710 662610 111800 662850
rect 112040 662610 112150 662850
rect 112390 662610 112480 662850
rect 112720 662610 112810 662850
rect 113050 662610 113140 662850
rect 113380 662610 113490 662850
rect 113730 662610 113820 662850
rect 114060 662610 114150 662850
rect 114390 662610 114480 662850
rect 114720 662610 114830 662850
rect 115070 662610 115160 662850
rect 115400 662610 115490 662850
rect 115730 662610 115820 662850
rect 116060 662610 116170 662850
rect 116410 662610 116500 662850
rect 116740 662610 116830 662850
rect 117070 662610 117160 662850
rect 117400 662610 117510 662850
rect 117750 662610 117840 662850
rect 118080 662610 118170 662850
rect 118410 662610 118500 662850
rect 118740 662610 118850 662850
rect 119090 662610 119180 662850
rect 119420 662610 119510 662850
rect 119750 662610 119840 662850
rect 120080 662610 120190 662850
rect 120430 662610 120520 662850
rect 120760 662610 120850 662850
rect 121090 662610 121180 662850
rect 121420 662610 121530 662850
rect 121770 662610 122190 662850
rect 122430 662610 122520 662850
rect 122760 662610 122850 662850
rect 123090 662610 123180 662850
rect 123420 662610 123530 662850
rect 123770 662610 123860 662850
rect 124100 662610 124190 662850
rect 124430 662610 124520 662850
rect 124760 662610 124870 662850
rect 125110 662610 125200 662850
rect 125440 662610 125530 662850
rect 125770 662610 125860 662850
rect 126100 662610 126210 662850
rect 126450 662610 126540 662850
rect 126780 662610 126870 662850
rect 127110 662610 127200 662850
rect 127440 662610 127550 662850
rect 127790 662610 127880 662850
rect 128120 662610 128210 662850
rect 128450 662610 128540 662850
rect 128780 662610 128890 662850
rect 129130 662610 129220 662850
rect 129460 662610 129550 662850
rect 129790 662610 129880 662850
rect 130120 662610 130230 662850
rect 130470 662610 130560 662850
rect 130800 662610 130890 662850
rect 131130 662610 131220 662850
rect 131460 662610 131570 662850
rect 131810 662610 131900 662850
rect 132140 662610 132230 662850
rect 132470 662610 132560 662850
rect 132800 662610 132910 662850
rect 133150 662610 133570 662850
rect 133810 662610 133900 662850
rect 134140 662610 134230 662850
rect 134470 662610 134560 662850
rect 134800 662610 134910 662850
rect 135150 662610 135240 662850
rect 135480 662610 135570 662850
rect 135810 662610 135900 662850
rect 136140 662610 136250 662850
rect 136490 662610 136580 662850
rect 136820 662610 136910 662850
rect 137150 662610 137240 662850
rect 137480 662610 137590 662850
rect 137830 662610 137920 662850
rect 138160 662610 138250 662850
rect 138490 662610 138580 662850
rect 138820 662610 138930 662850
rect 139170 662610 139260 662850
rect 139500 662610 139590 662850
rect 139830 662610 139920 662850
rect 140160 662610 140270 662850
rect 140510 662610 140600 662850
rect 140840 662610 140930 662850
rect 141170 662610 141260 662850
rect 141500 662610 141610 662850
rect 141850 662610 141940 662850
rect 142180 662610 142270 662850
rect 142510 662610 142600 662850
rect 142840 662610 142950 662850
rect 143190 662610 143280 662850
rect 143520 662610 143610 662850
rect 143850 662610 143940 662850
rect 144180 662610 144290 662850
rect 144530 662610 144950 662850
rect 145190 662610 145280 662850
rect 145520 662610 145610 662850
rect 145850 662610 145940 662850
rect 146180 662610 146290 662850
rect 146530 662610 146620 662850
rect 146860 662610 146950 662850
rect 147190 662610 147280 662850
rect 147520 662610 147630 662850
rect 147870 662610 147960 662850
rect 148200 662610 148290 662850
rect 148530 662610 148620 662850
rect 148860 662610 148970 662850
rect 149210 662610 149300 662850
rect 149540 662610 149630 662850
rect 149870 662610 149960 662850
rect 150200 662610 150310 662850
rect 150550 662610 150640 662850
rect 150880 662610 150970 662850
rect 151210 662610 151300 662850
rect 151540 662610 151650 662850
rect 151890 662610 151980 662850
rect 152220 662610 152310 662850
rect 152550 662610 152640 662850
rect 152880 662610 152990 662850
rect 153230 662610 153320 662850
rect 153560 662610 153650 662850
rect 153890 662610 153980 662850
rect 154220 662610 154330 662850
rect 154570 662610 154660 662850
rect 154900 662610 154990 662850
rect 155230 662610 155320 662850
rect 155560 662610 155670 662850
rect 155910 662610 164457 662850
rect 2500 662520 164457 662610
rect 2500 662280 110810 662520
rect 111050 662280 111140 662520
rect 111380 662280 111470 662520
rect 111710 662280 111800 662520
rect 112040 662280 112150 662520
rect 112390 662280 112480 662520
rect 112720 662280 112810 662520
rect 113050 662280 113140 662520
rect 113380 662280 113490 662520
rect 113730 662280 113820 662520
rect 114060 662280 114150 662520
rect 114390 662280 114480 662520
rect 114720 662280 114830 662520
rect 115070 662280 115160 662520
rect 115400 662280 115490 662520
rect 115730 662280 115820 662520
rect 116060 662280 116170 662520
rect 116410 662280 116500 662520
rect 116740 662280 116830 662520
rect 117070 662280 117160 662520
rect 117400 662280 117510 662520
rect 117750 662280 117840 662520
rect 118080 662280 118170 662520
rect 118410 662280 118500 662520
rect 118740 662280 118850 662520
rect 119090 662280 119180 662520
rect 119420 662280 119510 662520
rect 119750 662280 119840 662520
rect 120080 662280 120190 662520
rect 120430 662280 120520 662520
rect 120760 662280 120850 662520
rect 121090 662280 121180 662520
rect 121420 662280 121530 662520
rect 121770 662280 122190 662520
rect 122430 662280 122520 662520
rect 122760 662280 122850 662520
rect 123090 662280 123180 662520
rect 123420 662280 123530 662520
rect 123770 662280 123860 662520
rect 124100 662280 124190 662520
rect 124430 662280 124520 662520
rect 124760 662280 124870 662520
rect 125110 662280 125200 662520
rect 125440 662280 125530 662520
rect 125770 662280 125860 662520
rect 126100 662280 126210 662520
rect 126450 662280 126540 662520
rect 126780 662280 126870 662520
rect 127110 662280 127200 662520
rect 127440 662280 127550 662520
rect 127790 662280 127880 662520
rect 128120 662280 128210 662520
rect 128450 662280 128540 662520
rect 128780 662280 128890 662520
rect 129130 662280 129220 662520
rect 129460 662280 129550 662520
rect 129790 662280 129880 662520
rect 130120 662280 130230 662520
rect 130470 662280 130560 662520
rect 130800 662280 130890 662520
rect 131130 662280 131220 662520
rect 131460 662280 131570 662520
rect 131810 662280 131900 662520
rect 132140 662280 132230 662520
rect 132470 662280 132560 662520
rect 132800 662280 132910 662520
rect 133150 662280 133570 662520
rect 133810 662280 133900 662520
rect 134140 662280 134230 662520
rect 134470 662280 134560 662520
rect 134800 662280 134910 662520
rect 135150 662280 135240 662520
rect 135480 662280 135570 662520
rect 135810 662280 135900 662520
rect 136140 662280 136250 662520
rect 136490 662280 136580 662520
rect 136820 662280 136910 662520
rect 137150 662280 137240 662520
rect 137480 662280 137590 662520
rect 137830 662280 137920 662520
rect 138160 662280 138250 662520
rect 138490 662280 138580 662520
rect 138820 662280 138930 662520
rect 139170 662280 139260 662520
rect 139500 662280 139590 662520
rect 139830 662280 139920 662520
rect 140160 662280 140270 662520
rect 140510 662280 140600 662520
rect 140840 662280 140930 662520
rect 141170 662280 141260 662520
rect 141500 662280 141610 662520
rect 141850 662280 141940 662520
rect 142180 662280 142270 662520
rect 142510 662280 142600 662520
rect 142840 662280 142950 662520
rect 143190 662280 143280 662520
rect 143520 662280 143610 662520
rect 143850 662280 143940 662520
rect 144180 662280 144290 662520
rect 144530 662280 144950 662520
rect 145190 662280 145280 662520
rect 145520 662280 145610 662520
rect 145850 662280 145940 662520
rect 146180 662280 146290 662520
rect 146530 662280 146620 662520
rect 146860 662280 146950 662520
rect 147190 662280 147280 662520
rect 147520 662280 147630 662520
rect 147870 662280 147960 662520
rect 148200 662280 148290 662520
rect 148530 662280 148620 662520
rect 148860 662280 148970 662520
rect 149210 662280 149300 662520
rect 149540 662280 149630 662520
rect 149870 662280 149960 662520
rect 150200 662280 150310 662520
rect 150550 662280 150640 662520
rect 150880 662280 150970 662520
rect 151210 662280 151300 662520
rect 151540 662280 151650 662520
rect 151890 662280 151980 662520
rect 152220 662280 152310 662520
rect 152550 662280 152640 662520
rect 152880 662280 152990 662520
rect 153230 662280 153320 662520
rect 153560 662280 153650 662520
rect 153890 662280 153980 662520
rect 154220 662280 154330 662520
rect 154570 662280 154660 662520
rect 154900 662280 154990 662520
rect 155230 662280 155320 662520
rect 155560 662280 155670 662520
rect 155910 662280 164457 662520
rect 2500 662170 164457 662280
rect 2500 661930 110810 662170
rect 111050 661930 111140 662170
rect 111380 661930 111470 662170
rect 111710 661930 111800 662170
rect 112040 661930 112150 662170
rect 112390 661930 112480 662170
rect 112720 661930 112810 662170
rect 113050 661930 113140 662170
rect 113380 661930 113490 662170
rect 113730 661930 113820 662170
rect 114060 661930 114150 662170
rect 114390 661930 114480 662170
rect 114720 661930 114830 662170
rect 115070 661930 115160 662170
rect 115400 661930 115490 662170
rect 115730 661930 115820 662170
rect 116060 661930 116170 662170
rect 116410 661930 116500 662170
rect 116740 661930 116830 662170
rect 117070 661930 117160 662170
rect 117400 661930 117510 662170
rect 117750 661930 117840 662170
rect 118080 661930 118170 662170
rect 118410 661930 118500 662170
rect 118740 661930 118850 662170
rect 119090 661930 119180 662170
rect 119420 661930 119510 662170
rect 119750 661930 119840 662170
rect 120080 661930 120190 662170
rect 120430 661930 120520 662170
rect 120760 661930 120850 662170
rect 121090 661930 121180 662170
rect 121420 661930 121530 662170
rect 121770 661930 122190 662170
rect 122430 661930 122520 662170
rect 122760 661930 122850 662170
rect 123090 661930 123180 662170
rect 123420 661930 123530 662170
rect 123770 661930 123860 662170
rect 124100 661930 124190 662170
rect 124430 661930 124520 662170
rect 124760 661930 124870 662170
rect 125110 661930 125200 662170
rect 125440 661930 125530 662170
rect 125770 661930 125860 662170
rect 126100 661930 126210 662170
rect 126450 661930 126540 662170
rect 126780 661930 126870 662170
rect 127110 661930 127200 662170
rect 127440 661930 127550 662170
rect 127790 661930 127880 662170
rect 128120 661930 128210 662170
rect 128450 661930 128540 662170
rect 128780 661930 128890 662170
rect 129130 661930 129220 662170
rect 129460 661930 129550 662170
rect 129790 661930 129880 662170
rect 130120 661930 130230 662170
rect 130470 661930 130560 662170
rect 130800 661930 130890 662170
rect 131130 661930 131220 662170
rect 131460 661930 131570 662170
rect 131810 661930 131900 662170
rect 132140 661930 132230 662170
rect 132470 661930 132560 662170
rect 132800 661930 132910 662170
rect 133150 661930 133570 662170
rect 133810 661930 133900 662170
rect 134140 661930 134230 662170
rect 134470 661930 134560 662170
rect 134800 661930 134910 662170
rect 135150 661930 135240 662170
rect 135480 661930 135570 662170
rect 135810 661930 135900 662170
rect 136140 661930 136250 662170
rect 136490 661930 136580 662170
rect 136820 661930 136910 662170
rect 137150 661930 137240 662170
rect 137480 661930 137590 662170
rect 137830 661930 137920 662170
rect 138160 661930 138250 662170
rect 138490 661930 138580 662170
rect 138820 661930 138930 662170
rect 139170 661930 139260 662170
rect 139500 661930 139590 662170
rect 139830 661930 139920 662170
rect 140160 661930 140270 662170
rect 140510 661930 140600 662170
rect 140840 661930 140930 662170
rect 141170 661930 141260 662170
rect 141500 661930 141610 662170
rect 141850 661930 141940 662170
rect 142180 661930 142270 662170
rect 142510 661930 142600 662170
rect 142840 661930 142950 662170
rect 143190 661930 143280 662170
rect 143520 661930 143610 662170
rect 143850 661930 143940 662170
rect 144180 661930 144290 662170
rect 144530 661930 144950 662170
rect 145190 661930 145280 662170
rect 145520 661930 145610 662170
rect 145850 661930 145940 662170
rect 146180 661930 146290 662170
rect 146530 661930 146620 662170
rect 146860 661930 146950 662170
rect 147190 661930 147280 662170
rect 147520 661930 147630 662170
rect 147870 661930 147960 662170
rect 148200 661930 148290 662170
rect 148530 661930 148620 662170
rect 148860 661930 148970 662170
rect 149210 661930 149300 662170
rect 149540 661930 149630 662170
rect 149870 661930 149960 662170
rect 150200 661930 150310 662170
rect 150550 661930 150640 662170
rect 150880 661930 150970 662170
rect 151210 661930 151300 662170
rect 151540 661930 151650 662170
rect 151890 661930 151980 662170
rect 152220 661930 152310 662170
rect 152550 661930 152640 662170
rect 152880 661930 152990 662170
rect 153230 661930 153320 662170
rect 153560 661930 153650 662170
rect 153890 661930 153980 662170
rect 154220 661930 154330 662170
rect 154570 661930 154660 662170
rect 154900 661930 154990 662170
rect 155230 661930 155320 662170
rect 155560 661930 155670 662170
rect 155910 661930 164457 662170
rect 2500 661840 164457 661930
rect 2500 661600 110810 661840
rect 111050 661600 111140 661840
rect 111380 661600 111470 661840
rect 111710 661600 111800 661840
rect 112040 661600 112150 661840
rect 112390 661600 112480 661840
rect 112720 661600 112810 661840
rect 113050 661600 113140 661840
rect 113380 661600 113490 661840
rect 113730 661600 113820 661840
rect 114060 661600 114150 661840
rect 114390 661600 114480 661840
rect 114720 661600 114830 661840
rect 115070 661600 115160 661840
rect 115400 661600 115490 661840
rect 115730 661600 115820 661840
rect 116060 661600 116170 661840
rect 116410 661600 116500 661840
rect 116740 661600 116830 661840
rect 117070 661600 117160 661840
rect 117400 661600 117510 661840
rect 117750 661600 117840 661840
rect 118080 661600 118170 661840
rect 118410 661600 118500 661840
rect 118740 661600 118850 661840
rect 119090 661600 119180 661840
rect 119420 661600 119510 661840
rect 119750 661600 119840 661840
rect 120080 661600 120190 661840
rect 120430 661600 120520 661840
rect 120760 661600 120850 661840
rect 121090 661600 121180 661840
rect 121420 661600 121530 661840
rect 121770 661600 122190 661840
rect 122430 661600 122520 661840
rect 122760 661600 122850 661840
rect 123090 661600 123180 661840
rect 123420 661600 123530 661840
rect 123770 661600 123860 661840
rect 124100 661600 124190 661840
rect 124430 661600 124520 661840
rect 124760 661600 124870 661840
rect 125110 661600 125200 661840
rect 125440 661600 125530 661840
rect 125770 661600 125860 661840
rect 126100 661600 126210 661840
rect 126450 661600 126540 661840
rect 126780 661600 126870 661840
rect 127110 661600 127200 661840
rect 127440 661600 127550 661840
rect 127790 661600 127880 661840
rect 128120 661600 128210 661840
rect 128450 661600 128540 661840
rect 128780 661600 128890 661840
rect 129130 661600 129220 661840
rect 129460 661600 129550 661840
rect 129790 661600 129880 661840
rect 130120 661600 130230 661840
rect 130470 661600 130560 661840
rect 130800 661600 130890 661840
rect 131130 661600 131220 661840
rect 131460 661600 131570 661840
rect 131810 661600 131900 661840
rect 132140 661600 132230 661840
rect 132470 661600 132560 661840
rect 132800 661600 132910 661840
rect 133150 661600 133570 661840
rect 133810 661600 133900 661840
rect 134140 661600 134230 661840
rect 134470 661600 134560 661840
rect 134800 661600 134910 661840
rect 135150 661600 135240 661840
rect 135480 661600 135570 661840
rect 135810 661600 135900 661840
rect 136140 661600 136250 661840
rect 136490 661600 136580 661840
rect 136820 661600 136910 661840
rect 137150 661600 137240 661840
rect 137480 661600 137590 661840
rect 137830 661600 137920 661840
rect 138160 661600 138250 661840
rect 138490 661600 138580 661840
rect 138820 661600 138930 661840
rect 139170 661600 139260 661840
rect 139500 661600 139590 661840
rect 139830 661600 139920 661840
rect 140160 661600 140270 661840
rect 140510 661600 140600 661840
rect 140840 661600 140930 661840
rect 141170 661600 141260 661840
rect 141500 661600 141610 661840
rect 141850 661600 141940 661840
rect 142180 661600 142270 661840
rect 142510 661600 142600 661840
rect 142840 661600 142950 661840
rect 143190 661600 143280 661840
rect 143520 661600 143610 661840
rect 143850 661600 143940 661840
rect 144180 661600 144290 661840
rect 144530 661600 144950 661840
rect 145190 661600 145280 661840
rect 145520 661600 145610 661840
rect 145850 661600 145940 661840
rect 146180 661600 146290 661840
rect 146530 661600 146620 661840
rect 146860 661600 146950 661840
rect 147190 661600 147280 661840
rect 147520 661600 147630 661840
rect 147870 661600 147960 661840
rect 148200 661600 148290 661840
rect 148530 661600 148620 661840
rect 148860 661600 148970 661840
rect 149210 661600 149300 661840
rect 149540 661600 149630 661840
rect 149870 661600 149960 661840
rect 150200 661600 150310 661840
rect 150550 661600 150640 661840
rect 150880 661600 150970 661840
rect 151210 661600 151300 661840
rect 151540 661600 151650 661840
rect 151890 661600 151980 661840
rect 152220 661600 152310 661840
rect 152550 661600 152640 661840
rect 152880 661600 152990 661840
rect 153230 661600 153320 661840
rect 153560 661600 153650 661840
rect 153890 661600 153980 661840
rect 154220 661600 154330 661840
rect 154570 661600 154660 661840
rect 154900 661600 154990 661840
rect 155230 661600 155320 661840
rect 155560 661600 155670 661840
rect 155910 661600 164457 661840
rect 2500 661510 164457 661600
rect 2500 661270 110810 661510
rect 111050 661270 111140 661510
rect 111380 661270 111470 661510
rect 111710 661270 111800 661510
rect 112040 661270 112150 661510
rect 112390 661270 112480 661510
rect 112720 661270 112810 661510
rect 113050 661270 113140 661510
rect 113380 661270 113490 661510
rect 113730 661270 113820 661510
rect 114060 661270 114150 661510
rect 114390 661270 114480 661510
rect 114720 661270 114830 661510
rect 115070 661270 115160 661510
rect 115400 661270 115490 661510
rect 115730 661270 115820 661510
rect 116060 661270 116170 661510
rect 116410 661270 116500 661510
rect 116740 661270 116830 661510
rect 117070 661270 117160 661510
rect 117400 661270 117510 661510
rect 117750 661270 117840 661510
rect 118080 661270 118170 661510
rect 118410 661270 118500 661510
rect 118740 661270 118850 661510
rect 119090 661270 119180 661510
rect 119420 661270 119510 661510
rect 119750 661270 119840 661510
rect 120080 661270 120190 661510
rect 120430 661270 120520 661510
rect 120760 661270 120850 661510
rect 121090 661270 121180 661510
rect 121420 661270 121530 661510
rect 121770 661270 122190 661510
rect 122430 661270 122520 661510
rect 122760 661270 122850 661510
rect 123090 661270 123180 661510
rect 123420 661270 123530 661510
rect 123770 661270 123860 661510
rect 124100 661270 124190 661510
rect 124430 661270 124520 661510
rect 124760 661270 124870 661510
rect 125110 661270 125200 661510
rect 125440 661270 125530 661510
rect 125770 661270 125860 661510
rect 126100 661270 126210 661510
rect 126450 661270 126540 661510
rect 126780 661270 126870 661510
rect 127110 661270 127200 661510
rect 127440 661270 127550 661510
rect 127790 661270 127880 661510
rect 128120 661270 128210 661510
rect 128450 661270 128540 661510
rect 128780 661270 128890 661510
rect 129130 661270 129220 661510
rect 129460 661270 129550 661510
rect 129790 661270 129880 661510
rect 130120 661270 130230 661510
rect 130470 661270 130560 661510
rect 130800 661270 130890 661510
rect 131130 661270 131220 661510
rect 131460 661270 131570 661510
rect 131810 661270 131900 661510
rect 132140 661270 132230 661510
rect 132470 661270 132560 661510
rect 132800 661270 132910 661510
rect 133150 661270 133570 661510
rect 133810 661270 133900 661510
rect 134140 661270 134230 661510
rect 134470 661270 134560 661510
rect 134800 661270 134910 661510
rect 135150 661270 135240 661510
rect 135480 661270 135570 661510
rect 135810 661270 135900 661510
rect 136140 661270 136250 661510
rect 136490 661270 136580 661510
rect 136820 661270 136910 661510
rect 137150 661270 137240 661510
rect 137480 661270 137590 661510
rect 137830 661270 137920 661510
rect 138160 661270 138250 661510
rect 138490 661270 138580 661510
rect 138820 661270 138930 661510
rect 139170 661270 139260 661510
rect 139500 661270 139590 661510
rect 139830 661270 139920 661510
rect 140160 661270 140270 661510
rect 140510 661270 140600 661510
rect 140840 661270 140930 661510
rect 141170 661270 141260 661510
rect 141500 661270 141610 661510
rect 141850 661270 141940 661510
rect 142180 661270 142270 661510
rect 142510 661270 142600 661510
rect 142840 661270 142950 661510
rect 143190 661270 143280 661510
rect 143520 661270 143610 661510
rect 143850 661270 143940 661510
rect 144180 661270 144290 661510
rect 144530 661270 144950 661510
rect 145190 661270 145280 661510
rect 145520 661270 145610 661510
rect 145850 661270 145940 661510
rect 146180 661270 146290 661510
rect 146530 661270 146620 661510
rect 146860 661270 146950 661510
rect 147190 661270 147280 661510
rect 147520 661270 147630 661510
rect 147870 661270 147960 661510
rect 148200 661270 148290 661510
rect 148530 661270 148620 661510
rect 148860 661270 148970 661510
rect 149210 661270 149300 661510
rect 149540 661270 149630 661510
rect 149870 661270 149960 661510
rect 150200 661270 150310 661510
rect 150550 661270 150640 661510
rect 150880 661270 150970 661510
rect 151210 661270 151300 661510
rect 151540 661270 151650 661510
rect 151890 661270 151980 661510
rect 152220 661270 152310 661510
rect 152550 661270 152640 661510
rect 152880 661270 152990 661510
rect 153230 661270 153320 661510
rect 153560 661270 153650 661510
rect 153890 661270 153980 661510
rect 154220 661270 154330 661510
rect 154570 661270 154660 661510
rect 154900 661270 154990 661510
rect 155230 661270 155320 661510
rect 155560 661270 155670 661510
rect 155910 661270 164457 661510
rect 2500 661180 164457 661270
rect 2500 660940 110810 661180
rect 111050 660940 111140 661180
rect 111380 660940 111470 661180
rect 111710 660940 111800 661180
rect 112040 660940 112150 661180
rect 112390 660940 112480 661180
rect 112720 660940 112810 661180
rect 113050 660940 113140 661180
rect 113380 660940 113490 661180
rect 113730 660940 113820 661180
rect 114060 660940 114150 661180
rect 114390 660940 114480 661180
rect 114720 660940 114830 661180
rect 115070 660940 115160 661180
rect 115400 660940 115490 661180
rect 115730 660940 115820 661180
rect 116060 660940 116170 661180
rect 116410 660940 116500 661180
rect 116740 660940 116830 661180
rect 117070 660940 117160 661180
rect 117400 660940 117510 661180
rect 117750 660940 117840 661180
rect 118080 660940 118170 661180
rect 118410 660940 118500 661180
rect 118740 660940 118850 661180
rect 119090 660940 119180 661180
rect 119420 660940 119510 661180
rect 119750 660940 119840 661180
rect 120080 660940 120190 661180
rect 120430 660940 120520 661180
rect 120760 660940 120850 661180
rect 121090 660940 121180 661180
rect 121420 660940 121530 661180
rect 121770 660940 122190 661180
rect 122430 660940 122520 661180
rect 122760 660940 122850 661180
rect 123090 660940 123180 661180
rect 123420 660940 123530 661180
rect 123770 660940 123860 661180
rect 124100 660940 124190 661180
rect 124430 660940 124520 661180
rect 124760 660940 124870 661180
rect 125110 660940 125200 661180
rect 125440 660940 125530 661180
rect 125770 660940 125860 661180
rect 126100 660940 126210 661180
rect 126450 660940 126540 661180
rect 126780 660940 126870 661180
rect 127110 660940 127200 661180
rect 127440 660940 127550 661180
rect 127790 660940 127880 661180
rect 128120 660940 128210 661180
rect 128450 660940 128540 661180
rect 128780 660940 128890 661180
rect 129130 660940 129220 661180
rect 129460 660940 129550 661180
rect 129790 660940 129880 661180
rect 130120 660940 130230 661180
rect 130470 660940 130560 661180
rect 130800 660940 130890 661180
rect 131130 660940 131220 661180
rect 131460 660940 131570 661180
rect 131810 660940 131900 661180
rect 132140 660940 132230 661180
rect 132470 660940 132560 661180
rect 132800 660940 132910 661180
rect 133150 660940 133570 661180
rect 133810 660940 133900 661180
rect 134140 660940 134230 661180
rect 134470 660940 134560 661180
rect 134800 660940 134910 661180
rect 135150 660940 135240 661180
rect 135480 660940 135570 661180
rect 135810 660940 135900 661180
rect 136140 660940 136250 661180
rect 136490 660940 136580 661180
rect 136820 660940 136910 661180
rect 137150 660940 137240 661180
rect 137480 660940 137590 661180
rect 137830 660940 137920 661180
rect 138160 660940 138250 661180
rect 138490 660940 138580 661180
rect 138820 660940 138930 661180
rect 139170 660940 139260 661180
rect 139500 660940 139590 661180
rect 139830 660940 139920 661180
rect 140160 660940 140270 661180
rect 140510 660940 140600 661180
rect 140840 660940 140930 661180
rect 141170 660940 141260 661180
rect 141500 660940 141610 661180
rect 141850 660940 141940 661180
rect 142180 660940 142270 661180
rect 142510 660940 142600 661180
rect 142840 660940 142950 661180
rect 143190 660940 143280 661180
rect 143520 660940 143610 661180
rect 143850 660940 143940 661180
rect 144180 660940 144290 661180
rect 144530 660940 144950 661180
rect 145190 660940 145280 661180
rect 145520 660940 145610 661180
rect 145850 660940 145940 661180
rect 146180 660940 146290 661180
rect 146530 660940 146620 661180
rect 146860 660940 146950 661180
rect 147190 660940 147280 661180
rect 147520 660940 147630 661180
rect 147870 660940 147960 661180
rect 148200 660940 148290 661180
rect 148530 660940 148620 661180
rect 148860 660940 148970 661180
rect 149210 660940 149300 661180
rect 149540 660940 149630 661180
rect 149870 660940 149960 661180
rect 150200 660940 150310 661180
rect 150550 660940 150640 661180
rect 150880 660940 150970 661180
rect 151210 660940 151300 661180
rect 151540 660940 151650 661180
rect 151890 660940 151980 661180
rect 152220 660940 152310 661180
rect 152550 660940 152640 661180
rect 152880 660940 152990 661180
rect 153230 660940 153320 661180
rect 153560 660940 153650 661180
rect 153890 660940 153980 661180
rect 154220 660940 154330 661180
rect 154570 660940 154660 661180
rect 154900 660940 154990 661180
rect 155230 660940 155320 661180
rect 155560 660940 155670 661180
rect 155910 660940 164457 661180
rect 2500 660760 164457 660940
rect 2500 660520 110890 660760
rect 111130 660520 111220 660760
rect 111460 660520 111550 660760
rect 111790 660520 111880 660760
rect 112120 660520 112210 660760
rect 112450 660520 112540 660760
rect 112780 660520 112870 660760
rect 113110 660520 113200 660760
rect 113440 660520 113530 660760
rect 113770 660520 113860 660760
rect 114100 660520 114190 660760
rect 114430 660520 114520 660760
rect 114760 660520 114850 660760
rect 115090 660520 115180 660760
rect 115420 660520 115510 660760
rect 115750 660520 115840 660760
rect 116080 660520 116170 660760
rect 116410 660520 116500 660760
rect 116740 660520 116830 660760
rect 117070 660520 117160 660760
rect 117400 660520 117490 660760
rect 117730 660520 117820 660760
rect 118060 660520 118150 660760
rect 118390 660520 118480 660760
rect 118720 660520 118810 660760
rect 119050 660520 119140 660760
rect 119380 660520 119470 660760
rect 119710 660520 119800 660760
rect 120040 660520 120130 660760
rect 120370 660520 120460 660760
rect 120700 660520 120790 660760
rect 121030 660520 121120 660760
rect 121360 660520 121450 660760
rect 121690 660520 122270 660760
rect 122510 660520 122600 660760
rect 122840 660520 122930 660760
rect 123170 660520 123260 660760
rect 123500 660520 123590 660760
rect 123830 660520 123920 660760
rect 124160 660520 124250 660760
rect 124490 660520 124580 660760
rect 124820 660520 124910 660760
rect 125150 660520 125240 660760
rect 125480 660520 125570 660760
rect 125810 660520 125900 660760
rect 126140 660520 126230 660760
rect 126470 660520 126560 660760
rect 126800 660520 126890 660760
rect 127130 660520 127220 660760
rect 127460 660520 127550 660760
rect 127790 660520 127880 660760
rect 128120 660520 128210 660760
rect 128450 660520 128540 660760
rect 128780 660520 128870 660760
rect 129110 660520 129200 660760
rect 129440 660520 129530 660760
rect 129770 660520 129860 660760
rect 130100 660520 130190 660760
rect 130430 660520 130520 660760
rect 130760 660520 130850 660760
rect 131090 660520 131180 660760
rect 131420 660520 131510 660760
rect 131750 660520 131840 660760
rect 132080 660520 132170 660760
rect 132410 660520 132500 660760
rect 132740 660520 132830 660760
rect 133070 660520 133650 660760
rect 133890 660520 133980 660760
rect 134220 660520 134310 660760
rect 134550 660520 134640 660760
rect 134880 660520 134970 660760
rect 135210 660520 135300 660760
rect 135540 660520 135630 660760
rect 135870 660520 135960 660760
rect 136200 660520 136290 660760
rect 136530 660520 136620 660760
rect 136860 660520 136950 660760
rect 137190 660520 137280 660760
rect 137520 660520 137610 660760
rect 137850 660520 137940 660760
rect 138180 660520 138270 660760
rect 138510 660520 138600 660760
rect 138840 660520 138930 660760
rect 139170 660520 139260 660760
rect 139500 660520 139590 660760
rect 139830 660520 139920 660760
rect 140160 660520 140250 660760
rect 140490 660520 140580 660760
rect 140820 660520 140910 660760
rect 141150 660520 141240 660760
rect 141480 660520 141570 660760
rect 141810 660520 141900 660760
rect 142140 660520 142230 660760
rect 142470 660520 142560 660760
rect 142800 660520 142890 660760
rect 143130 660520 143220 660760
rect 143460 660520 143550 660760
rect 143790 660520 143880 660760
rect 144120 660520 144210 660760
rect 144450 660520 145030 660760
rect 145270 660520 145360 660760
rect 145600 660520 145690 660760
rect 145930 660520 146020 660760
rect 146260 660520 146350 660760
rect 146590 660520 146680 660760
rect 146920 660520 147010 660760
rect 147250 660520 147340 660760
rect 147580 660520 147670 660760
rect 147910 660520 148000 660760
rect 148240 660520 148330 660760
rect 148570 660520 148660 660760
rect 148900 660520 148990 660760
rect 149230 660520 149320 660760
rect 149560 660520 149650 660760
rect 149890 660520 149980 660760
rect 150220 660520 150310 660760
rect 150550 660520 150640 660760
rect 150880 660520 150970 660760
rect 151210 660520 151300 660760
rect 151540 660520 151630 660760
rect 151870 660520 151960 660760
rect 152200 660520 152290 660760
rect 152530 660520 152620 660760
rect 152860 660520 152950 660760
rect 153190 660520 153280 660760
rect 153520 660520 153610 660760
rect 153850 660520 153940 660760
rect 154180 660520 154270 660760
rect 154510 660520 154600 660760
rect 154840 660520 154930 660760
rect 155170 660520 155260 660760
rect 155500 660520 155590 660760
rect 155830 660520 164457 660760
rect 2500 660505 164457 660520
rect 110760 660340 155960 660505
rect 110760 660100 110810 660340
rect 111050 660100 111160 660340
rect 111400 660100 111490 660340
rect 111730 660100 111820 660340
rect 112060 660100 112150 660340
rect 112390 660100 112500 660340
rect 112740 660100 112830 660340
rect 113070 660100 113160 660340
rect 113400 660100 113490 660340
rect 113730 660100 113840 660340
rect 114080 660100 114170 660340
rect 114410 660100 114500 660340
rect 114740 660100 114830 660340
rect 115070 660100 115180 660340
rect 115420 660100 115510 660340
rect 115750 660100 115840 660340
rect 116080 660100 116170 660340
rect 116410 660100 116520 660340
rect 116760 660100 116850 660340
rect 117090 660100 117180 660340
rect 117420 660100 117510 660340
rect 117750 660100 117860 660340
rect 118100 660100 118190 660340
rect 118430 660100 118520 660340
rect 118760 660100 118850 660340
rect 119090 660100 119200 660340
rect 119440 660100 119530 660340
rect 119770 660100 119860 660340
rect 120100 660100 120190 660340
rect 120430 660100 120540 660340
rect 120780 660100 120870 660340
rect 121110 660100 121200 660340
rect 121440 660100 121530 660340
rect 121770 660100 122190 660340
rect 122430 660100 122540 660340
rect 122780 660100 122870 660340
rect 123110 660100 123200 660340
rect 123440 660100 123530 660340
rect 123770 660100 123880 660340
rect 124120 660100 124210 660340
rect 124450 660100 124540 660340
rect 124780 660100 124870 660340
rect 125110 660100 125220 660340
rect 125460 660100 125550 660340
rect 125790 660100 125880 660340
rect 126120 660100 126210 660340
rect 126450 660100 126560 660340
rect 126800 660100 126890 660340
rect 127130 660100 127220 660340
rect 127460 660100 127550 660340
rect 127790 660100 127900 660340
rect 128140 660100 128230 660340
rect 128470 660100 128560 660340
rect 128800 660100 128890 660340
rect 129130 660100 129240 660340
rect 129480 660100 129570 660340
rect 129810 660100 129900 660340
rect 130140 660100 130230 660340
rect 130470 660100 130580 660340
rect 130820 660100 130910 660340
rect 131150 660100 131240 660340
rect 131480 660100 131570 660340
rect 131810 660100 131920 660340
rect 132160 660100 132250 660340
rect 132490 660100 132580 660340
rect 132820 660100 132910 660340
rect 133150 660100 133570 660340
rect 133810 660100 133920 660340
rect 134160 660100 134250 660340
rect 134490 660100 134580 660340
rect 134820 660100 134910 660340
rect 135150 660100 135260 660340
rect 135500 660100 135590 660340
rect 135830 660100 135920 660340
rect 136160 660100 136250 660340
rect 136490 660100 136600 660340
rect 136840 660100 136930 660340
rect 137170 660100 137260 660340
rect 137500 660100 137590 660340
rect 137830 660100 137940 660340
rect 138180 660100 138270 660340
rect 138510 660100 138600 660340
rect 138840 660100 138930 660340
rect 139170 660100 139280 660340
rect 139520 660100 139610 660340
rect 139850 660100 139940 660340
rect 140180 660100 140270 660340
rect 140510 660100 140620 660340
rect 140860 660100 140950 660340
rect 141190 660100 141280 660340
rect 141520 660100 141610 660340
rect 141850 660100 141960 660340
rect 142200 660100 142290 660340
rect 142530 660100 142620 660340
rect 142860 660100 142950 660340
rect 143190 660100 143300 660340
rect 143540 660100 143630 660340
rect 143870 660100 143960 660340
rect 144200 660100 144290 660340
rect 144530 660100 144950 660340
rect 145190 660100 145300 660340
rect 145540 660100 145630 660340
rect 145870 660100 145960 660340
rect 146200 660100 146290 660340
rect 146530 660100 146640 660340
rect 146880 660100 146970 660340
rect 147210 660100 147300 660340
rect 147540 660100 147630 660340
rect 147870 660100 147980 660340
rect 148220 660100 148310 660340
rect 148550 660100 148640 660340
rect 148880 660100 148970 660340
rect 149210 660100 149320 660340
rect 149560 660100 149650 660340
rect 149890 660100 149980 660340
rect 150220 660100 150310 660340
rect 150550 660100 150660 660340
rect 150900 660100 150990 660340
rect 151230 660100 151320 660340
rect 151560 660100 151650 660340
rect 151890 660100 152000 660340
rect 152240 660100 152330 660340
rect 152570 660100 152660 660340
rect 152900 660100 152990 660340
rect 153230 660100 153340 660340
rect 153580 660100 153670 660340
rect 153910 660100 154000 660340
rect 154240 660100 154330 660340
rect 154570 660100 154680 660340
rect 154920 660100 155010 660340
rect 155250 660100 155340 660340
rect 155580 660100 155670 660340
rect 155910 660100 155960 660340
rect 110760 660010 155960 660100
rect 110760 659770 110810 660010
rect 111050 659770 111160 660010
rect 111400 659770 111490 660010
rect 111730 659770 111820 660010
rect 112060 659770 112150 660010
rect 112390 659770 112500 660010
rect 112740 659770 112830 660010
rect 113070 659770 113160 660010
rect 113400 659770 113490 660010
rect 113730 659770 113840 660010
rect 114080 659770 114170 660010
rect 114410 659770 114500 660010
rect 114740 659770 114830 660010
rect 115070 659770 115180 660010
rect 115420 659770 115510 660010
rect 115750 659770 115840 660010
rect 116080 659770 116170 660010
rect 116410 659770 116520 660010
rect 116760 659770 116850 660010
rect 117090 659770 117180 660010
rect 117420 659770 117510 660010
rect 117750 659770 117860 660010
rect 118100 659770 118190 660010
rect 118430 659770 118520 660010
rect 118760 659770 118850 660010
rect 119090 659770 119200 660010
rect 119440 659770 119530 660010
rect 119770 659770 119860 660010
rect 120100 659770 120190 660010
rect 120430 659770 120540 660010
rect 120780 659770 120870 660010
rect 121110 659770 121200 660010
rect 121440 659770 121530 660010
rect 121770 659770 122190 660010
rect 122430 659770 122540 660010
rect 122780 659770 122870 660010
rect 123110 659770 123200 660010
rect 123440 659770 123530 660010
rect 123770 659770 123880 660010
rect 124120 659770 124210 660010
rect 124450 659770 124540 660010
rect 124780 659770 124870 660010
rect 125110 659770 125220 660010
rect 125460 659770 125550 660010
rect 125790 659770 125880 660010
rect 126120 659770 126210 660010
rect 126450 659770 126560 660010
rect 126800 659770 126890 660010
rect 127130 659770 127220 660010
rect 127460 659770 127550 660010
rect 127790 659770 127900 660010
rect 128140 659770 128230 660010
rect 128470 659770 128560 660010
rect 128800 659770 128890 660010
rect 129130 659770 129240 660010
rect 129480 659770 129570 660010
rect 129810 659770 129900 660010
rect 130140 659770 130230 660010
rect 130470 659770 130580 660010
rect 130820 659770 130910 660010
rect 131150 659770 131240 660010
rect 131480 659770 131570 660010
rect 131810 659770 131920 660010
rect 132160 659770 132250 660010
rect 132490 659770 132580 660010
rect 132820 659770 132910 660010
rect 133150 659770 133570 660010
rect 133810 659770 133920 660010
rect 134160 659770 134250 660010
rect 134490 659770 134580 660010
rect 134820 659770 134910 660010
rect 135150 659770 135260 660010
rect 135500 659770 135590 660010
rect 135830 659770 135920 660010
rect 136160 659770 136250 660010
rect 136490 659770 136600 660010
rect 136840 659770 136930 660010
rect 137170 659770 137260 660010
rect 137500 659770 137590 660010
rect 137830 659770 137940 660010
rect 138180 659770 138270 660010
rect 138510 659770 138600 660010
rect 138840 659770 138930 660010
rect 139170 659770 139280 660010
rect 139520 659770 139610 660010
rect 139850 659770 139940 660010
rect 140180 659770 140270 660010
rect 140510 659770 140620 660010
rect 140860 659770 140950 660010
rect 141190 659770 141280 660010
rect 141520 659770 141610 660010
rect 141850 659770 141960 660010
rect 142200 659770 142290 660010
rect 142530 659770 142620 660010
rect 142860 659770 142950 660010
rect 143190 659770 143300 660010
rect 143540 659770 143630 660010
rect 143870 659770 143960 660010
rect 144200 659770 144290 660010
rect 144530 659770 144950 660010
rect 145190 659770 145300 660010
rect 145540 659770 145630 660010
rect 145870 659770 145960 660010
rect 146200 659770 146290 660010
rect 146530 659770 146640 660010
rect 146880 659770 146970 660010
rect 147210 659770 147300 660010
rect 147540 659770 147630 660010
rect 147870 659770 147980 660010
rect 148220 659770 148310 660010
rect 148550 659770 148640 660010
rect 148880 659770 148970 660010
rect 149210 659770 149320 660010
rect 149560 659770 149650 660010
rect 149890 659770 149980 660010
rect 150220 659770 150310 660010
rect 150550 659770 150660 660010
rect 150900 659770 150990 660010
rect 151230 659770 151320 660010
rect 151560 659770 151650 660010
rect 151890 659770 152000 660010
rect 152240 659770 152330 660010
rect 152570 659770 152660 660010
rect 152900 659770 152990 660010
rect 153230 659770 153340 660010
rect 153580 659770 153670 660010
rect 153910 659770 154000 660010
rect 154240 659770 154330 660010
rect 154570 659770 154680 660010
rect 154920 659770 155010 660010
rect 155250 659770 155340 660010
rect 155580 659770 155670 660010
rect 155910 659770 155960 660010
rect 110760 659680 155960 659770
rect 110760 659440 110810 659680
rect 111050 659440 111160 659680
rect 111400 659440 111490 659680
rect 111730 659440 111820 659680
rect 112060 659440 112150 659680
rect 112390 659440 112500 659680
rect 112740 659440 112830 659680
rect 113070 659440 113160 659680
rect 113400 659440 113490 659680
rect 113730 659440 113840 659680
rect 114080 659440 114170 659680
rect 114410 659440 114500 659680
rect 114740 659440 114830 659680
rect 115070 659440 115180 659680
rect 115420 659440 115510 659680
rect 115750 659440 115840 659680
rect 116080 659440 116170 659680
rect 116410 659440 116520 659680
rect 116760 659440 116850 659680
rect 117090 659440 117180 659680
rect 117420 659440 117510 659680
rect 117750 659440 117860 659680
rect 118100 659440 118190 659680
rect 118430 659440 118520 659680
rect 118760 659440 118850 659680
rect 119090 659440 119200 659680
rect 119440 659440 119530 659680
rect 119770 659440 119860 659680
rect 120100 659440 120190 659680
rect 120430 659440 120540 659680
rect 120780 659440 120870 659680
rect 121110 659440 121200 659680
rect 121440 659440 121530 659680
rect 121770 659440 122190 659680
rect 122430 659440 122540 659680
rect 122780 659440 122870 659680
rect 123110 659440 123200 659680
rect 123440 659440 123530 659680
rect 123770 659440 123880 659680
rect 124120 659440 124210 659680
rect 124450 659440 124540 659680
rect 124780 659440 124870 659680
rect 125110 659440 125220 659680
rect 125460 659440 125550 659680
rect 125790 659440 125880 659680
rect 126120 659440 126210 659680
rect 126450 659440 126560 659680
rect 126800 659440 126890 659680
rect 127130 659440 127220 659680
rect 127460 659440 127550 659680
rect 127790 659440 127900 659680
rect 128140 659440 128230 659680
rect 128470 659440 128560 659680
rect 128800 659440 128890 659680
rect 129130 659440 129240 659680
rect 129480 659440 129570 659680
rect 129810 659440 129900 659680
rect 130140 659440 130230 659680
rect 130470 659440 130580 659680
rect 130820 659440 130910 659680
rect 131150 659440 131240 659680
rect 131480 659440 131570 659680
rect 131810 659440 131920 659680
rect 132160 659440 132250 659680
rect 132490 659440 132580 659680
rect 132820 659440 132910 659680
rect 133150 659440 133570 659680
rect 133810 659440 133920 659680
rect 134160 659440 134250 659680
rect 134490 659440 134580 659680
rect 134820 659440 134910 659680
rect 135150 659440 135260 659680
rect 135500 659440 135590 659680
rect 135830 659440 135920 659680
rect 136160 659440 136250 659680
rect 136490 659440 136600 659680
rect 136840 659440 136930 659680
rect 137170 659440 137260 659680
rect 137500 659440 137590 659680
rect 137830 659440 137940 659680
rect 138180 659440 138270 659680
rect 138510 659440 138600 659680
rect 138840 659440 138930 659680
rect 139170 659440 139280 659680
rect 139520 659440 139610 659680
rect 139850 659440 139940 659680
rect 140180 659440 140270 659680
rect 140510 659440 140620 659680
rect 140860 659440 140950 659680
rect 141190 659440 141280 659680
rect 141520 659440 141610 659680
rect 141850 659440 141960 659680
rect 142200 659440 142290 659680
rect 142530 659440 142620 659680
rect 142860 659440 142950 659680
rect 143190 659440 143300 659680
rect 143540 659440 143630 659680
rect 143870 659440 143960 659680
rect 144200 659440 144290 659680
rect 144530 659440 144950 659680
rect 145190 659440 145300 659680
rect 145540 659440 145630 659680
rect 145870 659440 145960 659680
rect 146200 659440 146290 659680
rect 146530 659440 146640 659680
rect 146880 659440 146970 659680
rect 147210 659440 147300 659680
rect 147540 659440 147630 659680
rect 147870 659440 147980 659680
rect 148220 659440 148310 659680
rect 148550 659440 148640 659680
rect 148880 659440 148970 659680
rect 149210 659440 149320 659680
rect 149560 659440 149650 659680
rect 149890 659440 149980 659680
rect 150220 659440 150310 659680
rect 150550 659440 150660 659680
rect 150900 659440 150990 659680
rect 151230 659440 151320 659680
rect 151560 659440 151650 659680
rect 151890 659440 152000 659680
rect 152240 659440 152330 659680
rect 152570 659440 152660 659680
rect 152900 659440 152990 659680
rect 153230 659440 153340 659680
rect 153580 659440 153670 659680
rect 153910 659440 154000 659680
rect 154240 659440 154330 659680
rect 154570 659440 154680 659680
rect 154920 659440 155010 659680
rect 155250 659440 155340 659680
rect 155580 659440 155670 659680
rect 155910 659440 155960 659680
rect 110760 659350 155960 659440
rect 110760 659110 110810 659350
rect 111050 659110 111160 659350
rect 111400 659110 111490 659350
rect 111730 659110 111820 659350
rect 112060 659110 112150 659350
rect 112390 659110 112500 659350
rect 112740 659110 112830 659350
rect 113070 659110 113160 659350
rect 113400 659110 113490 659350
rect 113730 659110 113840 659350
rect 114080 659110 114170 659350
rect 114410 659110 114500 659350
rect 114740 659110 114830 659350
rect 115070 659110 115180 659350
rect 115420 659110 115510 659350
rect 115750 659110 115840 659350
rect 116080 659110 116170 659350
rect 116410 659110 116520 659350
rect 116760 659110 116850 659350
rect 117090 659110 117180 659350
rect 117420 659110 117510 659350
rect 117750 659110 117860 659350
rect 118100 659110 118190 659350
rect 118430 659110 118520 659350
rect 118760 659110 118850 659350
rect 119090 659110 119200 659350
rect 119440 659110 119530 659350
rect 119770 659110 119860 659350
rect 120100 659110 120190 659350
rect 120430 659110 120540 659350
rect 120780 659110 120870 659350
rect 121110 659110 121200 659350
rect 121440 659110 121530 659350
rect 121770 659110 122190 659350
rect 122430 659110 122540 659350
rect 122780 659110 122870 659350
rect 123110 659110 123200 659350
rect 123440 659110 123530 659350
rect 123770 659110 123880 659350
rect 124120 659110 124210 659350
rect 124450 659110 124540 659350
rect 124780 659110 124870 659350
rect 125110 659110 125220 659350
rect 125460 659110 125550 659350
rect 125790 659110 125880 659350
rect 126120 659110 126210 659350
rect 126450 659110 126560 659350
rect 126800 659110 126890 659350
rect 127130 659110 127220 659350
rect 127460 659110 127550 659350
rect 127790 659110 127900 659350
rect 128140 659110 128230 659350
rect 128470 659110 128560 659350
rect 128800 659110 128890 659350
rect 129130 659110 129240 659350
rect 129480 659110 129570 659350
rect 129810 659110 129900 659350
rect 130140 659110 130230 659350
rect 130470 659110 130580 659350
rect 130820 659110 130910 659350
rect 131150 659110 131240 659350
rect 131480 659110 131570 659350
rect 131810 659110 131920 659350
rect 132160 659110 132250 659350
rect 132490 659110 132580 659350
rect 132820 659110 132910 659350
rect 133150 659110 133570 659350
rect 133810 659110 133920 659350
rect 134160 659110 134250 659350
rect 134490 659110 134580 659350
rect 134820 659110 134910 659350
rect 135150 659110 135260 659350
rect 135500 659110 135590 659350
rect 135830 659110 135920 659350
rect 136160 659110 136250 659350
rect 136490 659110 136600 659350
rect 136840 659110 136930 659350
rect 137170 659110 137260 659350
rect 137500 659110 137590 659350
rect 137830 659110 137940 659350
rect 138180 659110 138270 659350
rect 138510 659110 138600 659350
rect 138840 659110 138930 659350
rect 139170 659110 139280 659350
rect 139520 659110 139610 659350
rect 139850 659110 139940 659350
rect 140180 659110 140270 659350
rect 140510 659110 140620 659350
rect 140860 659110 140950 659350
rect 141190 659110 141280 659350
rect 141520 659110 141610 659350
rect 141850 659110 141960 659350
rect 142200 659110 142290 659350
rect 142530 659110 142620 659350
rect 142860 659110 142950 659350
rect 143190 659110 143300 659350
rect 143540 659110 143630 659350
rect 143870 659110 143960 659350
rect 144200 659110 144290 659350
rect 144530 659110 144950 659350
rect 145190 659110 145300 659350
rect 145540 659110 145630 659350
rect 145870 659110 145960 659350
rect 146200 659110 146290 659350
rect 146530 659110 146640 659350
rect 146880 659110 146970 659350
rect 147210 659110 147300 659350
rect 147540 659110 147630 659350
rect 147870 659110 147980 659350
rect 148220 659110 148310 659350
rect 148550 659110 148640 659350
rect 148880 659110 148970 659350
rect 149210 659110 149320 659350
rect 149560 659110 149650 659350
rect 149890 659110 149980 659350
rect 150220 659110 150310 659350
rect 150550 659110 150660 659350
rect 150900 659110 150990 659350
rect 151230 659110 151320 659350
rect 151560 659110 151650 659350
rect 151890 659110 152000 659350
rect 152240 659110 152330 659350
rect 152570 659110 152660 659350
rect 152900 659110 152990 659350
rect 153230 659110 153340 659350
rect 153580 659110 153670 659350
rect 153910 659110 154000 659350
rect 154240 659110 154330 659350
rect 154570 659110 154680 659350
rect 154920 659110 155010 659350
rect 155250 659110 155340 659350
rect 155580 659110 155670 659350
rect 155910 659110 155960 659350
rect 110760 659000 155960 659110
rect 110760 658760 110810 659000
rect 111050 658760 111160 659000
rect 111400 658760 111490 659000
rect 111730 658760 111820 659000
rect 112060 658760 112150 659000
rect 112390 658760 112500 659000
rect 112740 658760 112830 659000
rect 113070 658760 113160 659000
rect 113400 658760 113490 659000
rect 113730 658760 113840 659000
rect 114080 658760 114170 659000
rect 114410 658760 114500 659000
rect 114740 658760 114830 659000
rect 115070 658760 115180 659000
rect 115420 658760 115510 659000
rect 115750 658760 115840 659000
rect 116080 658760 116170 659000
rect 116410 658760 116520 659000
rect 116760 658760 116850 659000
rect 117090 658760 117180 659000
rect 117420 658760 117510 659000
rect 117750 658760 117860 659000
rect 118100 658760 118190 659000
rect 118430 658760 118520 659000
rect 118760 658760 118850 659000
rect 119090 658760 119200 659000
rect 119440 658760 119530 659000
rect 119770 658760 119860 659000
rect 120100 658760 120190 659000
rect 120430 658760 120540 659000
rect 120780 658760 120870 659000
rect 121110 658760 121200 659000
rect 121440 658760 121530 659000
rect 121770 658760 122190 659000
rect 122430 658760 122540 659000
rect 122780 658760 122870 659000
rect 123110 658760 123200 659000
rect 123440 658760 123530 659000
rect 123770 658760 123880 659000
rect 124120 658760 124210 659000
rect 124450 658760 124540 659000
rect 124780 658760 124870 659000
rect 125110 658760 125220 659000
rect 125460 658760 125550 659000
rect 125790 658760 125880 659000
rect 126120 658760 126210 659000
rect 126450 658760 126560 659000
rect 126800 658760 126890 659000
rect 127130 658760 127220 659000
rect 127460 658760 127550 659000
rect 127790 658760 127900 659000
rect 128140 658760 128230 659000
rect 128470 658760 128560 659000
rect 128800 658760 128890 659000
rect 129130 658760 129240 659000
rect 129480 658760 129570 659000
rect 129810 658760 129900 659000
rect 130140 658760 130230 659000
rect 130470 658760 130580 659000
rect 130820 658760 130910 659000
rect 131150 658760 131240 659000
rect 131480 658760 131570 659000
rect 131810 658760 131920 659000
rect 132160 658760 132250 659000
rect 132490 658760 132580 659000
rect 132820 658760 132910 659000
rect 133150 658760 133570 659000
rect 133810 658760 133920 659000
rect 134160 658760 134250 659000
rect 134490 658760 134580 659000
rect 134820 658760 134910 659000
rect 135150 658760 135260 659000
rect 135500 658760 135590 659000
rect 135830 658760 135920 659000
rect 136160 658760 136250 659000
rect 136490 658760 136600 659000
rect 136840 658760 136930 659000
rect 137170 658760 137260 659000
rect 137500 658760 137590 659000
rect 137830 658760 137940 659000
rect 138180 658760 138270 659000
rect 138510 658760 138600 659000
rect 138840 658760 138930 659000
rect 139170 658760 139280 659000
rect 139520 658760 139610 659000
rect 139850 658760 139940 659000
rect 140180 658760 140270 659000
rect 140510 658760 140620 659000
rect 140860 658760 140950 659000
rect 141190 658760 141280 659000
rect 141520 658760 141610 659000
rect 141850 658760 141960 659000
rect 142200 658760 142290 659000
rect 142530 658760 142620 659000
rect 142860 658760 142950 659000
rect 143190 658760 143300 659000
rect 143540 658760 143630 659000
rect 143870 658760 143960 659000
rect 144200 658760 144290 659000
rect 144530 658760 144950 659000
rect 145190 658760 145300 659000
rect 145540 658760 145630 659000
rect 145870 658760 145960 659000
rect 146200 658760 146290 659000
rect 146530 658760 146640 659000
rect 146880 658760 146970 659000
rect 147210 658760 147300 659000
rect 147540 658760 147630 659000
rect 147870 658760 147980 659000
rect 148220 658760 148310 659000
rect 148550 658760 148640 659000
rect 148880 658760 148970 659000
rect 149210 658760 149320 659000
rect 149560 658760 149650 659000
rect 149890 658760 149980 659000
rect 150220 658760 150310 659000
rect 150550 658760 150660 659000
rect 150900 658760 150990 659000
rect 151230 658760 151320 659000
rect 151560 658760 151650 659000
rect 151890 658760 152000 659000
rect 152240 658760 152330 659000
rect 152570 658760 152660 659000
rect 152900 658760 152990 659000
rect 153230 658760 153340 659000
rect 153580 658760 153670 659000
rect 153910 658760 154000 659000
rect 154240 658760 154330 659000
rect 154570 658760 154680 659000
rect 154920 658760 155010 659000
rect 155250 658760 155340 659000
rect 155580 658760 155670 659000
rect 155910 658760 155960 659000
rect 110760 658670 155960 658760
rect 110760 658430 110810 658670
rect 111050 658430 111160 658670
rect 111400 658430 111490 658670
rect 111730 658430 111820 658670
rect 112060 658430 112150 658670
rect 112390 658430 112500 658670
rect 112740 658430 112830 658670
rect 113070 658430 113160 658670
rect 113400 658430 113490 658670
rect 113730 658430 113840 658670
rect 114080 658430 114170 658670
rect 114410 658430 114500 658670
rect 114740 658430 114830 658670
rect 115070 658430 115180 658670
rect 115420 658430 115510 658670
rect 115750 658430 115840 658670
rect 116080 658430 116170 658670
rect 116410 658430 116520 658670
rect 116760 658430 116850 658670
rect 117090 658430 117180 658670
rect 117420 658430 117510 658670
rect 117750 658430 117860 658670
rect 118100 658430 118190 658670
rect 118430 658430 118520 658670
rect 118760 658430 118850 658670
rect 119090 658430 119200 658670
rect 119440 658430 119530 658670
rect 119770 658430 119860 658670
rect 120100 658430 120190 658670
rect 120430 658430 120540 658670
rect 120780 658430 120870 658670
rect 121110 658430 121200 658670
rect 121440 658430 121530 658670
rect 121770 658430 122190 658670
rect 122430 658430 122540 658670
rect 122780 658430 122870 658670
rect 123110 658430 123200 658670
rect 123440 658430 123530 658670
rect 123770 658430 123880 658670
rect 124120 658430 124210 658670
rect 124450 658430 124540 658670
rect 124780 658430 124870 658670
rect 125110 658430 125220 658670
rect 125460 658430 125550 658670
rect 125790 658430 125880 658670
rect 126120 658430 126210 658670
rect 126450 658430 126560 658670
rect 126800 658430 126890 658670
rect 127130 658430 127220 658670
rect 127460 658430 127550 658670
rect 127790 658430 127900 658670
rect 128140 658430 128230 658670
rect 128470 658430 128560 658670
rect 128800 658430 128890 658670
rect 129130 658430 129240 658670
rect 129480 658430 129570 658670
rect 129810 658430 129900 658670
rect 130140 658430 130230 658670
rect 130470 658430 130580 658670
rect 130820 658430 130910 658670
rect 131150 658430 131240 658670
rect 131480 658430 131570 658670
rect 131810 658430 131920 658670
rect 132160 658430 132250 658670
rect 132490 658430 132580 658670
rect 132820 658430 132910 658670
rect 133150 658430 133570 658670
rect 133810 658430 133920 658670
rect 134160 658430 134250 658670
rect 134490 658430 134580 658670
rect 134820 658430 134910 658670
rect 135150 658430 135260 658670
rect 135500 658430 135590 658670
rect 135830 658430 135920 658670
rect 136160 658430 136250 658670
rect 136490 658430 136600 658670
rect 136840 658430 136930 658670
rect 137170 658430 137260 658670
rect 137500 658430 137590 658670
rect 137830 658430 137940 658670
rect 138180 658430 138270 658670
rect 138510 658430 138600 658670
rect 138840 658430 138930 658670
rect 139170 658430 139280 658670
rect 139520 658430 139610 658670
rect 139850 658430 139940 658670
rect 140180 658430 140270 658670
rect 140510 658430 140620 658670
rect 140860 658430 140950 658670
rect 141190 658430 141280 658670
rect 141520 658430 141610 658670
rect 141850 658430 141960 658670
rect 142200 658430 142290 658670
rect 142530 658430 142620 658670
rect 142860 658430 142950 658670
rect 143190 658430 143300 658670
rect 143540 658430 143630 658670
rect 143870 658430 143960 658670
rect 144200 658430 144290 658670
rect 144530 658430 144950 658670
rect 145190 658430 145300 658670
rect 145540 658430 145630 658670
rect 145870 658430 145960 658670
rect 146200 658430 146290 658670
rect 146530 658430 146640 658670
rect 146880 658430 146970 658670
rect 147210 658430 147300 658670
rect 147540 658430 147630 658670
rect 147870 658430 147980 658670
rect 148220 658430 148310 658670
rect 148550 658430 148640 658670
rect 148880 658430 148970 658670
rect 149210 658430 149320 658670
rect 149560 658430 149650 658670
rect 149890 658430 149980 658670
rect 150220 658430 150310 658670
rect 150550 658430 150660 658670
rect 150900 658430 150990 658670
rect 151230 658430 151320 658670
rect 151560 658430 151650 658670
rect 151890 658430 152000 658670
rect 152240 658430 152330 658670
rect 152570 658430 152660 658670
rect 152900 658430 152990 658670
rect 153230 658430 153340 658670
rect 153580 658430 153670 658670
rect 153910 658430 154000 658670
rect 154240 658430 154330 658670
rect 154570 658430 154680 658670
rect 154920 658430 155010 658670
rect 155250 658430 155340 658670
rect 155580 658430 155670 658670
rect 155910 658430 155960 658670
rect 110760 658340 155960 658430
rect 110760 658100 110810 658340
rect 111050 658100 111160 658340
rect 111400 658100 111490 658340
rect 111730 658100 111820 658340
rect 112060 658100 112150 658340
rect 112390 658100 112500 658340
rect 112740 658100 112830 658340
rect 113070 658100 113160 658340
rect 113400 658100 113490 658340
rect 113730 658100 113840 658340
rect 114080 658100 114170 658340
rect 114410 658100 114500 658340
rect 114740 658100 114830 658340
rect 115070 658100 115180 658340
rect 115420 658100 115510 658340
rect 115750 658100 115840 658340
rect 116080 658100 116170 658340
rect 116410 658100 116520 658340
rect 116760 658100 116850 658340
rect 117090 658100 117180 658340
rect 117420 658100 117510 658340
rect 117750 658100 117860 658340
rect 118100 658100 118190 658340
rect 118430 658100 118520 658340
rect 118760 658100 118850 658340
rect 119090 658100 119200 658340
rect 119440 658100 119530 658340
rect 119770 658100 119860 658340
rect 120100 658100 120190 658340
rect 120430 658100 120540 658340
rect 120780 658100 120870 658340
rect 121110 658100 121200 658340
rect 121440 658100 121530 658340
rect 121770 658100 122190 658340
rect 122430 658100 122540 658340
rect 122780 658100 122870 658340
rect 123110 658100 123200 658340
rect 123440 658100 123530 658340
rect 123770 658100 123880 658340
rect 124120 658100 124210 658340
rect 124450 658100 124540 658340
rect 124780 658100 124870 658340
rect 125110 658100 125220 658340
rect 125460 658100 125550 658340
rect 125790 658100 125880 658340
rect 126120 658100 126210 658340
rect 126450 658100 126560 658340
rect 126800 658100 126890 658340
rect 127130 658100 127220 658340
rect 127460 658100 127550 658340
rect 127790 658100 127900 658340
rect 128140 658100 128230 658340
rect 128470 658100 128560 658340
rect 128800 658100 128890 658340
rect 129130 658100 129240 658340
rect 129480 658100 129570 658340
rect 129810 658100 129900 658340
rect 130140 658100 130230 658340
rect 130470 658100 130580 658340
rect 130820 658100 130910 658340
rect 131150 658100 131240 658340
rect 131480 658100 131570 658340
rect 131810 658100 131920 658340
rect 132160 658100 132250 658340
rect 132490 658100 132580 658340
rect 132820 658100 132910 658340
rect 133150 658100 133570 658340
rect 133810 658100 133920 658340
rect 134160 658100 134250 658340
rect 134490 658100 134580 658340
rect 134820 658100 134910 658340
rect 135150 658100 135260 658340
rect 135500 658100 135590 658340
rect 135830 658100 135920 658340
rect 136160 658100 136250 658340
rect 136490 658100 136600 658340
rect 136840 658100 136930 658340
rect 137170 658100 137260 658340
rect 137500 658100 137590 658340
rect 137830 658100 137940 658340
rect 138180 658100 138270 658340
rect 138510 658100 138600 658340
rect 138840 658100 138930 658340
rect 139170 658100 139280 658340
rect 139520 658100 139610 658340
rect 139850 658100 139940 658340
rect 140180 658100 140270 658340
rect 140510 658100 140620 658340
rect 140860 658100 140950 658340
rect 141190 658100 141280 658340
rect 141520 658100 141610 658340
rect 141850 658100 141960 658340
rect 142200 658100 142290 658340
rect 142530 658100 142620 658340
rect 142860 658100 142950 658340
rect 143190 658100 143300 658340
rect 143540 658100 143630 658340
rect 143870 658100 143960 658340
rect 144200 658100 144290 658340
rect 144530 658100 144950 658340
rect 145190 658100 145300 658340
rect 145540 658100 145630 658340
rect 145870 658100 145960 658340
rect 146200 658100 146290 658340
rect 146530 658100 146640 658340
rect 146880 658100 146970 658340
rect 147210 658100 147300 658340
rect 147540 658100 147630 658340
rect 147870 658100 147980 658340
rect 148220 658100 148310 658340
rect 148550 658100 148640 658340
rect 148880 658100 148970 658340
rect 149210 658100 149320 658340
rect 149560 658100 149650 658340
rect 149890 658100 149980 658340
rect 150220 658100 150310 658340
rect 150550 658100 150660 658340
rect 150900 658100 150990 658340
rect 151230 658100 151320 658340
rect 151560 658100 151650 658340
rect 151890 658100 152000 658340
rect 152240 658100 152330 658340
rect 152570 658100 152660 658340
rect 152900 658100 152990 658340
rect 153230 658100 153340 658340
rect 153580 658100 153670 658340
rect 153910 658100 154000 658340
rect 154240 658100 154330 658340
rect 154570 658100 154680 658340
rect 154920 658100 155010 658340
rect 155250 658100 155340 658340
rect 155580 658100 155670 658340
rect 155910 658100 155960 658340
rect 110760 658010 155960 658100
rect 110760 657770 110810 658010
rect 111050 657770 111160 658010
rect 111400 657770 111490 658010
rect 111730 657770 111820 658010
rect 112060 657770 112150 658010
rect 112390 657770 112500 658010
rect 112740 657770 112830 658010
rect 113070 657770 113160 658010
rect 113400 657770 113490 658010
rect 113730 657770 113840 658010
rect 114080 657770 114170 658010
rect 114410 657770 114500 658010
rect 114740 657770 114830 658010
rect 115070 657770 115180 658010
rect 115420 657770 115510 658010
rect 115750 657770 115840 658010
rect 116080 657770 116170 658010
rect 116410 657770 116520 658010
rect 116760 657770 116850 658010
rect 117090 657770 117180 658010
rect 117420 657770 117510 658010
rect 117750 657770 117860 658010
rect 118100 657770 118190 658010
rect 118430 657770 118520 658010
rect 118760 657770 118850 658010
rect 119090 657770 119200 658010
rect 119440 657770 119530 658010
rect 119770 657770 119860 658010
rect 120100 657770 120190 658010
rect 120430 657770 120540 658010
rect 120780 657770 120870 658010
rect 121110 657770 121200 658010
rect 121440 657770 121530 658010
rect 121770 657770 122190 658010
rect 122430 657770 122540 658010
rect 122780 657770 122870 658010
rect 123110 657770 123200 658010
rect 123440 657770 123530 658010
rect 123770 657770 123880 658010
rect 124120 657770 124210 658010
rect 124450 657770 124540 658010
rect 124780 657770 124870 658010
rect 125110 657770 125220 658010
rect 125460 657770 125550 658010
rect 125790 657770 125880 658010
rect 126120 657770 126210 658010
rect 126450 657770 126560 658010
rect 126800 657770 126890 658010
rect 127130 657770 127220 658010
rect 127460 657770 127550 658010
rect 127790 657770 127900 658010
rect 128140 657770 128230 658010
rect 128470 657770 128560 658010
rect 128800 657770 128890 658010
rect 129130 657770 129240 658010
rect 129480 657770 129570 658010
rect 129810 657770 129900 658010
rect 130140 657770 130230 658010
rect 130470 657770 130580 658010
rect 130820 657770 130910 658010
rect 131150 657770 131240 658010
rect 131480 657770 131570 658010
rect 131810 657770 131920 658010
rect 132160 657770 132250 658010
rect 132490 657770 132580 658010
rect 132820 657770 132910 658010
rect 133150 657770 133570 658010
rect 133810 657770 133920 658010
rect 134160 657770 134250 658010
rect 134490 657770 134580 658010
rect 134820 657770 134910 658010
rect 135150 657770 135260 658010
rect 135500 657770 135590 658010
rect 135830 657770 135920 658010
rect 136160 657770 136250 658010
rect 136490 657770 136600 658010
rect 136840 657770 136930 658010
rect 137170 657770 137260 658010
rect 137500 657770 137590 658010
rect 137830 657770 137940 658010
rect 138180 657770 138270 658010
rect 138510 657770 138600 658010
rect 138840 657770 138930 658010
rect 139170 657770 139280 658010
rect 139520 657770 139610 658010
rect 139850 657770 139940 658010
rect 140180 657770 140270 658010
rect 140510 657770 140620 658010
rect 140860 657770 140950 658010
rect 141190 657770 141280 658010
rect 141520 657770 141610 658010
rect 141850 657770 141960 658010
rect 142200 657770 142290 658010
rect 142530 657770 142620 658010
rect 142860 657770 142950 658010
rect 143190 657770 143300 658010
rect 143540 657770 143630 658010
rect 143870 657770 143960 658010
rect 144200 657770 144290 658010
rect 144530 657770 144950 658010
rect 145190 657770 145300 658010
rect 145540 657770 145630 658010
rect 145870 657770 145960 658010
rect 146200 657770 146290 658010
rect 146530 657770 146640 658010
rect 146880 657770 146970 658010
rect 147210 657770 147300 658010
rect 147540 657770 147630 658010
rect 147870 657770 147980 658010
rect 148220 657770 148310 658010
rect 148550 657770 148640 658010
rect 148880 657770 148970 658010
rect 149210 657770 149320 658010
rect 149560 657770 149650 658010
rect 149890 657770 149980 658010
rect 150220 657770 150310 658010
rect 150550 657770 150660 658010
rect 150900 657770 150990 658010
rect 151230 657770 151320 658010
rect 151560 657770 151650 658010
rect 151890 657770 152000 658010
rect 152240 657770 152330 658010
rect 152570 657770 152660 658010
rect 152900 657770 152990 658010
rect 153230 657770 153340 658010
rect 153580 657770 153670 658010
rect 153910 657770 154000 658010
rect 154240 657770 154330 658010
rect 154570 657770 154680 658010
rect 154920 657770 155010 658010
rect 155250 657770 155340 658010
rect 155580 657770 155670 658010
rect 155910 657770 155960 658010
rect 110760 657660 155960 657770
rect 110760 657420 110810 657660
rect 111050 657420 111160 657660
rect 111400 657420 111490 657660
rect 111730 657420 111820 657660
rect 112060 657420 112150 657660
rect 112390 657420 112500 657660
rect 112740 657420 112830 657660
rect 113070 657420 113160 657660
rect 113400 657420 113490 657660
rect 113730 657420 113840 657660
rect 114080 657420 114170 657660
rect 114410 657420 114500 657660
rect 114740 657420 114830 657660
rect 115070 657420 115180 657660
rect 115420 657420 115510 657660
rect 115750 657420 115840 657660
rect 116080 657420 116170 657660
rect 116410 657420 116520 657660
rect 116760 657420 116850 657660
rect 117090 657420 117180 657660
rect 117420 657420 117510 657660
rect 117750 657420 117860 657660
rect 118100 657420 118190 657660
rect 118430 657420 118520 657660
rect 118760 657420 118850 657660
rect 119090 657420 119200 657660
rect 119440 657420 119530 657660
rect 119770 657420 119860 657660
rect 120100 657420 120190 657660
rect 120430 657420 120540 657660
rect 120780 657420 120870 657660
rect 121110 657420 121200 657660
rect 121440 657420 121530 657660
rect 121770 657420 122190 657660
rect 122430 657420 122540 657660
rect 122780 657420 122870 657660
rect 123110 657420 123200 657660
rect 123440 657420 123530 657660
rect 123770 657420 123880 657660
rect 124120 657420 124210 657660
rect 124450 657420 124540 657660
rect 124780 657420 124870 657660
rect 125110 657420 125220 657660
rect 125460 657420 125550 657660
rect 125790 657420 125880 657660
rect 126120 657420 126210 657660
rect 126450 657420 126560 657660
rect 126800 657420 126890 657660
rect 127130 657420 127220 657660
rect 127460 657420 127550 657660
rect 127790 657420 127900 657660
rect 128140 657420 128230 657660
rect 128470 657420 128560 657660
rect 128800 657420 128890 657660
rect 129130 657420 129240 657660
rect 129480 657420 129570 657660
rect 129810 657420 129900 657660
rect 130140 657420 130230 657660
rect 130470 657420 130580 657660
rect 130820 657420 130910 657660
rect 131150 657420 131240 657660
rect 131480 657420 131570 657660
rect 131810 657420 131920 657660
rect 132160 657420 132250 657660
rect 132490 657420 132580 657660
rect 132820 657420 132910 657660
rect 133150 657420 133570 657660
rect 133810 657420 133920 657660
rect 134160 657420 134250 657660
rect 134490 657420 134580 657660
rect 134820 657420 134910 657660
rect 135150 657420 135260 657660
rect 135500 657420 135590 657660
rect 135830 657420 135920 657660
rect 136160 657420 136250 657660
rect 136490 657420 136600 657660
rect 136840 657420 136930 657660
rect 137170 657420 137260 657660
rect 137500 657420 137590 657660
rect 137830 657420 137940 657660
rect 138180 657420 138270 657660
rect 138510 657420 138600 657660
rect 138840 657420 138930 657660
rect 139170 657420 139280 657660
rect 139520 657420 139610 657660
rect 139850 657420 139940 657660
rect 140180 657420 140270 657660
rect 140510 657420 140620 657660
rect 140860 657420 140950 657660
rect 141190 657420 141280 657660
rect 141520 657420 141610 657660
rect 141850 657420 141960 657660
rect 142200 657420 142290 657660
rect 142530 657420 142620 657660
rect 142860 657420 142950 657660
rect 143190 657420 143300 657660
rect 143540 657420 143630 657660
rect 143870 657420 143960 657660
rect 144200 657420 144290 657660
rect 144530 657420 144950 657660
rect 145190 657420 145300 657660
rect 145540 657420 145630 657660
rect 145870 657420 145960 657660
rect 146200 657420 146290 657660
rect 146530 657420 146640 657660
rect 146880 657420 146970 657660
rect 147210 657420 147300 657660
rect 147540 657420 147630 657660
rect 147870 657420 147980 657660
rect 148220 657420 148310 657660
rect 148550 657420 148640 657660
rect 148880 657420 148970 657660
rect 149210 657420 149320 657660
rect 149560 657420 149650 657660
rect 149890 657420 149980 657660
rect 150220 657420 150310 657660
rect 150550 657420 150660 657660
rect 150900 657420 150990 657660
rect 151230 657420 151320 657660
rect 151560 657420 151650 657660
rect 151890 657420 152000 657660
rect 152240 657420 152330 657660
rect 152570 657420 152660 657660
rect 152900 657420 152990 657660
rect 153230 657420 153340 657660
rect 153580 657420 153670 657660
rect 153910 657420 154000 657660
rect 154240 657420 154330 657660
rect 154570 657420 154680 657660
rect 154920 657420 155010 657660
rect 155250 657420 155340 657660
rect 155580 657420 155670 657660
rect 155910 657420 155960 657660
rect 110760 657330 155960 657420
rect 110760 657090 110810 657330
rect 111050 657090 111160 657330
rect 111400 657090 111490 657330
rect 111730 657090 111820 657330
rect 112060 657090 112150 657330
rect 112390 657090 112500 657330
rect 112740 657090 112830 657330
rect 113070 657090 113160 657330
rect 113400 657090 113490 657330
rect 113730 657090 113840 657330
rect 114080 657090 114170 657330
rect 114410 657090 114500 657330
rect 114740 657090 114830 657330
rect 115070 657090 115180 657330
rect 115420 657090 115510 657330
rect 115750 657090 115840 657330
rect 116080 657090 116170 657330
rect 116410 657090 116520 657330
rect 116760 657090 116850 657330
rect 117090 657090 117180 657330
rect 117420 657090 117510 657330
rect 117750 657090 117860 657330
rect 118100 657090 118190 657330
rect 118430 657090 118520 657330
rect 118760 657090 118850 657330
rect 119090 657090 119200 657330
rect 119440 657090 119530 657330
rect 119770 657090 119860 657330
rect 120100 657090 120190 657330
rect 120430 657090 120540 657330
rect 120780 657090 120870 657330
rect 121110 657090 121200 657330
rect 121440 657090 121530 657330
rect 121770 657090 122190 657330
rect 122430 657090 122540 657330
rect 122780 657090 122870 657330
rect 123110 657090 123200 657330
rect 123440 657090 123530 657330
rect 123770 657090 123880 657330
rect 124120 657090 124210 657330
rect 124450 657090 124540 657330
rect 124780 657090 124870 657330
rect 125110 657090 125220 657330
rect 125460 657090 125550 657330
rect 125790 657090 125880 657330
rect 126120 657090 126210 657330
rect 126450 657090 126560 657330
rect 126800 657090 126890 657330
rect 127130 657090 127220 657330
rect 127460 657090 127550 657330
rect 127790 657090 127900 657330
rect 128140 657090 128230 657330
rect 128470 657090 128560 657330
rect 128800 657090 128890 657330
rect 129130 657090 129240 657330
rect 129480 657090 129570 657330
rect 129810 657090 129900 657330
rect 130140 657090 130230 657330
rect 130470 657090 130580 657330
rect 130820 657090 130910 657330
rect 131150 657090 131240 657330
rect 131480 657090 131570 657330
rect 131810 657090 131920 657330
rect 132160 657090 132250 657330
rect 132490 657090 132580 657330
rect 132820 657090 132910 657330
rect 133150 657090 133570 657330
rect 133810 657090 133920 657330
rect 134160 657090 134250 657330
rect 134490 657090 134580 657330
rect 134820 657090 134910 657330
rect 135150 657090 135260 657330
rect 135500 657090 135590 657330
rect 135830 657090 135920 657330
rect 136160 657090 136250 657330
rect 136490 657090 136600 657330
rect 136840 657090 136930 657330
rect 137170 657090 137260 657330
rect 137500 657090 137590 657330
rect 137830 657090 137940 657330
rect 138180 657090 138270 657330
rect 138510 657090 138600 657330
rect 138840 657090 138930 657330
rect 139170 657090 139280 657330
rect 139520 657090 139610 657330
rect 139850 657090 139940 657330
rect 140180 657090 140270 657330
rect 140510 657090 140620 657330
rect 140860 657090 140950 657330
rect 141190 657090 141280 657330
rect 141520 657090 141610 657330
rect 141850 657090 141960 657330
rect 142200 657090 142290 657330
rect 142530 657090 142620 657330
rect 142860 657090 142950 657330
rect 143190 657090 143300 657330
rect 143540 657090 143630 657330
rect 143870 657090 143960 657330
rect 144200 657090 144290 657330
rect 144530 657090 144950 657330
rect 145190 657090 145300 657330
rect 145540 657090 145630 657330
rect 145870 657090 145960 657330
rect 146200 657090 146290 657330
rect 146530 657090 146640 657330
rect 146880 657090 146970 657330
rect 147210 657090 147300 657330
rect 147540 657090 147630 657330
rect 147870 657090 147980 657330
rect 148220 657090 148310 657330
rect 148550 657090 148640 657330
rect 148880 657090 148970 657330
rect 149210 657090 149320 657330
rect 149560 657090 149650 657330
rect 149890 657090 149980 657330
rect 150220 657090 150310 657330
rect 150550 657090 150660 657330
rect 150900 657090 150990 657330
rect 151230 657090 151320 657330
rect 151560 657090 151650 657330
rect 151890 657090 152000 657330
rect 152240 657090 152330 657330
rect 152570 657090 152660 657330
rect 152900 657090 152990 657330
rect 153230 657090 153340 657330
rect 153580 657090 153670 657330
rect 153910 657090 154000 657330
rect 154240 657090 154330 657330
rect 154570 657090 154680 657330
rect 154920 657090 155010 657330
rect 155250 657090 155340 657330
rect 155580 657090 155670 657330
rect 155910 657090 155960 657330
rect 110760 657000 155960 657090
rect 110760 656760 110810 657000
rect 111050 656760 111160 657000
rect 111400 656760 111490 657000
rect 111730 656760 111820 657000
rect 112060 656760 112150 657000
rect 112390 656760 112500 657000
rect 112740 656760 112830 657000
rect 113070 656760 113160 657000
rect 113400 656760 113490 657000
rect 113730 656760 113840 657000
rect 114080 656760 114170 657000
rect 114410 656760 114500 657000
rect 114740 656760 114830 657000
rect 115070 656760 115180 657000
rect 115420 656760 115510 657000
rect 115750 656760 115840 657000
rect 116080 656760 116170 657000
rect 116410 656760 116520 657000
rect 116760 656760 116850 657000
rect 117090 656760 117180 657000
rect 117420 656760 117510 657000
rect 117750 656760 117860 657000
rect 118100 656760 118190 657000
rect 118430 656760 118520 657000
rect 118760 656760 118850 657000
rect 119090 656760 119200 657000
rect 119440 656760 119530 657000
rect 119770 656760 119860 657000
rect 120100 656760 120190 657000
rect 120430 656760 120540 657000
rect 120780 656760 120870 657000
rect 121110 656760 121200 657000
rect 121440 656760 121530 657000
rect 121770 656760 122190 657000
rect 122430 656760 122540 657000
rect 122780 656760 122870 657000
rect 123110 656760 123200 657000
rect 123440 656760 123530 657000
rect 123770 656760 123880 657000
rect 124120 656760 124210 657000
rect 124450 656760 124540 657000
rect 124780 656760 124870 657000
rect 125110 656760 125220 657000
rect 125460 656760 125550 657000
rect 125790 656760 125880 657000
rect 126120 656760 126210 657000
rect 126450 656760 126560 657000
rect 126800 656760 126890 657000
rect 127130 656760 127220 657000
rect 127460 656760 127550 657000
rect 127790 656760 127900 657000
rect 128140 656760 128230 657000
rect 128470 656760 128560 657000
rect 128800 656760 128890 657000
rect 129130 656760 129240 657000
rect 129480 656760 129570 657000
rect 129810 656760 129900 657000
rect 130140 656760 130230 657000
rect 130470 656760 130580 657000
rect 130820 656760 130910 657000
rect 131150 656760 131240 657000
rect 131480 656760 131570 657000
rect 131810 656760 131920 657000
rect 132160 656760 132250 657000
rect 132490 656760 132580 657000
rect 132820 656760 132910 657000
rect 133150 656760 133570 657000
rect 133810 656760 133920 657000
rect 134160 656760 134250 657000
rect 134490 656760 134580 657000
rect 134820 656760 134910 657000
rect 135150 656760 135260 657000
rect 135500 656760 135590 657000
rect 135830 656760 135920 657000
rect 136160 656760 136250 657000
rect 136490 656760 136600 657000
rect 136840 656760 136930 657000
rect 137170 656760 137260 657000
rect 137500 656760 137590 657000
rect 137830 656760 137940 657000
rect 138180 656760 138270 657000
rect 138510 656760 138600 657000
rect 138840 656760 138930 657000
rect 139170 656760 139280 657000
rect 139520 656760 139610 657000
rect 139850 656760 139940 657000
rect 140180 656760 140270 657000
rect 140510 656760 140620 657000
rect 140860 656760 140950 657000
rect 141190 656760 141280 657000
rect 141520 656760 141610 657000
rect 141850 656760 141960 657000
rect 142200 656760 142290 657000
rect 142530 656760 142620 657000
rect 142860 656760 142950 657000
rect 143190 656760 143300 657000
rect 143540 656760 143630 657000
rect 143870 656760 143960 657000
rect 144200 656760 144290 657000
rect 144530 656760 144950 657000
rect 145190 656760 145300 657000
rect 145540 656760 145630 657000
rect 145870 656760 145960 657000
rect 146200 656760 146290 657000
rect 146530 656760 146640 657000
rect 146880 656760 146970 657000
rect 147210 656760 147300 657000
rect 147540 656760 147630 657000
rect 147870 656760 147980 657000
rect 148220 656760 148310 657000
rect 148550 656760 148640 657000
rect 148880 656760 148970 657000
rect 149210 656760 149320 657000
rect 149560 656760 149650 657000
rect 149890 656760 149980 657000
rect 150220 656760 150310 657000
rect 150550 656760 150660 657000
rect 150900 656760 150990 657000
rect 151230 656760 151320 657000
rect 151560 656760 151650 657000
rect 151890 656760 152000 657000
rect 152240 656760 152330 657000
rect 152570 656760 152660 657000
rect 152900 656760 152990 657000
rect 153230 656760 153340 657000
rect 153580 656760 153670 657000
rect 153910 656760 154000 657000
rect 154240 656760 154330 657000
rect 154570 656760 154680 657000
rect 154920 656760 155010 657000
rect 155250 656760 155340 657000
rect 155580 656760 155670 657000
rect 155910 656760 155960 657000
rect 110760 656670 155960 656760
rect 110760 656430 110810 656670
rect 111050 656430 111160 656670
rect 111400 656430 111490 656670
rect 111730 656430 111820 656670
rect 112060 656430 112150 656670
rect 112390 656430 112500 656670
rect 112740 656430 112830 656670
rect 113070 656430 113160 656670
rect 113400 656430 113490 656670
rect 113730 656430 113840 656670
rect 114080 656430 114170 656670
rect 114410 656430 114500 656670
rect 114740 656430 114830 656670
rect 115070 656430 115180 656670
rect 115420 656430 115510 656670
rect 115750 656430 115840 656670
rect 116080 656430 116170 656670
rect 116410 656430 116520 656670
rect 116760 656430 116850 656670
rect 117090 656430 117180 656670
rect 117420 656430 117510 656670
rect 117750 656430 117860 656670
rect 118100 656430 118190 656670
rect 118430 656430 118520 656670
rect 118760 656430 118850 656670
rect 119090 656430 119200 656670
rect 119440 656430 119530 656670
rect 119770 656430 119860 656670
rect 120100 656430 120190 656670
rect 120430 656430 120540 656670
rect 120780 656430 120870 656670
rect 121110 656430 121200 656670
rect 121440 656430 121530 656670
rect 121770 656430 122190 656670
rect 122430 656430 122540 656670
rect 122780 656430 122870 656670
rect 123110 656430 123200 656670
rect 123440 656430 123530 656670
rect 123770 656430 123880 656670
rect 124120 656430 124210 656670
rect 124450 656430 124540 656670
rect 124780 656430 124870 656670
rect 125110 656430 125220 656670
rect 125460 656430 125550 656670
rect 125790 656430 125880 656670
rect 126120 656430 126210 656670
rect 126450 656430 126560 656670
rect 126800 656430 126890 656670
rect 127130 656430 127220 656670
rect 127460 656430 127550 656670
rect 127790 656430 127900 656670
rect 128140 656430 128230 656670
rect 128470 656430 128560 656670
rect 128800 656430 128890 656670
rect 129130 656430 129240 656670
rect 129480 656430 129570 656670
rect 129810 656430 129900 656670
rect 130140 656430 130230 656670
rect 130470 656430 130580 656670
rect 130820 656430 130910 656670
rect 131150 656430 131240 656670
rect 131480 656430 131570 656670
rect 131810 656430 131920 656670
rect 132160 656430 132250 656670
rect 132490 656430 132580 656670
rect 132820 656430 132910 656670
rect 133150 656430 133570 656670
rect 133810 656430 133920 656670
rect 134160 656430 134250 656670
rect 134490 656430 134580 656670
rect 134820 656430 134910 656670
rect 135150 656430 135260 656670
rect 135500 656430 135590 656670
rect 135830 656430 135920 656670
rect 136160 656430 136250 656670
rect 136490 656430 136600 656670
rect 136840 656430 136930 656670
rect 137170 656430 137260 656670
rect 137500 656430 137590 656670
rect 137830 656430 137940 656670
rect 138180 656430 138270 656670
rect 138510 656430 138600 656670
rect 138840 656430 138930 656670
rect 139170 656430 139280 656670
rect 139520 656430 139610 656670
rect 139850 656430 139940 656670
rect 140180 656430 140270 656670
rect 140510 656430 140620 656670
rect 140860 656430 140950 656670
rect 141190 656430 141280 656670
rect 141520 656430 141610 656670
rect 141850 656430 141960 656670
rect 142200 656430 142290 656670
rect 142530 656430 142620 656670
rect 142860 656430 142950 656670
rect 143190 656430 143300 656670
rect 143540 656430 143630 656670
rect 143870 656430 143960 656670
rect 144200 656430 144290 656670
rect 144530 656430 144950 656670
rect 145190 656430 145300 656670
rect 145540 656430 145630 656670
rect 145870 656430 145960 656670
rect 146200 656430 146290 656670
rect 146530 656430 146640 656670
rect 146880 656430 146970 656670
rect 147210 656430 147300 656670
rect 147540 656430 147630 656670
rect 147870 656430 147980 656670
rect 148220 656430 148310 656670
rect 148550 656430 148640 656670
rect 148880 656430 148970 656670
rect 149210 656430 149320 656670
rect 149560 656430 149650 656670
rect 149890 656430 149980 656670
rect 150220 656430 150310 656670
rect 150550 656430 150660 656670
rect 150900 656430 150990 656670
rect 151230 656430 151320 656670
rect 151560 656430 151650 656670
rect 151890 656430 152000 656670
rect 152240 656430 152330 656670
rect 152570 656430 152660 656670
rect 152900 656430 152990 656670
rect 153230 656430 153340 656670
rect 153580 656430 153670 656670
rect 153910 656430 154000 656670
rect 154240 656430 154330 656670
rect 154570 656430 154680 656670
rect 154920 656430 155010 656670
rect 155250 656430 155340 656670
rect 155580 656430 155670 656670
rect 155910 656430 155960 656670
rect 110760 656320 155960 656430
rect 110760 656080 110810 656320
rect 111050 656080 111160 656320
rect 111400 656080 111490 656320
rect 111730 656080 111820 656320
rect 112060 656080 112150 656320
rect 112390 656080 112500 656320
rect 112740 656080 112830 656320
rect 113070 656080 113160 656320
rect 113400 656080 113490 656320
rect 113730 656080 113840 656320
rect 114080 656080 114170 656320
rect 114410 656080 114500 656320
rect 114740 656080 114830 656320
rect 115070 656080 115180 656320
rect 115420 656080 115510 656320
rect 115750 656080 115840 656320
rect 116080 656080 116170 656320
rect 116410 656080 116520 656320
rect 116760 656080 116850 656320
rect 117090 656080 117180 656320
rect 117420 656080 117510 656320
rect 117750 656080 117860 656320
rect 118100 656080 118190 656320
rect 118430 656080 118520 656320
rect 118760 656080 118850 656320
rect 119090 656080 119200 656320
rect 119440 656080 119530 656320
rect 119770 656080 119860 656320
rect 120100 656080 120190 656320
rect 120430 656080 120540 656320
rect 120780 656080 120870 656320
rect 121110 656080 121200 656320
rect 121440 656080 121530 656320
rect 121770 656080 122190 656320
rect 122430 656080 122540 656320
rect 122780 656080 122870 656320
rect 123110 656080 123200 656320
rect 123440 656080 123530 656320
rect 123770 656080 123880 656320
rect 124120 656080 124210 656320
rect 124450 656080 124540 656320
rect 124780 656080 124870 656320
rect 125110 656080 125220 656320
rect 125460 656080 125550 656320
rect 125790 656080 125880 656320
rect 126120 656080 126210 656320
rect 126450 656080 126560 656320
rect 126800 656080 126890 656320
rect 127130 656080 127220 656320
rect 127460 656080 127550 656320
rect 127790 656080 127900 656320
rect 128140 656080 128230 656320
rect 128470 656080 128560 656320
rect 128800 656080 128890 656320
rect 129130 656080 129240 656320
rect 129480 656080 129570 656320
rect 129810 656080 129900 656320
rect 130140 656080 130230 656320
rect 130470 656080 130580 656320
rect 130820 656080 130910 656320
rect 131150 656080 131240 656320
rect 131480 656080 131570 656320
rect 131810 656080 131920 656320
rect 132160 656080 132250 656320
rect 132490 656080 132580 656320
rect 132820 656080 132910 656320
rect 133150 656080 133570 656320
rect 133810 656080 133920 656320
rect 134160 656080 134250 656320
rect 134490 656080 134580 656320
rect 134820 656080 134910 656320
rect 135150 656080 135260 656320
rect 135500 656080 135590 656320
rect 135830 656080 135920 656320
rect 136160 656080 136250 656320
rect 136490 656080 136600 656320
rect 136840 656080 136930 656320
rect 137170 656080 137260 656320
rect 137500 656080 137590 656320
rect 137830 656080 137940 656320
rect 138180 656080 138270 656320
rect 138510 656080 138600 656320
rect 138840 656080 138930 656320
rect 139170 656080 139280 656320
rect 139520 656080 139610 656320
rect 139850 656080 139940 656320
rect 140180 656080 140270 656320
rect 140510 656080 140620 656320
rect 140860 656080 140950 656320
rect 141190 656080 141280 656320
rect 141520 656080 141610 656320
rect 141850 656080 141960 656320
rect 142200 656080 142290 656320
rect 142530 656080 142620 656320
rect 142860 656080 142950 656320
rect 143190 656080 143300 656320
rect 143540 656080 143630 656320
rect 143870 656080 143960 656320
rect 144200 656080 144290 656320
rect 144530 656080 144950 656320
rect 145190 656080 145300 656320
rect 145540 656080 145630 656320
rect 145870 656080 145960 656320
rect 146200 656080 146290 656320
rect 146530 656080 146640 656320
rect 146880 656080 146970 656320
rect 147210 656080 147300 656320
rect 147540 656080 147630 656320
rect 147870 656080 147980 656320
rect 148220 656080 148310 656320
rect 148550 656080 148640 656320
rect 148880 656080 148970 656320
rect 149210 656080 149320 656320
rect 149560 656080 149650 656320
rect 149890 656080 149980 656320
rect 150220 656080 150310 656320
rect 150550 656080 150660 656320
rect 150900 656080 150990 656320
rect 151230 656080 151320 656320
rect 151560 656080 151650 656320
rect 151890 656080 152000 656320
rect 152240 656080 152330 656320
rect 152570 656080 152660 656320
rect 152900 656080 152990 656320
rect 153230 656080 153340 656320
rect 153580 656080 153670 656320
rect 153910 656080 154000 656320
rect 154240 656080 154330 656320
rect 154570 656080 154680 656320
rect 154920 656080 155010 656320
rect 155250 656080 155340 656320
rect 155580 656080 155670 656320
rect 155910 656080 155960 656320
rect 110760 655990 155960 656080
rect 110760 655750 110810 655990
rect 111050 655750 111160 655990
rect 111400 655750 111490 655990
rect 111730 655750 111820 655990
rect 112060 655750 112150 655990
rect 112390 655750 112500 655990
rect 112740 655750 112830 655990
rect 113070 655750 113160 655990
rect 113400 655750 113490 655990
rect 113730 655750 113840 655990
rect 114080 655750 114170 655990
rect 114410 655750 114500 655990
rect 114740 655750 114830 655990
rect 115070 655750 115180 655990
rect 115420 655750 115510 655990
rect 115750 655750 115840 655990
rect 116080 655750 116170 655990
rect 116410 655750 116520 655990
rect 116760 655750 116850 655990
rect 117090 655750 117180 655990
rect 117420 655750 117510 655990
rect 117750 655750 117860 655990
rect 118100 655750 118190 655990
rect 118430 655750 118520 655990
rect 118760 655750 118850 655990
rect 119090 655750 119200 655990
rect 119440 655750 119530 655990
rect 119770 655750 119860 655990
rect 120100 655750 120190 655990
rect 120430 655750 120540 655990
rect 120780 655750 120870 655990
rect 121110 655750 121200 655990
rect 121440 655750 121530 655990
rect 121770 655750 122190 655990
rect 122430 655750 122540 655990
rect 122780 655750 122870 655990
rect 123110 655750 123200 655990
rect 123440 655750 123530 655990
rect 123770 655750 123880 655990
rect 124120 655750 124210 655990
rect 124450 655750 124540 655990
rect 124780 655750 124870 655990
rect 125110 655750 125220 655990
rect 125460 655750 125550 655990
rect 125790 655750 125880 655990
rect 126120 655750 126210 655990
rect 126450 655750 126560 655990
rect 126800 655750 126890 655990
rect 127130 655750 127220 655990
rect 127460 655750 127550 655990
rect 127790 655750 127900 655990
rect 128140 655750 128230 655990
rect 128470 655750 128560 655990
rect 128800 655750 128890 655990
rect 129130 655750 129240 655990
rect 129480 655750 129570 655990
rect 129810 655750 129900 655990
rect 130140 655750 130230 655990
rect 130470 655750 130580 655990
rect 130820 655750 130910 655990
rect 131150 655750 131240 655990
rect 131480 655750 131570 655990
rect 131810 655750 131920 655990
rect 132160 655750 132250 655990
rect 132490 655750 132580 655990
rect 132820 655750 132910 655990
rect 133150 655750 133570 655990
rect 133810 655750 133920 655990
rect 134160 655750 134250 655990
rect 134490 655750 134580 655990
rect 134820 655750 134910 655990
rect 135150 655750 135260 655990
rect 135500 655750 135590 655990
rect 135830 655750 135920 655990
rect 136160 655750 136250 655990
rect 136490 655750 136600 655990
rect 136840 655750 136930 655990
rect 137170 655750 137260 655990
rect 137500 655750 137590 655990
rect 137830 655750 137940 655990
rect 138180 655750 138270 655990
rect 138510 655750 138600 655990
rect 138840 655750 138930 655990
rect 139170 655750 139280 655990
rect 139520 655750 139610 655990
rect 139850 655750 139940 655990
rect 140180 655750 140270 655990
rect 140510 655750 140620 655990
rect 140860 655750 140950 655990
rect 141190 655750 141280 655990
rect 141520 655750 141610 655990
rect 141850 655750 141960 655990
rect 142200 655750 142290 655990
rect 142530 655750 142620 655990
rect 142860 655750 142950 655990
rect 143190 655750 143300 655990
rect 143540 655750 143630 655990
rect 143870 655750 143960 655990
rect 144200 655750 144290 655990
rect 144530 655750 144950 655990
rect 145190 655750 145300 655990
rect 145540 655750 145630 655990
rect 145870 655750 145960 655990
rect 146200 655750 146290 655990
rect 146530 655750 146640 655990
rect 146880 655750 146970 655990
rect 147210 655750 147300 655990
rect 147540 655750 147630 655990
rect 147870 655750 147980 655990
rect 148220 655750 148310 655990
rect 148550 655750 148640 655990
rect 148880 655750 148970 655990
rect 149210 655750 149320 655990
rect 149560 655750 149650 655990
rect 149890 655750 149980 655990
rect 150220 655750 150310 655990
rect 150550 655750 150660 655990
rect 150900 655750 150990 655990
rect 151230 655750 151320 655990
rect 151560 655750 151650 655990
rect 151890 655750 152000 655990
rect 152240 655750 152330 655990
rect 152570 655750 152660 655990
rect 152900 655750 152990 655990
rect 153230 655750 153340 655990
rect 153580 655750 153670 655990
rect 153910 655750 154000 655990
rect 154240 655750 154330 655990
rect 154570 655750 154680 655990
rect 154920 655750 155010 655990
rect 155250 655750 155340 655990
rect 155580 655750 155670 655990
rect 155910 655750 155960 655990
rect 110760 655660 155960 655750
rect 110760 655420 110810 655660
rect 111050 655420 111160 655660
rect 111400 655420 111490 655660
rect 111730 655420 111820 655660
rect 112060 655420 112150 655660
rect 112390 655420 112500 655660
rect 112740 655420 112830 655660
rect 113070 655420 113160 655660
rect 113400 655420 113490 655660
rect 113730 655420 113840 655660
rect 114080 655420 114170 655660
rect 114410 655420 114500 655660
rect 114740 655420 114830 655660
rect 115070 655420 115180 655660
rect 115420 655420 115510 655660
rect 115750 655420 115840 655660
rect 116080 655420 116170 655660
rect 116410 655420 116520 655660
rect 116760 655420 116850 655660
rect 117090 655420 117180 655660
rect 117420 655420 117510 655660
rect 117750 655420 117860 655660
rect 118100 655420 118190 655660
rect 118430 655420 118520 655660
rect 118760 655420 118850 655660
rect 119090 655420 119200 655660
rect 119440 655420 119530 655660
rect 119770 655420 119860 655660
rect 120100 655420 120190 655660
rect 120430 655420 120540 655660
rect 120780 655420 120870 655660
rect 121110 655420 121200 655660
rect 121440 655420 121530 655660
rect 121770 655420 122190 655660
rect 122430 655420 122540 655660
rect 122780 655420 122870 655660
rect 123110 655420 123200 655660
rect 123440 655420 123530 655660
rect 123770 655420 123880 655660
rect 124120 655420 124210 655660
rect 124450 655420 124540 655660
rect 124780 655420 124870 655660
rect 125110 655420 125220 655660
rect 125460 655420 125550 655660
rect 125790 655420 125880 655660
rect 126120 655420 126210 655660
rect 126450 655420 126560 655660
rect 126800 655420 126890 655660
rect 127130 655420 127220 655660
rect 127460 655420 127550 655660
rect 127790 655420 127900 655660
rect 128140 655420 128230 655660
rect 128470 655420 128560 655660
rect 128800 655420 128890 655660
rect 129130 655420 129240 655660
rect 129480 655420 129570 655660
rect 129810 655420 129900 655660
rect 130140 655420 130230 655660
rect 130470 655420 130580 655660
rect 130820 655420 130910 655660
rect 131150 655420 131240 655660
rect 131480 655420 131570 655660
rect 131810 655420 131920 655660
rect 132160 655420 132250 655660
rect 132490 655420 132580 655660
rect 132820 655420 132910 655660
rect 133150 655420 133570 655660
rect 133810 655420 133920 655660
rect 134160 655420 134250 655660
rect 134490 655420 134580 655660
rect 134820 655420 134910 655660
rect 135150 655420 135260 655660
rect 135500 655420 135590 655660
rect 135830 655420 135920 655660
rect 136160 655420 136250 655660
rect 136490 655420 136600 655660
rect 136840 655420 136930 655660
rect 137170 655420 137260 655660
rect 137500 655420 137590 655660
rect 137830 655420 137940 655660
rect 138180 655420 138270 655660
rect 138510 655420 138600 655660
rect 138840 655420 138930 655660
rect 139170 655420 139280 655660
rect 139520 655420 139610 655660
rect 139850 655420 139940 655660
rect 140180 655420 140270 655660
rect 140510 655420 140620 655660
rect 140860 655420 140950 655660
rect 141190 655420 141280 655660
rect 141520 655420 141610 655660
rect 141850 655420 141960 655660
rect 142200 655420 142290 655660
rect 142530 655420 142620 655660
rect 142860 655420 142950 655660
rect 143190 655420 143300 655660
rect 143540 655420 143630 655660
rect 143870 655420 143960 655660
rect 144200 655420 144290 655660
rect 144530 655420 144950 655660
rect 145190 655420 145300 655660
rect 145540 655420 145630 655660
rect 145870 655420 145960 655660
rect 146200 655420 146290 655660
rect 146530 655420 146640 655660
rect 146880 655420 146970 655660
rect 147210 655420 147300 655660
rect 147540 655420 147630 655660
rect 147870 655420 147980 655660
rect 148220 655420 148310 655660
rect 148550 655420 148640 655660
rect 148880 655420 148970 655660
rect 149210 655420 149320 655660
rect 149560 655420 149650 655660
rect 149890 655420 149980 655660
rect 150220 655420 150310 655660
rect 150550 655420 150660 655660
rect 150900 655420 150990 655660
rect 151230 655420 151320 655660
rect 151560 655420 151650 655660
rect 151890 655420 152000 655660
rect 152240 655420 152330 655660
rect 152570 655420 152660 655660
rect 152900 655420 152990 655660
rect 153230 655420 153340 655660
rect 153580 655420 153670 655660
rect 153910 655420 154000 655660
rect 154240 655420 154330 655660
rect 154570 655420 154680 655660
rect 154920 655420 155010 655660
rect 155250 655420 155340 655660
rect 155580 655420 155670 655660
rect 155910 655420 155960 655660
rect 110760 655330 155960 655420
rect 110760 655090 110810 655330
rect 111050 655090 111160 655330
rect 111400 655090 111490 655330
rect 111730 655090 111820 655330
rect 112060 655090 112150 655330
rect 112390 655090 112500 655330
rect 112740 655090 112830 655330
rect 113070 655090 113160 655330
rect 113400 655090 113490 655330
rect 113730 655090 113840 655330
rect 114080 655090 114170 655330
rect 114410 655090 114500 655330
rect 114740 655090 114830 655330
rect 115070 655090 115180 655330
rect 115420 655090 115510 655330
rect 115750 655090 115840 655330
rect 116080 655090 116170 655330
rect 116410 655090 116520 655330
rect 116760 655090 116850 655330
rect 117090 655090 117180 655330
rect 117420 655090 117510 655330
rect 117750 655090 117860 655330
rect 118100 655090 118190 655330
rect 118430 655090 118520 655330
rect 118760 655090 118850 655330
rect 119090 655090 119200 655330
rect 119440 655090 119530 655330
rect 119770 655090 119860 655330
rect 120100 655090 120190 655330
rect 120430 655090 120540 655330
rect 120780 655090 120870 655330
rect 121110 655090 121200 655330
rect 121440 655090 121530 655330
rect 121770 655090 122190 655330
rect 122430 655090 122540 655330
rect 122780 655090 122870 655330
rect 123110 655090 123200 655330
rect 123440 655090 123530 655330
rect 123770 655090 123880 655330
rect 124120 655090 124210 655330
rect 124450 655090 124540 655330
rect 124780 655090 124870 655330
rect 125110 655090 125220 655330
rect 125460 655090 125550 655330
rect 125790 655090 125880 655330
rect 126120 655090 126210 655330
rect 126450 655090 126560 655330
rect 126800 655090 126890 655330
rect 127130 655090 127220 655330
rect 127460 655090 127550 655330
rect 127790 655090 127900 655330
rect 128140 655090 128230 655330
rect 128470 655090 128560 655330
rect 128800 655090 128890 655330
rect 129130 655090 129240 655330
rect 129480 655090 129570 655330
rect 129810 655090 129900 655330
rect 130140 655090 130230 655330
rect 130470 655090 130580 655330
rect 130820 655090 130910 655330
rect 131150 655090 131240 655330
rect 131480 655090 131570 655330
rect 131810 655090 131920 655330
rect 132160 655090 132250 655330
rect 132490 655090 132580 655330
rect 132820 655090 132910 655330
rect 133150 655090 133570 655330
rect 133810 655090 133920 655330
rect 134160 655090 134250 655330
rect 134490 655090 134580 655330
rect 134820 655090 134910 655330
rect 135150 655090 135260 655330
rect 135500 655090 135590 655330
rect 135830 655090 135920 655330
rect 136160 655090 136250 655330
rect 136490 655090 136600 655330
rect 136840 655090 136930 655330
rect 137170 655090 137260 655330
rect 137500 655090 137590 655330
rect 137830 655090 137940 655330
rect 138180 655090 138270 655330
rect 138510 655090 138600 655330
rect 138840 655090 138930 655330
rect 139170 655090 139280 655330
rect 139520 655090 139610 655330
rect 139850 655090 139940 655330
rect 140180 655090 140270 655330
rect 140510 655090 140620 655330
rect 140860 655090 140950 655330
rect 141190 655090 141280 655330
rect 141520 655090 141610 655330
rect 141850 655090 141960 655330
rect 142200 655090 142290 655330
rect 142530 655090 142620 655330
rect 142860 655090 142950 655330
rect 143190 655090 143300 655330
rect 143540 655090 143630 655330
rect 143870 655090 143960 655330
rect 144200 655090 144290 655330
rect 144530 655090 144950 655330
rect 145190 655090 145300 655330
rect 145540 655090 145630 655330
rect 145870 655090 145960 655330
rect 146200 655090 146290 655330
rect 146530 655090 146640 655330
rect 146880 655090 146970 655330
rect 147210 655090 147300 655330
rect 147540 655090 147630 655330
rect 147870 655090 147980 655330
rect 148220 655090 148310 655330
rect 148550 655090 148640 655330
rect 148880 655090 148970 655330
rect 149210 655090 149320 655330
rect 149560 655090 149650 655330
rect 149890 655090 149980 655330
rect 150220 655090 150310 655330
rect 150550 655090 150660 655330
rect 150900 655090 150990 655330
rect 151230 655090 151320 655330
rect 151560 655090 151650 655330
rect 151890 655090 152000 655330
rect 152240 655090 152330 655330
rect 152570 655090 152660 655330
rect 152900 655090 152990 655330
rect 153230 655090 153340 655330
rect 153580 655090 153670 655330
rect 153910 655090 154000 655330
rect 154240 655090 154330 655330
rect 154570 655090 154680 655330
rect 154920 655090 155010 655330
rect 155250 655090 155340 655330
rect 155580 655090 155670 655330
rect 155910 655090 155960 655330
rect 110760 654980 155960 655090
rect 110760 654740 110810 654980
rect 111050 654740 111160 654980
rect 111400 654740 111490 654980
rect 111730 654740 111820 654980
rect 112060 654740 112150 654980
rect 112390 654740 112500 654980
rect 112740 654740 112830 654980
rect 113070 654740 113160 654980
rect 113400 654740 113490 654980
rect 113730 654740 113840 654980
rect 114080 654740 114170 654980
rect 114410 654740 114500 654980
rect 114740 654740 114830 654980
rect 115070 654740 115180 654980
rect 115420 654740 115510 654980
rect 115750 654740 115840 654980
rect 116080 654740 116170 654980
rect 116410 654740 116520 654980
rect 116760 654740 116850 654980
rect 117090 654740 117180 654980
rect 117420 654740 117510 654980
rect 117750 654740 117860 654980
rect 118100 654740 118190 654980
rect 118430 654740 118520 654980
rect 118760 654740 118850 654980
rect 119090 654740 119200 654980
rect 119440 654740 119530 654980
rect 119770 654740 119860 654980
rect 120100 654740 120190 654980
rect 120430 654740 120540 654980
rect 120780 654740 120870 654980
rect 121110 654740 121200 654980
rect 121440 654740 121530 654980
rect 121770 654740 122190 654980
rect 122430 654740 122540 654980
rect 122780 654740 122870 654980
rect 123110 654740 123200 654980
rect 123440 654740 123530 654980
rect 123770 654740 123880 654980
rect 124120 654740 124210 654980
rect 124450 654740 124540 654980
rect 124780 654740 124870 654980
rect 125110 654740 125220 654980
rect 125460 654740 125550 654980
rect 125790 654740 125880 654980
rect 126120 654740 126210 654980
rect 126450 654740 126560 654980
rect 126800 654740 126890 654980
rect 127130 654740 127220 654980
rect 127460 654740 127550 654980
rect 127790 654740 127900 654980
rect 128140 654740 128230 654980
rect 128470 654740 128560 654980
rect 128800 654740 128890 654980
rect 129130 654740 129240 654980
rect 129480 654740 129570 654980
rect 129810 654740 129900 654980
rect 130140 654740 130230 654980
rect 130470 654740 130580 654980
rect 130820 654740 130910 654980
rect 131150 654740 131240 654980
rect 131480 654740 131570 654980
rect 131810 654740 131920 654980
rect 132160 654740 132250 654980
rect 132490 654740 132580 654980
rect 132820 654740 132910 654980
rect 133150 654740 133570 654980
rect 133810 654740 133920 654980
rect 134160 654740 134250 654980
rect 134490 654740 134580 654980
rect 134820 654740 134910 654980
rect 135150 654740 135260 654980
rect 135500 654740 135590 654980
rect 135830 654740 135920 654980
rect 136160 654740 136250 654980
rect 136490 654740 136600 654980
rect 136840 654740 136930 654980
rect 137170 654740 137260 654980
rect 137500 654740 137590 654980
rect 137830 654740 137940 654980
rect 138180 654740 138270 654980
rect 138510 654740 138600 654980
rect 138840 654740 138930 654980
rect 139170 654740 139280 654980
rect 139520 654740 139610 654980
rect 139850 654740 139940 654980
rect 140180 654740 140270 654980
rect 140510 654740 140620 654980
rect 140860 654740 140950 654980
rect 141190 654740 141280 654980
rect 141520 654740 141610 654980
rect 141850 654740 141960 654980
rect 142200 654740 142290 654980
rect 142530 654740 142620 654980
rect 142860 654740 142950 654980
rect 143190 654740 143300 654980
rect 143540 654740 143630 654980
rect 143870 654740 143960 654980
rect 144200 654740 144290 654980
rect 144530 654740 144950 654980
rect 145190 654740 145300 654980
rect 145540 654740 145630 654980
rect 145870 654740 145960 654980
rect 146200 654740 146290 654980
rect 146530 654740 146640 654980
rect 146880 654740 146970 654980
rect 147210 654740 147300 654980
rect 147540 654740 147630 654980
rect 147870 654740 147980 654980
rect 148220 654740 148310 654980
rect 148550 654740 148640 654980
rect 148880 654740 148970 654980
rect 149210 654740 149320 654980
rect 149560 654740 149650 654980
rect 149890 654740 149980 654980
rect 150220 654740 150310 654980
rect 150550 654740 150660 654980
rect 150900 654740 150990 654980
rect 151230 654740 151320 654980
rect 151560 654740 151650 654980
rect 151890 654740 152000 654980
rect 152240 654740 152330 654980
rect 152570 654740 152660 654980
rect 152900 654740 152990 654980
rect 153230 654740 153340 654980
rect 153580 654740 153670 654980
rect 153910 654740 154000 654980
rect 154240 654740 154330 654980
rect 154570 654740 154680 654980
rect 154920 654740 155010 654980
rect 155250 654740 155340 654980
rect 155580 654740 155670 654980
rect 155910 654740 155960 654980
rect 110760 654650 155960 654740
rect 110760 654410 110810 654650
rect 111050 654410 111160 654650
rect 111400 654410 111490 654650
rect 111730 654410 111820 654650
rect 112060 654410 112150 654650
rect 112390 654410 112500 654650
rect 112740 654410 112830 654650
rect 113070 654410 113160 654650
rect 113400 654410 113490 654650
rect 113730 654410 113840 654650
rect 114080 654410 114170 654650
rect 114410 654410 114500 654650
rect 114740 654410 114830 654650
rect 115070 654410 115180 654650
rect 115420 654410 115510 654650
rect 115750 654410 115840 654650
rect 116080 654410 116170 654650
rect 116410 654410 116520 654650
rect 116760 654410 116850 654650
rect 117090 654410 117180 654650
rect 117420 654410 117510 654650
rect 117750 654410 117860 654650
rect 118100 654410 118190 654650
rect 118430 654410 118520 654650
rect 118760 654410 118850 654650
rect 119090 654410 119200 654650
rect 119440 654410 119530 654650
rect 119770 654410 119860 654650
rect 120100 654410 120190 654650
rect 120430 654410 120540 654650
rect 120780 654410 120870 654650
rect 121110 654410 121200 654650
rect 121440 654410 121530 654650
rect 121770 654410 122190 654650
rect 122430 654410 122540 654650
rect 122780 654410 122870 654650
rect 123110 654410 123200 654650
rect 123440 654410 123530 654650
rect 123770 654410 123880 654650
rect 124120 654410 124210 654650
rect 124450 654410 124540 654650
rect 124780 654410 124870 654650
rect 125110 654410 125220 654650
rect 125460 654410 125550 654650
rect 125790 654410 125880 654650
rect 126120 654410 126210 654650
rect 126450 654410 126560 654650
rect 126800 654410 126890 654650
rect 127130 654410 127220 654650
rect 127460 654410 127550 654650
rect 127790 654410 127900 654650
rect 128140 654410 128230 654650
rect 128470 654410 128560 654650
rect 128800 654410 128890 654650
rect 129130 654410 129240 654650
rect 129480 654410 129570 654650
rect 129810 654410 129900 654650
rect 130140 654410 130230 654650
rect 130470 654410 130580 654650
rect 130820 654410 130910 654650
rect 131150 654410 131240 654650
rect 131480 654410 131570 654650
rect 131810 654410 131920 654650
rect 132160 654410 132250 654650
rect 132490 654410 132580 654650
rect 132820 654410 132910 654650
rect 133150 654410 133570 654650
rect 133810 654410 133920 654650
rect 134160 654410 134250 654650
rect 134490 654410 134580 654650
rect 134820 654410 134910 654650
rect 135150 654410 135260 654650
rect 135500 654410 135590 654650
rect 135830 654410 135920 654650
rect 136160 654410 136250 654650
rect 136490 654410 136600 654650
rect 136840 654410 136930 654650
rect 137170 654410 137260 654650
rect 137500 654410 137590 654650
rect 137830 654410 137940 654650
rect 138180 654410 138270 654650
rect 138510 654410 138600 654650
rect 138840 654410 138930 654650
rect 139170 654410 139280 654650
rect 139520 654410 139610 654650
rect 139850 654410 139940 654650
rect 140180 654410 140270 654650
rect 140510 654410 140620 654650
rect 140860 654410 140950 654650
rect 141190 654410 141280 654650
rect 141520 654410 141610 654650
rect 141850 654410 141960 654650
rect 142200 654410 142290 654650
rect 142530 654410 142620 654650
rect 142860 654410 142950 654650
rect 143190 654410 143300 654650
rect 143540 654410 143630 654650
rect 143870 654410 143960 654650
rect 144200 654410 144290 654650
rect 144530 654410 144950 654650
rect 145190 654410 145300 654650
rect 145540 654410 145630 654650
rect 145870 654410 145960 654650
rect 146200 654410 146290 654650
rect 146530 654410 146640 654650
rect 146880 654410 146970 654650
rect 147210 654410 147300 654650
rect 147540 654410 147630 654650
rect 147870 654410 147980 654650
rect 148220 654410 148310 654650
rect 148550 654410 148640 654650
rect 148880 654410 148970 654650
rect 149210 654410 149320 654650
rect 149560 654410 149650 654650
rect 149890 654410 149980 654650
rect 150220 654410 150310 654650
rect 150550 654410 150660 654650
rect 150900 654410 150990 654650
rect 151230 654410 151320 654650
rect 151560 654410 151650 654650
rect 151890 654410 152000 654650
rect 152240 654410 152330 654650
rect 152570 654410 152660 654650
rect 152900 654410 152990 654650
rect 153230 654410 153340 654650
rect 153580 654410 153670 654650
rect 153910 654410 154000 654650
rect 154240 654410 154330 654650
rect 154570 654410 154680 654650
rect 154920 654410 155010 654650
rect 155250 654410 155340 654650
rect 155580 654410 155670 654650
rect 155910 654410 155960 654650
rect 110760 654320 155960 654410
rect 110760 654080 110810 654320
rect 111050 654080 111160 654320
rect 111400 654080 111490 654320
rect 111730 654080 111820 654320
rect 112060 654080 112150 654320
rect 112390 654080 112500 654320
rect 112740 654080 112830 654320
rect 113070 654080 113160 654320
rect 113400 654080 113490 654320
rect 113730 654080 113840 654320
rect 114080 654080 114170 654320
rect 114410 654080 114500 654320
rect 114740 654080 114830 654320
rect 115070 654080 115180 654320
rect 115420 654080 115510 654320
rect 115750 654080 115840 654320
rect 116080 654080 116170 654320
rect 116410 654080 116520 654320
rect 116760 654080 116850 654320
rect 117090 654080 117180 654320
rect 117420 654080 117510 654320
rect 117750 654080 117860 654320
rect 118100 654080 118190 654320
rect 118430 654080 118520 654320
rect 118760 654080 118850 654320
rect 119090 654080 119200 654320
rect 119440 654080 119530 654320
rect 119770 654080 119860 654320
rect 120100 654080 120190 654320
rect 120430 654080 120540 654320
rect 120780 654080 120870 654320
rect 121110 654080 121200 654320
rect 121440 654080 121530 654320
rect 121770 654080 122190 654320
rect 122430 654080 122540 654320
rect 122780 654080 122870 654320
rect 123110 654080 123200 654320
rect 123440 654080 123530 654320
rect 123770 654080 123880 654320
rect 124120 654080 124210 654320
rect 124450 654080 124540 654320
rect 124780 654080 124870 654320
rect 125110 654080 125220 654320
rect 125460 654080 125550 654320
rect 125790 654080 125880 654320
rect 126120 654080 126210 654320
rect 126450 654080 126560 654320
rect 126800 654080 126890 654320
rect 127130 654080 127220 654320
rect 127460 654080 127550 654320
rect 127790 654080 127900 654320
rect 128140 654080 128230 654320
rect 128470 654080 128560 654320
rect 128800 654080 128890 654320
rect 129130 654080 129240 654320
rect 129480 654080 129570 654320
rect 129810 654080 129900 654320
rect 130140 654080 130230 654320
rect 130470 654080 130580 654320
rect 130820 654080 130910 654320
rect 131150 654080 131240 654320
rect 131480 654080 131570 654320
rect 131810 654080 131920 654320
rect 132160 654080 132250 654320
rect 132490 654080 132580 654320
rect 132820 654080 132910 654320
rect 133150 654080 133570 654320
rect 133810 654080 133920 654320
rect 134160 654080 134250 654320
rect 134490 654080 134580 654320
rect 134820 654080 134910 654320
rect 135150 654080 135260 654320
rect 135500 654080 135590 654320
rect 135830 654080 135920 654320
rect 136160 654080 136250 654320
rect 136490 654080 136600 654320
rect 136840 654080 136930 654320
rect 137170 654080 137260 654320
rect 137500 654080 137590 654320
rect 137830 654080 137940 654320
rect 138180 654080 138270 654320
rect 138510 654080 138600 654320
rect 138840 654080 138930 654320
rect 139170 654080 139280 654320
rect 139520 654080 139610 654320
rect 139850 654080 139940 654320
rect 140180 654080 140270 654320
rect 140510 654080 140620 654320
rect 140860 654080 140950 654320
rect 141190 654080 141280 654320
rect 141520 654080 141610 654320
rect 141850 654080 141960 654320
rect 142200 654080 142290 654320
rect 142530 654080 142620 654320
rect 142860 654080 142950 654320
rect 143190 654080 143300 654320
rect 143540 654080 143630 654320
rect 143870 654080 143960 654320
rect 144200 654080 144290 654320
rect 144530 654080 144950 654320
rect 145190 654080 145300 654320
rect 145540 654080 145630 654320
rect 145870 654080 145960 654320
rect 146200 654080 146290 654320
rect 146530 654080 146640 654320
rect 146880 654080 146970 654320
rect 147210 654080 147300 654320
rect 147540 654080 147630 654320
rect 147870 654080 147980 654320
rect 148220 654080 148310 654320
rect 148550 654080 148640 654320
rect 148880 654080 148970 654320
rect 149210 654080 149320 654320
rect 149560 654080 149650 654320
rect 149890 654080 149980 654320
rect 150220 654080 150310 654320
rect 150550 654080 150660 654320
rect 150900 654080 150990 654320
rect 151230 654080 151320 654320
rect 151560 654080 151650 654320
rect 151890 654080 152000 654320
rect 152240 654080 152330 654320
rect 152570 654080 152660 654320
rect 152900 654080 152990 654320
rect 153230 654080 153340 654320
rect 153580 654080 153670 654320
rect 153910 654080 154000 654320
rect 154240 654080 154330 654320
rect 154570 654080 154680 654320
rect 154920 654080 155010 654320
rect 155250 654080 155340 654320
rect 155580 654080 155670 654320
rect 155910 654080 155960 654320
rect 110760 653990 155960 654080
rect 110760 653750 110810 653990
rect 111050 653750 111160 653990
rect 111400 653750 111490 653990
rect 111730 653750 111820 653990
rect 112060 653750 112150 653990
rect 112390 653750 112500 653990
rect 112740 653750 112830 653990
rect 113070 653750 113160 653990
rect 113400 653750 113490 653990
rect 113730 653750 113840 653990
rect 114080 653750 114170 653990
rect 114410 653750 114500 653990
rect 114740 653750 114830 653990
rect 115070 653750 115180 653990
rect 115420 653750 115510 653990
rect 115750 653750 115840 653990
rect 116080 653750 116170 653990
rect 116410 653750 116520 653990
rect 116760 653750 116850 653990
rect 117090 653750 117180 653990
rect 117420 653750 117510 653990
rect 117750 653750 117860 653990
rect 118100 653750 118190 653990
rect 118430 653750 118520 653990
rect 118760 653750 118850 653990
rect 119090 653750 119200 653990
rect 119440 653750 119530 653990
rect 119770 653750 119860 653990
rect 120100 653750 120190 653990
rect 120430 653750 120540 653990
rect 120780 653750 120870 653990
rect 121110 653750 121200 653990
rect 121440 653750 121530 653990
rect 121770 653750 122190 653990
rect 122430 653750 122540 653990
rect 122780 653750 122870 653990
rect 123110 653750 123200 653990
rect 123440 653750 123530 653990
rect 123770 653750 123880 653990
rect 124120 653750 124210 653990
rect 124450 653750 124540 653990
rect 124780 653750 124870 653990
rect 125110 653750 125220 653990
rect 125460 653750 125550 653990
rect 125790 653750 125880 653990
rect 126120 653750 126210 653990
rect 126450 653750 126560 653990
rect 126800 653750 126890 653990
rect 127130 653750 127220 653990
rect 127460 653750 127550 653990
rect 127790 653750 127900 653990
rect 128140 653750 128230 653990
rect 128470 653750 128560 653990
rect 128800 653750 128890 653990
rect 129130 653750 129240 653990
rect 129480 653750 129570 653990
rect 129810 653750 129900 653990
rect 130140 653750 130230 653990
rect 130470 653750 130580 653990
rect 130820 653750 130910 653990
rect 131150 653750 131240 653990
rect 131480 653750 131570 653990
rect 131810 653750 131920 653990
rect 132160 653750 132250 653990
rect 132490 653750 132580 653990
rect 132820 653750 132910 653990
rect 133150 653750 133570 653990
rect 133810 653750 133920 653990
rect 134160 653750 134250 653990
rect 134490 653750 134580 653990
rect 134820 653750 134910 653990
rect 135150 653750 135260 653990
rect 135500 653750 135590 653990
rect 135830 653750 135920 653990
rect 136160 653750 136250 653990
rect 136490 653750 136600 653990
rect 136840 653750 136930 653990
rect 137170 653750 137260 653990
rect 137500 653750 137590 653990
rect 137830 653750 137940 653990
rect 138180 653750 138270 653990
rect 138510 653750 138600 653990
rect 138840 653750 138930 653990
rect 139170 653750 139280 653990
rect 139520 653750 139610 653990
rect 139850 653750 139940 653990
rect 140180 653750 140270 653990
rect 140510 653750 140620 653990
rect 140860 653750 140950 653990
rect 141190 653750 141280 653990
rect 141520 653750 141610 653990
rect 141850 653750 141960 653990
rect 142200 653750 142290 653990
rect 142530 653750 142620 653990
rect 142860 653750 142950 653990
rect 143190 653750 143300 653990
rect 143540 653750 143630 653990
rect 143870 653750 143960 653990
rect 144200 653750 144290 653990
rect 144530 653750 144950 653990
rect 145190 653750 145300 653990
rect 145540 653750 145630 653990
rect 145870 653750 145960 653990
rect 146200 653750 146290 653990
rect 146530 653750 146640 653990
rect 146880 653750 146970 653990
rect 147210 653750 147300 653990
rect 147540 653750 147630 653990
rect 147870 653750 147980 653990
rect 148220 653750 148310 653990
rect 148550 653750 148640 653990
rect 148880 653750 148970 653990
rect 149210 653750 149320 653990
rect 149560 653750 149650 653990
rect 149890 653750 149980 653990
rect 150220 653750 150310 653990
rect 150550 653750 150660 653990
rect 150900 653750 150990 653990
rect 151230 653750 151320 653990
rect 151560 653750 151650 653990
rect 151890 653750 152000 653990
rect 152240 653750 152330 653990
rect 152570 653750 152660 653990
rect 152900 653750 152990 653990
rect 153230 653750 153340 653990
rect 153580 653750 153670 653990
rect 153910 653750 154000 653990
rect 154240 653750 154330 653990
rect 154570 653750 154680 653990
rect 154920 653750 155010 653990
rect 155250 653750 155340 653990
rect 155580 653750 155670 653990
rect 155910 653750 155960 653990
rect 110760 653640 155960 653750
rect 110760 653400 110810 653640
rect 111050 653400 111160 653640
rect 111400 653400 111490 653640
rect 111730 653400 111820 653640
rect 112060 653400 112150 653640
rect 112390 653400 112500 653640
rect 112740 653400 112830 653640
rect 113070 653400 113160 653640
rect 113400 653400 113490 653640
rect 113730 653400 113840 653640
rect 114080 653400 114170 653640
rect 114410 653400 114500 653640
rect 114740 653400 114830 653640
rect 115070 653400 115180 653640
rect 115420 653400 115510 653640
rect 115750 653400 115840 653640
rect 116080 653400 116170 653640
rect 116410 653400 116520 653640
rect 116760 653400 116850 653640
rect 117090 653400 117180 653640
rect 117420 653400 117510 653640
rect 117750 653400 117860 653640
rect 118100 653400 118190 653640
rect 118430 653400 118520 653640
rect 118760 653400 118850 653640
rect 119090 653400 119200 653640
rect 119440 653400 119530 653640
rect 119770 653400 119860 653640
rect 120100 653400 120190 653640
rect 120430 653400 120540 653640
rect 120780 653400 120870 653640
rect 121110 653400 121200 653640
rect 121440 653400 121530 653640
rect 121770 653400 122190 653640
rect 122430 653400 122540 653640
rect 122780 653400 122870 653640
rect 123110 653400 123200 653640
rect 123440 653400 123530 653640
rect 123770 653400 123880 653640
rect 124120 653400 124210 653640
rect 124450 653400 124540 653640
rect 124780 653400 124870 653640
rect 125110 653400 125220 653640
rect 125460 653400 125550 653640
rect 125790 653400 125880 653640
rect 126120 653400 126210 653640
rect 126450 653400 126560 653640
rect 126800 653400 126890 653640
rect 127130 653400 127220 653640
rect 127460 653400 127550 653640
rect 127790 653400 127900 653640
rect 128140 653400 128230 653640
rect 128470 653400 128560 653640
rect 128800 653400 128890 653640
rect 129130 653400 129240 653640
rect 129480 653400 129570 653640
rect 129810 653400 129900 653640
rect 130140 653400 130230 653640
rect 130470 653400 130580 653640
rect 130820 653400 130910 653640
rect 131150 653400 131240 653640
rect 131480 653400 131570 653640
rect 131810 653400 131920 653640
rect 132160 653400 132250 653640
rect 132490 653400 132580 653640
rect 132820 653400 132910 653640
rect 133150 653400 133570 653640
rect 133810 653400 133920 653640
rect 134160 653400 134250 653640
rect 134490 653400 134580 653640
rect 134820 653400 134910 653640
rect 135150 653400 135260 653640
rect 135500 653400 135590 653640
rect 135830 653400 135920 653640
rect 136160 653400 136250 653640
rect 136490 653400 136600 653640
rect 136840 653400 136930 653640
rect 137170 653400 137260 653640
rect 137500 653400 137590 653640
rect 137830 653400 137940 653640
rect 138180 653400 138270 653640
rect 138510 653400 138600 653640
rect 138840 653400 138930 653640
rect 139170 653400 139280 653640
rect 139520 653400 139610 653640
rect 139850 653400 139940 653640
rect 140180 653400 140270 653640
rect 140510 653400 140620 653640
rect 140860 653400 140950 653640
rect 141190 653400 141280 653640
rect 141520 653400 141610 653640
rect 141850 653400 141960 653640
rect 142200 653400 142290 653640
rect 142530 653400 142620 653640
rect 142860 653400 142950 653640
rect 143190 653400 143300 653640
rect 143540 653400 143630 653640
rect 143870 653400 143960 653640
rect 144200 653400 144290 653640
rect 144530 653400 144950 653640
rect 145190 653400 145300 653640
rect 145540 653400 145630 653640
rect 145870 653400 145960 653640
rect 146200 653400 146290 653640
rect 146530 653400 146640 653640
rect 146880 653400 146970 653640
rect 147210 653400 147300 653640
rect 147540 653400 147630 653640
rect 147870 653400 147980 653640
rect 148220 653400 148310 653640
rect 148550 653400 148640 653640
rect 148880 653400 148970 653640
rect 149210 653400 149320 653640
rect 149560 653400 149650 653640
rect 149890 653400 149980 653640
rect 150220 653400 150310 653640
rect 150550 653400 150660 653640
rect 150900 653400 150990 653640
rect 151230 653400 151320 653640
rect 151560 653400 151650 653640
rect 151890 653400 152000 653640
rect 152240 653400 152330 653640
rect 152570 653400 152660 653640
rect 152900 653400 152990 653640
rect 153230 653400 153340 653640
rect 153580 653400 153670 653640
rect 153910 653400 154000 653640
rect 154240 653400 154330 653640
rect 154570 653400 154680 653640
rect 154920 653400 155010 653640
rect 155250 653400 155340 653640
rect 155580 653400 155670 653640
rect 155910 653400 155960 653640
rect 110760 653310 155960 653400
rect 110760 653070 110810 653310
rect 111050 653070 111160 653310
rect 111400 653070 111490 653310
rect 111730 653070 111820 653310
rect 112060 653070 112150 653310
rect 112390 653070 112500 653310
rect 112740 653070 112830 653310
rect 113070 653070 113160 653310
rect 113400 653070 113490 653310
rect 113730 653070 113840 653310
rect 114080 653070 114170 653310
rect 114410 653070 114500 653310
rect 114740 653070 114830 653310
rect 115070 653070 115180 653310
rect 115420 653070 115510 653310
rect 115750 653070 115840 653310
rect 116080 653070 116170 653310
rect 116410 653070 116520 653310
rect 116760 653070 116850 653310
rect 117090 653070 117180 653310
rect 117420 653070 117510 653310
rect 117750 653070 117860 653310
rect 118100 653070 118190 653310
rect 118430 653070 118520 653310
rect 118760 653070 118850 653310
rect 119090 653070 119200 653310
rect 119440 653070 119530 653310
rect 119770 653070 119860 653310
rect 120100 653070 120190 653310
rect 120430 653070 120540 653310
rect 120780 653070 120870 653310
rect 121110 653070 121200 653310
rect 121440 653070 121530 653310
rect 121770 653070 122190 653310
rect 122430 653070 122540 653310
rect 122780 653070 122870 653310
rect 123110 653070 123200 653310
rect 123440 653070 123530 653310
rect 123770 653070 123880 653310
rect 124120 653070 124210 653310
rect 124450 653070 124540 653310
rect 124780 653070 124870 653310
rect 125110 653070 125220 653310
rect 125460 653070 125550 653310
rect 125790 653070 125880 653310
rect 126120 653070 126210 653310
rect 126450 653070 126560 653310
rect 126800 653070 126890 653310
rect 127130 653070 127220 653310
rect 127460 653070 127550 653310
rect 127790 653070 127900 653310
rect 128140 653070 128230 653310
rect 128470 653070 128560 653310
rect 128800 653070 128890 653310
rect 129130 653070 129240 653310
rect 129480 653070 129570 653310
rect 129810 653070 129900 653310
rect 130140 653070 130230 653310
rect 130470 653070 130580 653310
rect 130820 653070 130910 653310
rect 131150 653070 131240 653310
rect 131480 653070 131570 653310
rect 131810 653070 131920 653310
rect 132160 653070 132250 653310
rect 132490 653070 132580 653310
rect 132820 653070 132910 653310
rect 133150 653070 133570 653310
rect 133810 653070 133920 653310
rect 134160 653070 134250 653310
rect 134490 653070 134580 653310
rect 134820 653070 134910 653310
rect 135150 653070 135260 653310
rect 135500 653070 135590 653310
rect 135830 653070 135920 653310
rect 136160 653070 136250 653310
rect 136490 653070 136600 653310
rect 136840 653070 136930 653310
rect 137170 653070 137260 653310
rect 137500 653070 137590 653310
rect 137830 653070 137940 653310
rect 138180 653070 138270 653310
rect 138510 653070 138600 653310
rect 138840 653070 138930 653310
rect 139170 653070 139280 653310
rect 139520 653070 139610 653310
rect 139850 653070 139940 653310
rect 140180 653070 140270 653310
rect 140510 653070 140620 653310
rect 140860 653070 140950 653310
rect 141190 653070 141280 653310
rect 141520 653070 141610 653310
rect 141850 653070 141960 653310
rect 142200 653070 142290 653310
rect 142530 653070 142620 653310
rect 142860 653070 142950 653310
rect 143190 653070 143300 653310
rect 143540 653070 143630 653310
rect 143870 653070 143960 653310
rect 144200 653070 144290 653310
rect 144530 653070 144950 653310
rect 145190 653070 145300 653310
rect 145540 653070 145630 653310
rect 145870 653070 145960 653310
rect 146200 653070 146290 653310
rect 146530 653070 146640 653310
rect 146880 653070 146970 653310
rect 147210 653070 147300 653310
rect 147540 653070 147630 653310
rect 147870 653070 147980 653310
rect 148220 653070 148310 653310
rect 148550 653070 148640 653310
rect 148880 653070 148970 653310
rect 149210 653070 149320 653310
rect 149560 653070 149650 653310
rect 149890 653070 149980 653310
rect 150220 653070 150310 653310
rect 150550 653070 150660 653310
rect 150900 653070 150990 653310
rect 151230 653070 151320 653310
rect 151560 653070 151650 653310
rect 151890 653070 152000 653310
rect 152240 653070 152330 653310
rect 152570 653070 152660 653310
rect 152900 653070 152990 653310
rect 153230 653070 153340 653310
rect 153580 653070 153670 653310
rect 153910 653070 154000 653310
rect 154240 653070 154330 653310
rect 154570 653070 154680 653310
rect 154920 653070 155010 653310
rect 155250 653070 155340 653310
rect 155580 653070 155670 653310
rect 155910 653070 155960 653310
rect 110760 652980 155960 653070
rect 110760 652740 110810 652980
rect 111050 652740 111160 652980
rect 111400 652740 111490 652980
rect 111730 652740 111820 652980
rect 112060 652740 112150 652980
rect 112390 652740 112500 652980
rect 112740 652740 112830 652980
rect 113070 652740 113160 652980
rect 113400 652740 113490 652980
rect 113730 652740 113840 652980
rect 114080 652740 114170 652980
rect 114410 652740 114500 652980
rect 114740 652740 114830 652980
rect 115070 652740 115180 652980
rect 115420 652740 115510 652980
rect 115750 652740 115840 652980
rect 116080 652740 116170 652980
rect 116410 652740 116520 652980
rect 116760 652740 116850 652980
rect 117090 652740 117180 652980
rect 117420 652740 117510 652980
rect 117750 652740 117860 652980
rect 118100 652740 118190 652980
rect 118430 652740 118520 652980
rect 118760 652740 118850 652980
rect 119090 652740 119200 652980
rect 119440 652740 119530 652980
rect 119770 652740 119860 652980
rect 120100 652740 120190 652980
rect 120430 652740 120540 652980
rect 120780 652740 120870 652980
rect 121110 652740 121200 652980
rect 121440 652740 121530 652980
rect 121770 652740 122190 652980
rect 122430 652740 122540 652980
rect 122780 652740 122870 652980
rect 123110 652740 123200 652980
rect 123440 652740 123530 652980
rect 123770 652740 123880 652980
rect 124120 652740 124210 652980
rect 124450 652740 124540 652980
rect 124780 652740 124870 652980
rect 125110 652740 125220 652980
rect 125460 652740 125550 652980
rect 125790 652740 125880 652980
rect 126120 652740 126210 652980
rect 126450 652740 126560 652980
rect 126800 652740 126890 652980
rect 127130 652740 127220 652980
rect 127460 652740 127550 652980
rect 127790 652740 127900 652980
rect 128140 652740 128230 652980
rect 128470 652740 128560 652980
rect 128800 652740 128890 652980
rect 129130 652740 129240 652980
rect 129480 652740 129570 652980
rect 129810 652740 129900 652980
rect 130140 652740 130230 652980
rect 130470 652740 130580 652980
rect 130820 652740 130910 652980
rect 131150 652740 131240 652980
rect 131480 652740 131570 652980
rect 131810 652740 131920 652980
rect 132160 652740 132250 652980
rect 132490 652740 132580 652980
rect 132820 652740 132910 652980
rect 133150 652740 133570 652980
rect 133810 652740 133920 652980
rect 134160 652740 134250 652980
rect 134490 652740 134580 652980
rect 134820 652740 134910 652980
rect 135150 652740 135260 652980
rect 135500 652740 135590 652980
rect 135830 652740 135920 652980
rect 136160 652740 136250 652980
rect 136490 652740 136600 652980
rect 136840 652740 136930 652980
rect 137170 652740 137260 652980
rect 137500 652740 137590 652980
rect 137830 652740 137940 652980
rect 138180 652740 138270 652980
rect 138510 652740 138600 652980
rect 138840 652740 138930 652980
rect 139170 652740 139280 652980
rect 139520 652740 139610 652980
rect 139850 652740 139940 652980
rect 140180 652740 140270 652980
rect 140510 652740 140620 652980
rect 140860 652740 140950 652980
rect 141190 652740 141280 652980
rect 141520 652740 141610 652980
rect 141850 652740 141960 652980
rect 142200 652740 142290 652980
rect 142530 652740 142620 652980
rect 142860 652740 142950 652980
rect 143190 652740 143300 652980
rect 143540 652740 143630 652980
rect 143870 652740 143960 652980
rect 144200 652740 144290 652980
rect 144530 652740 144950 652980
rect 145190 652740 145300 652980
rect 145540 652740 145630 652980
rect 145870 652740 145960 652980
rect 146200 652740 146290 652980
rect 146530 652740 146640 652980
rect 146880 652740 146970 652980
rect 147210 652740 147300 652980
rect 147540 652740 147630 652980
rect 147870 652740 147980 652980
rect 148220 652740 148310 652980
rect 148550 652740 148640 652980
rect 148880 652740 148970 652980
rect 149210 652740 149320 652980
rect 149560 652740 149650 652980
rect 149890 652740 149980 652980
rect 150220 652740 150310 652980
rect 150550 652740 150660 652980
rect 150900 652740 150990 652980
rect 151230 652740 151320 652980
rect 151560 652740 151650 652980
rect 151890 652740 152000 652980
rect 152240 652740 152330 652980
rect 152570 652740 152660 652980
rect 152900 652740 152990 652980
rect 153230 652740 153340 652980
rect 153580 652740 153670 652980
rect 153910 652740 154000 652980
rect 154240 652740 154330 652980
rect 154570 652740 154680 652980
rect 154920 652740 155010 652980
rect 155250 652740 155340 652980
rect 155580 652740 155670 652980
rect 155910 652740 155960 652980
rect 110760 652650 155960 652740
rect 110760 652410 110810 652650
rect 111050 652410 111160 652650
rect 111400 652410 111490 652650
rect 111730 652410 111820 652650
rect 112060 652410 112150 652650
rect 112390 652410 112500 652650
rect 112740 652410 112830 652650
rect 113070 652410 113160 652650
rect 113400 652410 113490 652650
rect 113730 652410 113840 652650
rect 114080 652410 114170 652650
rect 114410 652410 114500 652650
rect 114740 652410 114830 652650
rect 115070 652410 115180 652650
rect 115420 652410 115510 652650
rect 115750 652410 115840 652650
rect 116080 652410 116170 652650
rect 116410 652410 116520 652650
rect 116760 652410 116850 652650
rect 117090 652410 117180 652650
rect 117420 652410 117510 652650
rect 117750 652410 117860 652650
rect 118100 652410 118190 652650
rect 118430 652410 118520 652650
rect 118760 652410 118850 652650
rect 119090 652410 119200 652650
rect 119440 652410 119530 652650
rect 119770 652410 119860 652650
rect 120100 652410 120190 652650
rect 120430 652410 120540 652650
rect 120780 652410 120870 652650
rect 121110 652410 121200 652650
rect 121440 652410 121530 652650
rect 121770 652410 122190 652650
rect 122430 652410 122540 652650
rect 122780 652410 122870 652650
rect 123110 652410 123200 652650
rect 123440 652410 123530 652650
rect 123770 652410 123880 652650
rect 124120 652410 124210 652650
rect 124450 652410 124540 652650
rect 124780 652410 124870 652650
rect 125110 652410 125220 652650
rect 125460 652410 125550 652650
rect 125790 652410 125880 652650
rect 126120 652410 126210 652650
rect 126450 652410 126560 652650
rect 126800 652410 126890 652650
rect 127130 652410 127220 652650
rect 127460 652410 127550 652650
rect 127790 652410 127900 652650
rect 128140 652410 128230 652650
rect 128470 652410 128560 652650
rect 128800 652410 128890 652650
rect 129130 652410 129240 652650
rect 129480 652410 129570 652650
rect 129810 652410 129900 652650
rect 130140 652410 130230 652650
rect 130470 652410 130580 652650
rect 130820 652410 130910 652650
rect 131150 652410 131240 652650
rect 131480 652410 131570 652650
rect 131810 652410 131920 652650
rect 132160 652410 132250 652650
rect 132490 652410 132580 652650
rect 132820 652410 132910 652650
rect 133150 652410 133570 652650
rect 133810 652410 133920 652650
rect 134160 652410 134250 652650
rect 134490 652410 134580 652650
rect 134820 652410 134910 652650
rect 135150 652410 135260 652650
rect 135500 652410 135590 652650
rect 135830 652410 135920 652650
rect 136160 652410 136250 652650
rect 136490 652410 136600 652650
rect 136840 652410 136930 652650
rect 137170 652410 137260 652650
rect 137500 652410 137590 652650
rect 137830 652410 137940 652650
rect 138180 652410 138270 652650
rect 138510 652410 138600 652650
rect 138840 652410 138930 652650
rect 139170 652410 139280 652650
rect 139520 652410 139610 652650
rect 139850 652410 139940 652650
rect 140180 652410 140270 652650
rect 140510 652410 140620 652650
rect 140860 652410 140950 652650
rect 141190 652410 141280 652650
rect 141520 652410 141610 652650
rect 141850 652410 141960 652650
rect 142200 652410 142290 652650
rect 142530 652410 142620 652650
rect 142860 652410 142950 652650
rect 143190 652410 143300 652650
rect 143540 652410 143630 652650
rect 143870 652410 143960 652650
rect 144200 652410 144290 652650
rect 144530 652410 144950 652650
rect 145190 652410 145300 652650
rect 145540 652410 145630 652650
rect 145870 652410 145960 652650
rect 146200 652410 146290 652650
rect 146530 652410 146640 652650
rect 146880 652410 146970 652650
rect 147210 652410 147300 652650
rect 147540 652410 147630 652650
rect 147870 652410 147980 652650
rect 148220 652410 148310 652650
rect 148550 652410 148640 652650
rect 148880 652410 148970 652650
rect 149210 652410 149320 652650
rect 149560 652410 149650 652650
rect 149890 652410 149980 652650
rect 150220 652410 150310 652650
rect 150550 652410 150660 652650
rect 150900 652410 150990 652650
rect 151230 652410 151320 652650
rect 151560 652410 151650 652650
rect 151890 652410 152000 652650
rect 152240 652410 152330 652650
rect 152570 652410 152660 652650
rect 152900 652410 152990 652650
rect 153230 652410 153340 652650
rect 153580 652410 153670 652650
rect 153910 652410 154000 652650
rect 154240 652410 154330 652650
rect 154570 652410 154680 652650
rect 154920 652410 155010 652650
rect 155250 652410 155340 652650
rect 155580 652410 155670 652650
rect 155910 652410 155960 652650
rect 110760 652300 155960 652410
rect 110760 652060 110810 652300
rect 111050 652060 111160 652300
rect 111400 652060 111490 652300
rect 111730 652060 111820 652300
rect 112060 652060 112150 652300
rect 112390 652060 112500 652300
rect 112740 652060 112830 652300
rect 113070 652060 113160 652300
rect 113400 652060 113490 652300
rect 113730 652060 113840 652300
rect 114080 652060 114170 652300
rect 114410 652060 114500 652300
rect 114740 652060 114830 652300
rect 115070 652060 115180 652300
rect 115420 652060 115510 652300
rect 115750 652060 115840 652300
rect 116080 652060 116170 652300
rect 116410 652060 116520 652300
rect 116760 652060 116850 652300
rect 117090 652060 117180 652300
rect 117420 652060 117510 652300
rect 117750 652060 117860 652300
rect 118100 652060 118190 652300
rect 118430 652060 118520 652300
rect 118760 652060 118850 652300
rect 119090 652060 119200 652300
rect 119440 652060 119530 652300
rect 119770 652060 119860 652300
rect 120100 652060 120190 652300
rect 120430 652060 120540 652300
rect 120780 652060 120870 652300
rect 121110 652060 121200 652300
rect 121440 652060 121530 652300
rect 121770 652060 122190 652300
rect 122430 652060 122540 652300
rect 122780 652060 122870 652300
rect 123110 652060 123200 652300
rect 123440 652060 123530 652300
rect 123770 652060 123880 652300
rect 124120 652060 124210 652300
rect 124450 652060 124540 652300
rect 124780 652060 124870 652300
rect 125110 652060 125220 652300
rect 125460 652060 125550 652300
rect 125790 652060 125880 652300
rect 126120 652060 126210 652300
rect 126450 652060 126560 652300
rect 126800 652060 126890 652300
rect 127130 652060 127220 652300
rect 127460 652060 127550 652300
rect 127790 652060 127900 652300
rect 128140 652060 128230 652300
rect 128470 652060 128560 652300
rect 128800 652060 128890 652300
rect 129130 652060 129240 652300
rect 129480 652060 129570 652300
rect 129810 652060 129900 652300
rect 130140 652060 130230 652300
rect 130470 652060 130580 652300
rect 130820 652060 130910 652300
rect 131150 652060 131240 652300
rect 131480 652060 131570 652300
rect 131810 652060 131920 652300
rect 132160 652060 132250 652300
rect 132490 652060 132580 652300
rect 132820 652060 132910 652300
rect 133150 652060 133570 652300
rect 133810 652060 133920 652300
rect 134160 652060 134250 652300
rect 134490 652060 134580 652300
rect 134820 652060 134910 652300
rect 135150 652060 135260 652300
rect 135500 652060 135590 652300
rect 135830 652060 135920 652300
rect 136160 652060 136250 652300
rect 136490 652060 136600 652300
rect 136840 652060 136930 652300
rect 137170 652060 137260 652300
rect 137500 652060 137590 652300
rect 137830 652060 137940 652300
rect 138180 652060 138270 652300
rect 138510 652060 138600 652300
rect 138840 652060 138930 652300
rect 139170 652060 139280 652300
rect 139520 652060 139610 652300
rect 139850 652060 139940 652300
rect 140180 652060 140270 652300
rect 140510 652060 140620 652300
rect 140860 652060 140950 652300
rect 141190 652060 141280 652300
rect 141520 652060 141610 652300
rect 141850 652060 141960 652300
rect 142200 652060 142290 652300
rect 142530 652060 142620 652300
rect 142860 652060 142950 652300
rect 143190 652060 143300 652300
rect 143540 652060 143630 652300
rect 143870 652060 143960 652300
rect 144200 652060 144290 652300
rect 144530 652060 144950 652300
rect 145190 652060 145300 652300
rect 145540 652060 145630 652300
rect 145870 652060 145960 652300
rect 146200 652060 146290 652300
rect 146530 652060 146640 652300
rect 146880 652060 146970 652300
rect 147210 652060 147300 652300
rect 147540 652060 147630 652300
rect 147870 652060 147980 652300
rect 148220 652060 148310 652300
rect 148550 652060 148640 652300
rect 148880 652060 148970 652300
rect 149210 652060 149320 652300
rect 149560 652060 149650 652300
rect 149890 652060 149980 652300
rect 150220 652060 150310 652300
rect 150550 652060 150660 652300
rect 150900 652060 150990 652300
rect 151230 652060 151320 652300
rect 151560 652060 151650 652300
rect 151890 652060 152000 652300
rect 152240 652060 152330 652300
rect 152570 652060 152660 652300
rect 152900 652060 152990 652300
rect 153230 652060 153340 652300
rect 153580 652060 153670 652300
rect 153910 652060 154000 652300
rect 154240 652060 154330 652300
rect 154570 652060 154680 652300
rect 154920 652060 155010 652300
rect 155250 652060 155340 652300
rect 155580 652060 155670 652300
rect 155910 652060 155960 652300
rect 110760 651970 155960 652060
rect 110760 651730 110810 651970
rect 111050 651730 111160 651970
rect 111400 651730 111490 651970
rect 111730 651730 111820 651970
rect 112060 651730 112150 651970
rect 112390 651730 112500 651970
rect 112740 651730 112830 651970
rect 113070 651730 113160 651970
rect 113400 651730 113490 651970
rect 113730 651730 113840 651970
rect 114080 651730 114170 651970
rect 114410 651730 114500 651970
rect 114740 651730 114830 651970
rect 115070 651730 115180 651970
rect 115420 651730 115510 651970
rect 115750 651730 115840 651970
rect 116080 651730 116170 651970
rect 116410 651730 116520 651970
rect 116760 651730 116850 651970
rect 117090 651730 117180 651970
rect 117420 651730 117510 651970
rect 117750 651730 117860 651970
rect 118100 651730 118190 651970
rect 118430 651730 118520 651970
rect 118760 651730 118850 651970
rect 119090 651730 119200 651970
rect 119440 651730 119530 651970
rect 119770 651730 119860 651970
rect 120100 651730 120190 651970
rect 120430 651730 120540 651970
rect 120780 651730 120870 651970
rect 121110 651730 121200 651970
rect 121440 651730 121530 651970
rect 121770 651730 122190 651970
rect 122430 651730 122540 651970
rect 122780 651730 122870 651970
rect 123110 651730 123200 651970
rect 123440 651730 123530 651970
rect 123770 651730 123880 651970
rect 124120 651730 124210 651970
rect 124450 651730 124540 651970
rect 124780 651730 124870 651970
rect 125110 651730 125220 651970
rect 125460 651730 125550 651970
rect 125790 651730 125880 651970
rect 126120 651730 126210 651970
rect 126450 651730 126560 651970
rect 126800 651730 126890 651970
rect 127130 651730 127220 651970
rect 127460 651730 127550 651970
rect 127790 651730 127900 651970
rect 128140 651730 128230 651970
rect 128470 651730 128560 651970
rect 128800 651730 128890 651970
rect 129130 651730 129240 651970
rect 129480 651730 129570 651970
rect 129810 651730 129900 651970
rect 130140 651730 130230 651970
rect 130470 651730 130580 651970
rect 130820 651730 130910 651970
rect 131150 651730 131240 651970
rect 131480 651730 131570 651970
rect 131810 651730 131920 651970
rect 132160 651730 132250 651970
rect 132490 651730 132580 651970
rect 132820 651730 132910 651970
rect 133150 651730 133570 651970
rect 133810 651730 133920 651970
rect 134160 651730 134250 651970
rect 134490 651730 134580 651970
rect 134820 651730 134910 651970
rect 135150 651730 135260 651970
rect 135500 651730 135590 651970
rect 135830 651730 135920 651970
rect 136160 651730 136250 651970
rect 136490 651730 136600 651970
rect 136840 651730 136930 651970
rect 137170 651730 137260 651970
rect 137500 651730 137590 651970
rect 137830 651730 137940 651970
rect 138180 651730 138270 651970
rect 138510 651730 138600 651970
rect 138840 651730 138930 651970
rect 139170 651730 139280 651970
rect 139520 651730 139610 651970
rect 139850 651730 139940 651970
rect 140180 651730 140270 651970
rect 140510 651730 140620 651970
rect 140860 651730 140950 651970
rect 141190 651730 141280 651970
rect 141520 651730 141610 651970
rect 141850 651730 141960 651970
rect 142200 651730 142290 651970
rect 142530 651730 142620 651970
rect 142860 651730 142950 651970
rect 143190 651730 143300 651970
rect 143540 651730 143630 651970
rect 143870 651730 143960 651970
rect 144200 651730 144290 651970
rect 144530 651730 144950 651970
rect 145190 651730 145300 651970
rect 145540 651730 145630 651970
rect 145870 651730 145960 651970
rect 146200 651730 146290 651970
rect 146530 651730 146640 651970
rect 146880 651730 146970 651970
rect 147210 651730 147300 651970
rect 147540 651730 147630 651970
rect 147870 651730 147980 651970
rect 148220 651730 148310 651970
rect 148550 651730 148640 651970
rect 148880 651730 148970 651970
rect 149210 651730 149320 651970
rect 149560 651730 149650 651970
rect 149890 651730 149980 651970
rect 150220 651730 150310 651970
rect 150550 651730 150660 651970
rect 150900 651730 150990 651970
rect 151230 651730 151320 651970
rect 151560 651730 151650 651970
rect 151890 651730 152000 651970
rect 152240 651730 152330 651970
rect 152570 651730 152660 651970
rect 152900 651730 152990 651970
rect 153230 651730 153340 651970
rect 153580 651730 153670 651970
rect 153910 651730 154000 651970
rect 154240 651730 154330 651970
rect 154570 651730 154680 651970
rect 154920 651730 155010 651970
rect 155250 651730 155340 651970
rect 155580 651730 155670 651970
rect 155910 651730 155960 651970
rect 110760 651640 155960 651730
rect 110760 651400 110810 651640
rect 111050 651400 111160 651640
rect 111400 651400 111490 651640
rect 111730 651400 111820 651640
rect 112060 651400 112150 651640
rect 112390 651400 112500 651640
rect 112740 651400 112830 651640
rect 113070 651400 113160 651640
rect 113400 651400 113490 651640
rect 113730 651400 113840 651640
rect 114080 651400 114170 651640
rect 114410 651400 114500 651640
rect 114740 651400 114830 651640
rect 115070 651400 115180 651640
rect 115420 651400 115510 651640
rect 115750 651400 115840 651640
rect 116080 651400 116170 651640
rect 116410 651400 116520 651640
rect 116760 651400 116850 651640
rect 117090 651400 117180 651640
rect 117420 651400 117510 651640
rect 117750 651400 117860 651640
rect 118100 651400 118190 651640
rect 118430 651400 118520 651640
rect 118760 651400 118850 651640
rect 119090 651400 119200 651640
rect 119440 651400 119530 651640
rect 119770 651400 119860 651640
rect 120100 651400 120190 651640
rect 120430 651400 120540 651640
rect 120780 651400 120870 651640
rect 121110 651400 121200 651640
rect 121440 651400 121530 651640
rect 121770 651400 122190 651640
rect 122430 651400 122540 651640
rect 122780 651400 122870 651640
rect 123110 651400 123200 651640
rect 123440 651400 123530 651640
rect 123770 651400 123880 651640
rect 124120 651400 124210 651640
rect 124450 651400 124540 651640
rect 124780 651400 124870 651640
rect 125110 651400 125220 651640
rect 125460 651400 125550 651640
rect 125790 651400 125880 651640
rect 126120 651400 126210 651640
rect 126450 651400 126560 651640
rect 126800 651400 126890 651640
rect 127130 651400 127220 651640
rect 127460 651400 127550 651640
rect 127790 651400 127900 651640
rect 128140 651400 128230 651640
rect 128470 651400 128560 651640
rect 128800 651400 128890 651640
rect 129130 651400 129240 651640
rect 129480 651400 129570 651640
rect 129810 651400 129900 651640
rect 130140 651400 130230 651640
rect 130470 651400 130580 651640
rect 130820 651400 130910 651640
rect 131150 651400 131240 651640
rect 131480 651400 131570 651640
rect 131810 651400 131920 651640
rect 132160 651400 132250 651640
rect 132490 651400 132580 651640
rect 132820 651400 132910 651640
rect 133150 651400 133570 651640
rect 133810 651400 133920 651640
rect 134160 651400 134250 651640
rect 134490 651400 134580 651640
rect 134820 651400 134910 651640
rect 135150 651400 135260 651640
rect 135500 651400 135590 651640
rect 135830 651400 135920 651640
rect 136160 651400 136250 651640
rect 136490 651400 136600 651640
rect 136840 651400 136930 651640
rect 137170 651400 137260 651640
rect 137500 651400 137590 651640
rect 137830 651400 137940 651640
rect 138180 651400 138270 651640
rect 138510 651400 138600 651640
rect 138840 651400 138930 651640
rect 139170 651400 139280 651640
rect 139520 651400 139610 651640
rect 139850 651400 139940 651640
rect 140180 651400 140270 651640
rect 140510 651400 140620 651640
rect 140860 651400 140950 651640
rect 141190 651400 141280 651640
rect 141520 651400 141610 651640
rect 141850 651400 141960 651640
rect 142200 651400 142290 651640
rect 142530 651400 142620 651640
rect 142860 651400 142950 651640
rect 143190 651400 143300 651640
rect 143540 651400 143630 651640
rect 143870 651400 143960 651640
rect 144200 651400 144290 651640
rect 144530 651400 144950 651640
rect 145190 651400 145300 651640
rect 145540 651400 145630 651640
rect 145870 651400 145960 651640
rect 146200 651400 146290 651640
rect 146530 651400 146640 651640
rect 146880 651400 146970 651640
rect 147210 651400 147300 651640
rect 147540 651400 147630 651640
rect 147870 651400 147980 651640
rect 148220 651400 148310 651640
rect 148550 651400 148640 651640
rect 148880 651400 148970 651640
rect 149210 651400 149320 651640
rect 149560 651400 149650 651640
rect 149890 651400 149980 651640
rect 150220 651400 150310 651640
rect 150550 651400 150660 651640
rect 150900 651400 150990 651640
rect 151230 651400 151320 651640
rect 151560 651400 151650 651640
rect 151890 651400 152000 651640
rect 152240 651400 152330 651640
rect 152570 651400 152660 651640
rect 152900 651400 152990 651640
rect 153230 651400 153340 651640
rect 153580 651400 153670 651640
rect 153910 651400 154000 651640
rect 154240 651400 154330 651640
rect 154570 651400 154680 651640
rect 154920 651400 155010 651640
rect 155250 651400 155340 651640
rect 155580 651400 155670 651640
rect 155910 651400 155960 651640
rect 110760 651310 155960 651400
rect 110760 651070 110810 651310
rect 111050 651070 111160 651310
rect 111400 651070 111490 651310
rect 111730 651070 111820 651310
rect 112060 651070 112150 651310
rect 112390 651070 112500 651310
rect 112740 651070 112830 651310
rect 113070 651070 113160 651310
rect 113400 651070 113490 651310
rect 113730 651070 113840 651310
rect 114080 651070 114170 651310
rect 114410 651070 114500 651310
rect 114740 651070 114830 651310
rect 115070 651070 115180 651310
rect 115420 651070 115510 651310
rect 115750 651070 115840 651310
rect 116080 651070 116170 651310
rect 116410 651070 116520 651310
rect 116760 651070 116850 651310
rect 117090 651070 117180 651310
rect 117420 651070 117510 651310
rect 117750 651070 117860 651310
rect 118100 651070 118190 651310
rect 118430 651070 118520 651310
rect 118760 651070 118850 651310
rect 119090 651070 119200 651310
rect 119440 651070 119530 651310
rect 119770 651070 119860 651310
rect 120100 651070 120190 651310
rect 120430 651070 120540 651310
rect 120780 651070 120870 651310
rect 121110 651070 121200 651310
rect 121440 651070 121530 651310
rect 121770 651070 122190 651310
rect 122430 651070 122540 651310
rect 122780 651070 122870 651310
rect 123110 651070 123200 651310
rect 123440 651070 123530 651310
rect 123770 651070 123880 651310
rect 124120 651070 124210 651310
rect 124450 651070 124540 651310
rect 124780 651070 124870 651310
rect 125110 651070 125220 651310
rect 125460 651070 125550 651310
rect 125790 651070 125880 651310
rect 126120 651070 126210 651310
rect 126450 651070 126560 651310
rect 126800 651070 126890 651310
rect 127130 651070 127220 651310
rect 127460 651070 127550 651310
rect 127790 651070 127900 651310
rect 128140 651070 128230 651310
rect 128470 651070 128560 651310
rect 128800 651070 128890 651310
rect 129130 651070 129240 651310
rect 129480 651070 129570 651310
rect 129810 651070 129900 651310
rect 130140 651070 130230 651310
rect 130470 651070 130580 651310
rect 130820 651070 130910 651310
rect 131150 651070 131240 651310
rect 131480 651070 131570 651310
rect 131810 651070 131920 651310
rect 132160 651070 132250 651310
rect 132490 651070 132580 651310
rect 132820 651070 132910 651310
rect 133150 651070 133570 651310
rect 133810 651070 133920 651310
rect 134160 651070 134250 651310
rect 134490 651070 134580 651310
rect 134820 651070 134910 651310
rect 135150 651070 135260 651310
rect 135500 651070 135590 651310
rect 135830 651070 135920 651310
rect 136160 651070 136250 651310
rect 136490 651070 136600 651310
rect 136840 651070 136930 651310
rect 137170 651070 137260 651310
rect 137500 651070 137590 651310
rect 137830 651070 137940 651310
rect 138180 651070 138270 651310
rect 138510 651070 138600 651310
rect 138840 651070 138930 651310
rect 139170 651070 139280 651310
rect 139520 651070 139610 651310
rect 139850 651070 139940 651310
rect 140180 651070 140270 651310
rect 140510 651070 140620 651310
rect 140860 651070 140950 651310
rect 141190 651070 141280 651310
rect 141520 651070 141610 651310
rect 141850 651070 141960 651310
rect 142200 651070 142290 651310
rect 142530 651070 142620 651310
rect 142860 651070 142950 651310
rect 143190 651070 143300 651310
rect 143540 651070 143630 651310
rect 143870 651070 143960 651310
rect 144200 651070 144290 651310
rect 144530 651070 144950 651310
rect 145190 651070 145300 651310
rect 145540 651070 145630 651310
rect 145870 651070 145960 651310
rect 146200 651070 146290 651310
rect 146530 651070 146640 651310
rect 146880 651070 146970 651310
rect 147210 651070 147300 651310
rect 147540 651070 147630 651310
rect 147870 651070 147980 651310
rect 148220 651070 148310 651310
rect 148550 651070 148640 651310
rect 148880 651070 148970 651310
rect 149210 651070 149320 651310
rect 149560 651070 149650 651310
rect 149890 651070 149980 651310
rect 150220 651070 150310 651310
rect 150550 651070 150660 651310
rect 150900 651070 150990 651310
rect 151230 651070 151320 651310
rect 151560 651070 151650 651310
rect 151890 651070 152000 651310
rect 152240 651070 152330 651310
rect 152570 651070 152660 651310
rect 152900 651070 152990 651310
rect 153230 651070 153340 651310
rect 153580 651070 153670 651310
rect 153910 651070 154000 651310
rect 154240 651070 154330 651310
rect 154570 651070 154680 651310
rect 154920 651070 155010 651310
rect 155250 651070 155340 651310
rect 155580 651070 155670 651310
rect 155910 651070 155960 651310
rect 110760 650960 155960 651070
rect 110760 650720 110810 650960
rect 111050 650720 111160 650960
rect 111400 650720 111490 650960
rect 111730 650720 111820 650960
rect 112060 650720 112150 650960
rect 112390 650720 112500 650960
rect 112740 650720 112830 650960
rect 113070 650720 113160 650960
rect 113400 650720 113490 650960
rect 113730 650720 113840 650960
rect 114080 650720 114170 650960
rect 114410 650720 114500 650960
rect 114740 650720 114830 650960
rect 115070 650720 115180 650960
rect 115420 650720 115510 650960
rect 115750 650720 115840 650960
rect 116080 650720 116170 650960
rect 116410 650720 116520 650960
rect 116760 650720 116850 650960
rect 117090 650720 117180 650960
rect 117420 650720 117510 650960
rect 117750 650720 117860 650960
rect 118100 650720 118190 650960
rect 118430 650720 118520 650960
rect 118760 650720 118850 650960
rect 119090 650720 119200 650960
rect 119440 650720 119530 650960
rect 119770 650720 119860 650960
rect 120100 650720 120190 650960
rect 120430 650720 120540 650960
rect 120780 650720 120870 650960
rect 121110 650720 121200 650960
rect 121440 650720 121530 650960
rect 121770 650720 122190 650960
rect 122430 650720 122540 650960
rect 122780 650720 122870 650960
rect 123110 650720 123200 650960
rect 123440 650720 123530 650960
rect 123770 650720 123880 650960
rect 124120 650720 124210 650960
rect 124450 650720 124540 650960
rect 124780 650720 124870 650960
rect 125110 650720 125220 650960
rect 125460 650720 125550 650960
rect 125790 650720 125880 650960
rect 126120 650720 126210 650960
rect 126450 650720 126560 650960
rect 126800 650720 126890 650960
rect 127130 650720 127220 650960
rect 127460 650720 127550 650960
rect 127790 650720 127900 650960
rect 128140 650720 128230 650960
rect 128470 650720 128560 650960
rect 128800 650720 128890 650960
rect 129130 650720 129240 650960
rect 129480 650720 129570 650960
rect 129810 650720 129900 650960
rect 130140 650720 130230 650960
rect 130470 650720 130580 650960
rect 130820 650720 130910 650960
rect 131150 650720 131240 650960
rect 131480 650720 131570 650960
rect 131810 650720 131920 650960
rect 132160 650720 132250 650960
rect 132490 650720 132580 650960
rect 132820 650720 132910 650960
rect 133150 650720 133570 650960
rect 133810 650720 133920 650960
rect 134160 650720 134250 650960
rect 134490 650720 134580 650960
rect 134820 650720 134910 650960
rect 135150 650720 135260 650960
rect 135500 650720 135590 650960
rect 135830 650720 135920 650960
rect 136160 650720 136250 650960
rect 136490 650720 136600 650960
rect 136840 650720 136930 650960
rect 137170 650720 137260 650960
rect 137500 650720 137590 650960
rect 137830 650720 137940 650960
rect 138180 650720 138270 650960
rect 138510 650720 138600 650960
rect 138840 650720 138930 650960
rect 139170 650720 139280 650960
rect 139520 650720 139610 650960
rect 139850 650720 139940 650960
rect 140180 650720 140270 650960
rect 140510 650720 140620 650960
rect 140860 650720 140950 650960
rect 141190 650720 141280 650960
rect 141520 650720 141610 650960
rect 141850 650720 141960 650960
rect 142200 650720 142290 650960
rect 142530 650720 142620 650960
rect 142860 650720 142950 650960
rect 143190 650720 143300 650960
rect 143540 650720 143630 650960
rect 143870 650720 143960 650960
rect 144200 650720 144290 650960
rect 144530 650720 144950 650960
rect 145190 650720 145300 650960
rect 145540 650720 145630 650960
rect 145870 650720 145960 650960
rect 146200 650720 146290 650960
rect 146530 650720 146640 650960
rect 146880 650720 146970 650960
rect 147210 650720 147300 650960
rect 147540 650720 147630 650960
rect 147870 650720 147980 650960
rect 148220 650720 148310 650960
rect 148550 650720 148640 650960
rect 148880 650720 148970 650960
rect 149210 650720 149320 650960
rect 149560 650720 149650 650960
rect 149890 650720 149980 650960
rect 150220 650720 150310 650960
rect 150550 650720 150660 650960
rect 150900 650720 150990 650960
rect 151230 650720 151320 650960
rect 151560 650720 151650 650960
rect 151890 650720 152000 650960
rect 152240 650720 152330 650960
rect 152570 650720 152660 650960
rect 152900 650720 152990 650960
rect 153230 650720 153340 650960
rect 153580 650720 153670 650960
rect 153910 650720 154000 650960
rect 154240 650720 154330 650960
rect 154570 650720 154680 650960
rect 154920 650720 155010 650960
rect 155250 650720 155340 650960
rect 155580 650720 155670 650960
rect 155910 650720 155960 650960
rect 110760 650630 155960 650720
rect 110760 650390 110810 650630
rect 111050 650390 111160 650630
rect 111400 650390 111490 650630
rect 111730 650390 111820 650630
rect 112060 650390 112150 650630
rect 112390 650390 112500 650630
rect 112740 650390 112830 650630
rect 113070 650390 113160 650630
rect 113400 650390 113490 650630
rect 113730 650390 113840 650630
rect 114080 650390 114170 650630
rect 114410 650390 114500 650630
rect 114740 650390 114830 650630
rect 115070 650390 115180 650630
rect 115420 650390 115510 650630
rect 115750 650390 115840 650630
rect 116080 650390 116170 650630
rect 116410 650390 116520 650630
rect 116760 650390 116850 650630
rect 117090 650390 117180 650630
rect 117420 650390 117510 650630
rect 117750 650390 117860 650630
rect 118100 650390 118190 650630
rect 118430 650390 118520 650630
rect 118760 650390 118850 650630
rect 119090 650390 119200 650630
rect 119440 650390 119530 650630
rect 119770 650390 119860 650630
rect 120100 650390 120190 650630
rect 120430 650390 120540 650630
rect 120780 650390 120870 650630
rect 121110 650390 121200 650630
rect 121440 650390 121530 650630
rect 121770 650390 122190 650630
rect 122430 650390 122540 650630
rect 122780 650390 122870 650630
rect 123110 650390 123200 650630
rect 123440 650390 123530 650630
rect 123770 650390 123880 650630
rect 124120 650390 124210 650630
rect 124450 650390 124540 650630
rect 124780 650390 124870 650630
rect 125110 650390 125220 650630
rect 125460 650390 125550 650630
rect 125790 650390 125880 650630
rect 126120 650390 126210 650630
rect 126450 650390 126560 650630
rect 126800 650390 126890 650630
rect 127130 650390 127220 650630
rect 127460 650390 127550 650630
rect 127790 650390 127900 650630
rect 128140 650390 128230 650630
rect 128470 650390 128560 650630
rect 128800 650390 128890 650630
rect 129130 650390 129240 650630
rect 129480 650390 129570 650630
rect 129810 650390 129900 650630
rect 130140 650390 130230 650630
rect 130470 650390 130580 650630
rect 130820 650390 130910 650630
rect 131150 650390 131240 650630
rect 131480 650390 131570 650630
rect 131810 650390 131920 650630
rect 132160 650390 132250 650630
rect 132490 650390 132580 650630
rect 132820 650390 132910 650630
rect 133150 650390 133570 650630
rect 133810 650390 133920 650630
rect 134160 650390 134250 650630
rect 134490 650390 134580 650630
rect 134820 650390 134910 650630
rect 135150 650390 135260 650630
rect 135500 650390 135590 650630
rect 135830 650390 135920 650630
rect 136160 650390 136250 650630
rect 136490 650390 136600 650630
rect 136840 650390 136930 650630
rect 137170 650390 137260 650630
rect 137500 650390 137590 650630
rect 137830 650390 137940 650630
rect 138180 650390 138270 650630
rect 138510 650390 138600 650630
rect 138840 650390 138930 650630
rect 139170 650390 139280 650630
rect 139520 650390 139610 650630
rect 139850 650390 139940 650630
rect 140180 650390 140270 650630
rect 140510 650390 140620 650630
rect 140860 650390 140950 650630
rect 141190 650390 141280 650630
rect 141520 650390 141610 650630
rect 141850 650390 141960 650630
rect 142200 650390 142290 650630
rect 142530 650390 142620 650630
rect 142860 650390 142950 650630
rect 143190 650390 143300 650630
rect 143540 650390 143630 650630
rect 143870 650390 143960 650630
rect 144200 650390 144290 650630
rect 144530 650390 144950 650630
rect 145190 650390 145300 650630
rect 145540 650390 145630 650630
rect 145870 650390 145960 650630
rect 146200 650390 146290 650630
rect 146530 650390 146640 650630
rect 146880 650390 146970 650630
rect 147210 650390 147300 650630
rect 147540 650390 147630 650630
rect 147870 650390 147980 650630
rect 148220 650390 148310 650630
rect 148550 650390 148640 650630
rect 148880 650390 148970 650630
rect 149210 650390 149320 650630
rect 149560 650390 149650 650630
rect 149890 650390 149980 650630
rect 150220 650390 150310 650630
rect 150550 650390 150660 650630
rect 150900 650390 150990 650630
rect 151230 650390 151320 650630
rect 151560 650390 151650 650630
rect 151890 650390 152000 650630
rect 152240 650390 152330 650630
rect 152570 650390 152660 650630
rect 152900 650390 152990 650630
rect 153230 650390 153340 650630
rect 153580 650390 153670 650630
rect 153910 650390 154000 650630
rect 154240 650390 154330 650630
rect 154570 650390 154680 650630
rect 154920 650390 155010 650630
rect 155250 650390 155340 650630
rect 155580 650390 155670 650630
rect 155910 650390 155960 650630
rect 110760 650300 155960 650390
rect 110760 650060 110810 650300
rect 111050 650060 111160 650300
rect 111400 650060 111490 650300
rect 111730 650060 111820 650300
rect 112060 650060 112150 650300
rect 112390 650060 112500 650300
rect 112740 650060 112830 650300
rect 113070 650060 113160 650300
rect 113400 650060 113490 650300
rect 113730 650060 113840 650300
rect 114080 650060 114170 650300
rect 114410 650060 114500 650300
rect 114740 650060 114830 650300
rect 115070 650060 115180 650300
rect 115420 650060 115510 650300
rect 115750 650060 115840 650300
rect 116080 650060 116170 650300
rect 116410 650060 116520 650300
rect 116760 650060 116850 650300
rect 117090 650060 117180 650300
rect 117420 650060 117510 650300
rect 117750 650060 117860 650300
rect 118100 650060 118190 650300
rect 118430 650060 118520 650300
rect 118760 650060 118850 650300
rect 119090 650060 119200 650300
rect 119440 650060 119530 650300
rect 119770 650060 119860 650300
rect 120100 650060 120190 650300
rect 120430 650060 120540 650300
rect 120780 650060 120870 650300
rect 121110 650060 121200 650300
rect 121440 650060 121530 650300
rect 121770 650060 122190 650300
rect 122430 650060 122540 650300
rect 122780 650060 122870 650300
rect 123110 650060 123200 650300
rect 123440 650060 123530 650300
rect 123770 650060 123880 650300
rect 124120 650060 124210 650300
rect 124450 650060 124540 650300
rect 124780 650060 124870 650300
rect 125110 650060 125220 650300
rect 125460 650060 125550 650300
rect 125790 650060 125880 650300
rect 126120 650060 126210 650300
rect 126450 650060 126560 650300
rect 126800 650060 126890 650300
rect 127130 650060 127220 650300
rect 127460 650060 127550 650300
rect 127790 650060 127900 650300
rect 128140 650060 128230 650300
rect 128470 650060 128560 650300
rect 128800 650060 128890 650300
rect 129130 650060 129240 650300
rect 129480 650060 129570 650300
rect 129810 650060 129900 650300
rect 130140 650060 130230 650300
rect 130470 650060 130580 650300
rect 130820 650060 130910 650300
rect 131150 650060 131240 650300
rect 131480 650060 131570 650300
rect 131810 650060 131920 650300
rect 132160 650060 132250 650300
rect 132490 650060 132580 650300
rect 132820 650060 132910 650300
rect 133150 650060 133570 650300
rect 133810 650060 133920 650300
rect 134160 650060 134250 650300
rect 134490 650060 134580 650300
rect 134820 650060 134910 650300
rect 135150 650060 135260 650300
rect 135500 650060 135590 650300
rect 135830 650060 135920 650300
rect 136160 650060 136250 650300
rect 136490 650060 136600 650300
rect 136840 650060 136930 650300
rect 137170 650060 137260 650300
rect 137500 650060 137590 650300
rect 137830 650060 137940 650300
rect 138180 650060 138270 650300
rect 138510 650060 138600 650300
rect 138840 650060 138930 650300
rect 139170 650060 139280 650300
rect 139520 650060 139610 650300
rect 139850 650060 139940 650300
rect 140180 650060 140270 650300
rect 140510 650060 140620 650300
rect 140860 650060 140950 650300
rect 141190 650060 141280 650300
rect 141520 650060 141610 650300
rect 141850 650060 141960 650300
rect 142200 650060 142290 650300
rect 142530 650060 142620 650300
rect 142860 650060 142950 650300
rect 143190 650060 143300 650300
rect 143540 650060 143630 650300
rect 143870 650060 143960 650300
rect 144200 650060 144290 650300
rect 144530 650060 144950 650300
rect 145190 650060 145300 650300
rect 145540 650060 145630 650300
rect 145870 650060 145960 650300
rect 146200 650060 146290 650300
rect 146530 650060 146640 650300
rect 146880 650060 146970 650300
rect 147210 650060 147300 650300
rect 147540 650060 147630 650300
rect 147870 650060 147980 650300
rect 148220 650060 148310 650300
rect 148550 650060 148640 650300
rect 148880 650060 148970 650300
rect 149210 650060 149320 650300
rect 149560 650060 149650 650300
rect 149890 650060 149980 650300
rect 150220 650060 150310 650300
rect 150550 650060 150660 650300
rect 150900 650060 150990 650300
rect 151230 650060 151320 650300
rect 151560 650060 151650 650300
rect 151890 650060 152000 650300
rect 152240 650060 152330 650300
rect 152570 650060 152660 650300
rect 152900 650060 152990 650300
rect 153230 650060 153340 650300
rect 153580 650060 153670 650300
rect 153910 650060 154000 650300
rect 154240 650060 154330 650300
rect 154570 650060 154680 650300
rect 154920 650060 155010 650300
rect 155250 650060 155340 650300
rect 155580 650060 155670 650300
rect 155910 650060 155960 650300
rect 110760 649970 155960 650060
rect 110760 649730 110810 649970
rect 111050 649730 111160 649970
rect 111400 649730 111490 649970
rect 111730 649730 111820 649970
rect 112060 649730 112150 649970
rect 112390 649730 112500 649970
rect 112740 649730 112830 649970
rect 113070 649730 113160 649970
rect 113400 649730 113490 649970
rect 113730 649730 113840 649970
rect 114080 649730 114170 649970
rect 114410 649730 114500 649970
rect 114740 649730 114830 649970
rect 115070 649730 115180 649970
rect 115420 649730 115510 649970
rect 115750 649730 115840 649970
rect 116080 649730 116170 649970
rect 116410 649730 116520 649970
rect 116760 649730 116850 649970
rect 117090 649730 117180 649970
rect 117420 649730 117510 649970
rect 117750 649730 117860 649970
rect 118100 649730 118190 649970
rect 118430 649730 118520 649970
rect 118760 649730 118850 649970
rect 119090 649730 119200 649970
rect 119440 649730 119530 649970
rect 119770 649730 119860 649970
rect 120100 649730 120190 649970
rect 120430 649730 120540 649970
rect 120780 649730 120870 649970
rect 121110 649730 121200 649970
rect 121440 649730 121530 649970
rect 121770 649730 122190 649970
rect 122430 649730 122540 649970
rect 122780 649730 122870 649970
rect 123110 649730 123200 649970
rect 123440 649730 123530 649970
rect 123770 649730 123880 649970
rect 124120 649730 124210 649970
rect 124450 649730 124540 649970
rect 124780 649730 124870 649970
rect 125110 649730 125220 649970
rect 125460 649730 125550 649970
rect 125790 649730 125880 649970
rect 126120 649730 126210 649970
rect 126450 649730 126560 649970
rect 126800 649730 126890 649970
rect 127130 649730 127220 649970
rect 127460 649730 127550 649970
rect 127790 649730 127900 649970
rect 128140 649730 128230 649970
rect 128470 649730 128560 649970
rect 128800 649730 128890 649970
rect 129130 649730 129240 649970
rect 129480 649730 129570 649970
rect 129810 649730 129900 649970
rect 130140 649730 130230 649970
rect 130470 649730 130580 649970
rect 130820 649730 130910 649970
rect 131150 649730 131240 649970
rect 131480 649730 131570 649970
rect 131810 649730 131920 649970
rect 132160 649730 132250 649970
rect 132490 649730 132580 649970
rect 132820 649730 132910 649970
rect 133150 649730 133570 649970
rect 133810 649730 133920 649970
rect 134160 649730 134250 649970
rect 134490 649730 134580 649970
rect 134820 649730 134910 649970
rect 135150 649730 135260 649970
rect 135500 649730 135590 649970
rect 135830 649730 135920 649970
rect 136160 649730 136250 649970
rect 136490 649730 136600 649970
rect 136840 649730 136930 649970
rect 137170 649730 137260 649970
rect 137500 649730 137590 649970
rect 137830 649730 137940 649970
rect 138180 649730 138270 649970
rect 138510 649730 138600 649970
rect 138840 649730 138930 649970
rect 139170 649730 139280 649970
rect 139520 649730 139610 649970
rect 139850 649730 139940 649970
rect 140180 649730 140270 649970
rect 140510 649730 140620 649970
rect 140860 649730 140950 649970
rect 141190 649730 141280 649970
rect 141520 649730 141610 649970
rect 141850 649730 141960 649970
rect 142200 649730 142290 649970
rect 142530 649730 142620 649970
rect 142860 649730 142950 649970
rect 143190 649730 143300 649970
rect 143540 649730 143630 649970
rect 143870 649730 143960 649970
rect 144200 649730 144290 649970
rect 144530 649730 144950 649970
rect 145190 649730 145300 649970
rect 145540 649730 145630 649970
rect 145870 649730 145960 649970
rect 146200 649730 146290 649970
rect 146530 649730 146640 649970
rect 146880 649730 146970 649970
rect 147210 649730 147300 649970
rect 147540 649730 147630 649970
rect 147870 649730 147980 649970
rect 148220 649730 148310 649970
rect 148550 649730 148640 649970
rect 148880 649730 148970 649970
rect 149210 649730 149320 649970
rect 149560 649730 149650 649970
rect 149890 649730 149980 649970
rect 150220 649730 150310 649970
rect 150550 649730 150660 649970
rect 150900 649730 150990 649970
rect 151230 649730 151320 649970
rect 151560 649730 151650 649970
rect 151890 649730 152000 649970
rect 152240 649730 152330 649970
rect 152570 649730 152660 649970
rect 152900 649730 152990 649970
rect 153230 649730 153340 649970
rect 153580 649730 153670 649970
rect 153910 649730 154000 649970
rect 154240 649730 154330 649970
rect 154570 649730 154680 649970
rect 154920 649730 155010 649970
rect 155250 649730 155340 649970
rect 155580 649730 155670 649970
rect 155910 649730 155960 649970
rect 110760 649620 155960 649730
rect 110760 649380 110810 649620
rect 111050 649380 111160 649620
rect 111400 649380 111490 649620
rect 111730 649380 111820 649620
rect 112060 649380 112150 649620
rect 112390 649380 112500 649620
rect 112740 649380 112830 649620
rect 113070 649380 113160 649620
rect 113400 649380 113490 649620
rect 113730 649380 113840 649620
rect 114080 649380 114170 649620
rect 114410 649380 114500 649620
rect 114740 649380 114830 649620
rect 115070 649380 115180 649620
rect 115420 649380 115510 649620
rect 115750 649380 115840 649620
rect 116080 649380 116170 649620
rect 116410 649380 116520 649620
rect 116760 649380 116850 649620
rect 117090 649380 117180 649620
rect 117420 649380 117510 649620
rect 117750 649380 117860 649620
rect 118100 649380 118190 649620
rect 118430 649380 118520 649620
rect 118760 649380 118850 649620
rect 119090 649380 119200 649620
rect 119440 649380 119530 649620
rect 119770 649380 119860 649620
rect 120100 649380 120190 649620
rect 120430 649380 120540 649620
rect 120780 649380 120870 649620
rect 121110 649380 121200 649620
rect 121440 649380 121530 649620
rect 121770 649380 122190 649620
rect 122430 649380 122540 649620
rect 122780 649380 122870 649620
rect 123110 649380 123200 649620
rect 123440 649380 123530 649620
rect 123770 649380 123880 649620
rect 124120 649380 124210 649620
rect 124450 649380 124540 649620
rect 124780 649380 124870 649620
rect 125110 649380 125220 649620
rect 125460 649380 125550 649620
rect 125790 649380 125880 649620
rect 126120 649380 126210 649620
rect 126450 649380 126560 649620
rect 126800 649380 126890 649620
rect 127130 649380 127220 649620
rect 127460 649380 127550 649620
rect 127790 649380 127900 649620
rect 128140 649380 128230 649620
rect 128470 649380 128560 649620
rect 128800 649380 128890 649620
rect 129130 649380 129240 649620
rect 129480 649380 129570 649620
rect 129810 649380 129900 649620
rect 130140 649380 130230 649620
rect 130470 649380 130580 649620
rect 130820 649380 130910 649620
rect 131150 649380 131240 649620
rect 131480 649380 131570 649620
rect 131810 649380 131920 649620
rect 132160 649380 132250 649620
rect 132490 649380 132580 649620
rect 132820 649380 132910 649620
rect 133150 649380 133570 649620
rect 133810 649380 133920 649620
rect 134160 649380 134250 649620
rect 134490 649380 134580 649620
rect 134820 649380 134910 649620
rect 135150 649380 135260 649620
rect 135500 649380 135590 649620
rect 135830 649380 135920 649620
rect 136160 649380 136250 649620
rect 136490 649380 136600 649620
rect 136840 649380 136930 649620
rect 137170 649380 137260 649620
rect 137500 649380 137590 649620
rect 137830 649380 137940 649620
rect 138180 649380 138270 649620
rect 138510 649380 138600 649620
rect 138840 649380 138930 649620
rect 139170 649380 139280 649620
rect 139520 649380 139610 649620
rect 139850 649380 139940 649620
rect 140180 649380 140270 649620
rect 140510 649380 140620 649620
rect 140860 649380 140950 649620
rect 141190 649380 141280 649620
rect 141520 649380 141610 649620
rect 141850 649380 141960 649620
rect 142200 649380 142290 649620
rect 142530 649380 142620 649620
rect 142860 649380 142950 649620
rect 143190 649380 143300 649620
rect 143540 649380 143630 649620
rect 143870 649380 143960 649620
rect 144200 649380 144290 649620
rect 144530 649380 144950 649620
rect 145190 649380 145300 649620
rect 145540 649380 145630 649620
rect 145870 649380 145960 649620
rect 146200 649380 146290 649620
rect 146530 649380 146640 649620
rect 146880 649380 146970 649620
rect 147210 649380 147300 649620
rect 147540 649380 147630 649620
rect 147870 649380 147980 649620
rect 148220 649380 148310 649620
rect 148550 649380 148640 649620
rect 148880 649380 148970 649620
rect 149210 649380 149320 649620
rect 149560 649380 149650 649620
rect 149890 649380 149980 649620
rect 150220 649380 150310 649620
rect 150550 649380 150660 649620
rect 150900 649380 150990 649620
rect 151230 649380 151320 649620
rect 151560 649380 151650 649620
rect 151890 649380 152000 649620
rect 152240 649380 152330 649620
rect 152570 649380 152660 649620
rect 152900 649380 152990 649620
rect 153230 649380 153340 649620
rect 153580 649380 153670 649620
rect 153910 649380 154000 649620
rect 154240 649380 154330 649620
rect 154570 649380 154680 649620
rect 154920 649380 155010 649620
rect 155250 649380 155340 649620
rect 155580 649380 155670 649620
rect 155910 649380 155960 649620
rect 110760 649330 155960 649380
rect 159472 652735 164446 660505
rect 159472 647761 188604 652735
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use top  top_0
timestamp 1636213485
transform 1 0 191644 0 1 671360
box -6530 -24030 39650 21850
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
rlabel space 199094 693210 199094 693210 1 MIDDLE
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
