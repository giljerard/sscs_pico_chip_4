magic
tech sky130A
magscale 1 2
timestamp 1636588074
<< metal2 >>
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< metal3 >>
rect 16194 703650 21194 704800
rect 16194 703580 17270 703650
rect 17340 703580 17360 703650
rect 17430 703580 17450 703650
rect 17520 703580 17540 703650
rect 17610 703580 17630 703650
rect 17700 703580 17720 703650
rect 17790 703580 17810 703650
rect 17880 703580 17900 703650
rect 17970 703580 17990 703650
rect 18060 703580 18080 703650
rect 18150 703580 18170 703650
rect 18240 703580 18260 703650
rect 18330 703580 18350 703650
rect 18420 703580 18440 703650
rect 18510 703580 18530 703650
rect 18600 703580 18620 703650
rect 18690 703580 18710 703650
rect 18780 703580 18800 703650
rect 18870 703580 18890 703650
rect 18960 703580 18980 703650
rect 19050 703580 19070 703650
rect 19140 703580 19160 703650
rect 19230 703580 21194 703650
rect 16194 703560 21194 703580
rect 16194 703490 17270 703560
rect 17340 703490 17360 703560
rect 17430 703490 17450 703560
rect 17520 703490 17540 703560
rect 17610 703490 17630 703560
rect 17700 703490 17720 703560
rect 17790 703490 17810 703560
rect 17880 703490 17900 703560
rect 17970 703490 17990 703560
rect 18060 703490 18080 703560
rect 18150 703490 18170 703560
rect 18240 703490 18260 703560
rect 18330 703490 18350 703560
rect 18420 703490 18440 703560
rect 18510 703490 18530 703560
rect 18600 703490 18620 703560
rect 18690 703490 18710 703560
rect 18780 703490 18800 703560
rect 18870 703490 18890 703560
rect 18960 703490 18980 703560
rect 19050 703490 19070 703560
rect 19140 703490 19160 703560
rect 19230 703490 21194 703560
rect 16194 703470 21194 703490
rect 16194 703400 17270 703470
rect 17340 703400 17360 703470
rect 17430 703400 17450 703470
rect 17520 703400 17540 703470
rect 17610 703400 17630 703470
rect 17700 703400 17720 703470
rect 17790 703400 17810 703470
rect 17880 703400 17900 703470
rect 17970 703400 17990 703470
rect 18060 703400 18080 703470
rect 18150 703400 18170 703470
rect 18240 703400 18260 703470
rect 18330 703400 18350 703470
rect 18420 703400 18440 703470
rect 18510 703400 18530 703470
rect 18600 703400 18620 703470
rect 18690 703400 18710 703470
rect 18780 703400 18800 703470
rect 18870 703400 18890 703470
rect 18960 703400 18980 703470
rect 19050 703400 19070 703470
rect 19140 703400 19160 703470
rect 19230 703400 21194 703470
rect 16194 703380 21194 703400
rect 16194 703310 17270 703380
rect 17340 703310 17360 703380
rect 17430 703310 17450 703380
rect 17520 703310 17540 703380
rect 17610 703310 17630 703380
rect 17700 703310 17720 703380
rect 17790 703310 17810 703380
rect 17880 703310 17900 703380
rect 17970 703310 17990 703380
rect 18060 703310 18080 703380
rect 18150 703310 18170 703380
rect 18240 703310 18260 703380
rect 18330 703310 18350 703380
rect 18420 703310 18440 703380
rect 18510 703310 18530 703380
rect 18600 703310 18620 703380
rect 18690 703310 18710 703380
rect 18780 703310 18800 703380
rect 18870 703310 18890 703380
rect 18960 703310 18980 703380
rect 19050 703310 19070 703380
rect 19140 703310 19160 703380
rect 19230 703310 21194 703380
rect 16194 703290 21194 703310
rect 16194 703220 17270 703290
rect 17340 703220 17360 703290
rect 17430 703220 17450 703290
rect 17520 703220 17540 703290
rect 17610 703220 17630 703290
rect 17700 703220 17720 703290
rect 17790 703220 17810 703290
rect 17880 703220 17900 703290
rect 17970 703220 17990 703290
rect 18060 703220 18080 703290
rect 18150 703220 18170 703290
rect 18240 703220 18260 703290
rect 18330 703220 18350 703290
rect 18420 703220 18440 703290
rect 18510 703220 18530 703290
rect 18600 703220 18620 703290
rect 18690 703220 18710 703290
rect 18780 703220 18800 703290
rect 18870 703220 18890 703290
rect 18960 703220 18980 703290
rect 19050 703220 19070 703290
rect 19140 703220 19160 703290
rect 19230 703220 21194 703290
rect 16194 703200 21194 703220
rect 16194 703130 17270 703200
rect 17340 703130 17360 703200
rect 17430 703130 17450 703200
rect 17520 703130 17540 703200
rect 17610 703130 17630 703200
rect 17700 703130 17720 703200
rect 17790 703130 17810 703200
rect 17880 703130 17900 703200
rect 17970 703130 17990 703200
rect 18060 703130 18080 703200
rect 18150 703130 18170 703200
rect 18240 703130 18260 703200
rect 18330 703130 18350 703200
rect 18420 703130 18440 703200
rect 18510 703130 18530 703200
rect 18600 703130 18620 703200
rect 18690 703130 18710 703200
rect 18780 703130 18800 703200
rect 18870 703130 18890 703200
rect 18960 703130 18980 703200
rect 19050 703130 19070 703200
rect 19140 703130 19160 703200
rect 19230 703130 21194 703200
rect 16194 703110 21194 703130
rect 16194 703040 17270 703110
rect 17340 703040 17360 703110
rect 17430 703040 17450 703110
rect 17520 703040 17540 703110
rect 17610 703040 17630 703110
rect 17700 703040 17720 703110
rect 17790 703040 17810 703110
rect 17880 703040 17900 703110
rect 17970 703040 17990 703110
rect 18060 703040 18080 703110
rect 18150 703040 18170 703110
rect 18240 703040 18260 703110
rect 18330 703040 18350 703110
rect 18420 703040 18440 703110
rect 18510 703040 18530 703110
rect 18600 703040 18620 703110
rect 18690 703040 18710 703110
rect 18780 703040 18800 703110
rect 18870 703040 18890 703110
rect 18960 703040 18980 703110
rect 19050 703040 19070 703110
rect 19140 703040 19160 703110
rect 19230 703040 21194 703110
rect 16194 703020 21194 703040
rect 16194 702950 17270 703020
rect 17340 702950 17360 703020
rect 17430 702950 17450 703020
rect 17520 702950 17540 703020
rect 17610 702950 17630 703020
rect 17700 702950 17720 703020
rect 17790 702950 17810 703020
rect 17880 702950 17900 703020
rect 17970 702950 17990 703020
rect 18060 702950 18080 703020
rect 18150 702950 18170 703020
rect 18240 702950 18260 703020
rect 18330 702950 18350 703020
rect 18420 702950 18440 703020
rect 18510 702950 18530 703020
rect 18600 702950 18620 703020
rect 18690 702950 18710 703020
rect 18780 702950 18800 703020
rect 18870 702950 18890 703020
rect 18960 702950 18980 703020
rect 19050 702950 19070 703020
rect 19140 702950 19160 703020
rect 19230 702950 21194 703020
rect 16194 702930 21194 702950
rect 16194 702860 17270 702930
rect 17340 702860 17360 702930
rect 17430 702860 17450 702930
rect 17520 702860 17540 702930
rect 17610 702860 17630 702930
rect 17700 702860 17720 702930
rect 17790 702860 17810 702930
rect 17880 702860 17900 702930
rect 17970 702860 17990 702930
rect 18060 702860 18080 702930
rect 18150 702860 18170 702930
rect 18240 702860 18260 702930
rect 18330 702860 18350 702930
rect 18420 702860 18440 702930
rect 18510 702860 18530 702930
rect 18600 702860 18620 702930
rect 18690 702860 18710 702930
rect 18780 702860 18800 702930
rect 18870 702860 18890 702930
rect 18960 702860 18980 702930
rect 19050 702860 19070 702930
rect 19140 702860 19160 702930
rect 19230 702860 21194 702930
rect 16194 702840 21194 702860
rect 16194 702770 17270 702840
rect 17340 702770 17360 702840
rect 17430 702770 17450 702840
rect 17520 702770 17540 702840
rect 17610 702770 17630 702840
rect 17700 702770 17720 702840
rect 17790 702770 17810 702840
rect 17880 702770 17900 702840
rect 17970 702770 17990 702840
rect 18060 702770 18080 702840
rect 18150 702770 18170 702840
rect 18240 702770 18260 702840
rect 18330 702770 18350 702840
rect 18420 702770 18440 702840
rect 18510 702770 18530 702840
rect 18600 702770 18620 702840
rect 18690 702770 18710 702840
rect 18780 702770 18800 702840
rect 18870 702770 18890 702840
rect 18960 702770 18980 702840
rect 19050 702770 19070 702840
rect 19140 702770 19160 702840
rect 19230 702770 21194 702840
rect 16194 702750 21194 702770
rect 16194 702680 17270 702750
rect 17340 702680 17360 702750
rect 17430 702680 17450 702750
rect 17520 702680 17540 702750
rect 17610 702680 17630 702750
rect 17700 702680 17720 702750
rect 17790 702680 17810 702750
rect 17880 702680 17900 702750
rect 17970 702680 17990 702750
rect 18060 702680 18080 702750
rect 18150 702680 18170 702750
rect 18240 702680 18260 702750
rect 18330 702680 18350 702750
rect 18420 702680 18440 702750
rect 18510 702680 18530 702750
rect 18600 702680 18620 702750
rect 18690 702680 18710 702750
rect 18780 702680 18800 702750
rect 18870 702680 18890 702750
rect 18960 702680 18980 702750
rect 19050 702680 19070 702750
rect 19140 702680 19160 702750
rect 19230 702680 21194 702750
rect 16194 702660 21194 702680
rect 16194 702590 17270 702660
rect 17340 702590 17360 702660
rect 17430 702590 17450 702660
rect 17520 702590 17540 702660
rect 17610 702590 17630 702660
rect 17700 702590 17720 702660
rect 17790 702590 17810 702660
rect 17880 702590 17900 702660
rect 17970 702590 17990 702660
rect 18060 702590 18080 702660
rect 18150 702590 18170 702660
rect 18240 702590 18260 702660
rect 18330 702590 18350 702660
rect 18420 702590 18440 702660
rect 18510 702590 18530 702660
rect 18600 702590 18620 702660
rect 18690 702590 18710 702660
rect 18780 702590 18800 702660
rect 18870 702590 18890 702660
rect 18960 702590 18980 702660
rect 19050 702590 19070 702660
rect 19140 702590 19160 702660
rect 19230 702590 21194 702660
rect 16194 702570 21194 702590
rect 16194 702500 17270 702570
rect 17340 702500 17360 702570
rect 17430 702500 17450 702570
rect 17520 702500 17540 702570
rect 17610 702500 17630 702570
rect 17700 702500 17720 702570
rect 17790 702500 17810 702570
rect 17880 702500 17900 702570
rect 17970 702500 17990 702570
rect 18060 702500 18080 702570
rect 18150 702500 18170 702570
rect 18240 702500 18260 702570
rect 18330 702500 18350 702570
rect 18420 702500 18440 702570
rect 18510 702500 18530 702570
rect 18600 702500 18620 702570
rect 18690 702500 18710 702570
rect 18780 702500 18800 702570
rect 18870 702500 18890 702570
rect 18960 702500 18980 702570
rect 19050 702500 19070 702570
rect 19140 702500 19160 702570
rect 19230 702500 21194 702570
rect 16194 702480 21194 702500
rect 16194 702410 17270 702480
rect 17340 702410 17360 702480
rect 17430 702410 17450 702480
rect 17520 702410 17540 702480
rect 17610 702410 17630 702480
rect 17700 702410 17720 702480
rect 17790 702410 17810 702480
rect 17880 702410 17900 702480
rect 17970 702410 17990 702480
rect 18060 702410 18080 702480
rect 18150 702410 18170 702480
rect 18240 702410 18260 702480
rect 18330 702410 18350 702480
rect 18420 702410 18440 702480
rect 18510 702410 18530 702480
rect 18600 702410 18620 702480
rect 18690 702410 18710 702480
rect 18780 702410 18800 702480
rect 18870 702410 18890 702480
rect 18960 702410 18980 702480
rect 19050 702410 19070 702480
rect 19140 702410 19160 702480
rect 19230 702410 21194 702480
rect 16194 702390 21194 702410
rect 16194 702320 17270 702390
rect 17340 702320 17360 702390
rect 17430 702320 17450 702390
rect 17520 702320 17540 702390
rect 17610 702320 17630 702390
rect 17700 702320 17720 702390
rect 17790 702320 17810 702390
rect 17880 702320 17900 702390
rect 17970 702320 17990 702390
rect 18060 702320 18080 702390
rect 18150 702320 18170 702390
rect 18240 702320 18260 702390
rect 18330 702320 18350 702390
rect 18420 702320 18440 702390
rect 18510 702320 18530 702390
rect 18600 702320 18620 702390
rect 18690 702320 18710 702390
rect 18780 702320 18800 702390
rect 18870 702320 18890 702390
rect 18960 702320 18980 702390
rect 19050 702320 19070 702390
rect 19140 702320 19160 702390
rect 19230 702320 21194 702390
rect 16194 702300 21194 702320
rect 68194 703800 73194 704800
rect 68194 703500 68352 703800
rect 68652 703500 68852 703800
rect 69152 703500 69352 703800
rect 69652 703500 69852 703800
rect 70152 703500 70352 703800
rect 70652 703500 70852 703800
rect 71152 703500 71352 703800
rect 71652 703500 71852 703800
rect 72152 703500 72352 703800
rect 72652 703500 72852 703800
rect 73152 703500 73194 703800
rect 68194 703300 73194 703500
rect 68194 703000 68352 703300
rect 68652 703000 68852 703300
rect 69152 703000 69352 703300
rect 69652 703000 69852 703300
rect 70152 703000 70352 703300
rect 70652 703000 70852 703300
rect 71152 703000 71352 703300
rect 71652 703000 71852 703300
rect 72152 703000 72352 703300
rect 72652 703000 72852 703300
rect 73152 703000 73194 703300
rect 68194 702800 73194 703000
rect 68194 702500 68352 702800
rect 68652 702500 68852 702800
rect 69152 702500 69352 702800
rect 69652 702500 69852 702800
rect 70152 702500 70352 702800
rect 70652 702500 70852 702800
rect 71152 702500 71352 702800
rect 71652 702500 71852 702800
rect 72152 702500 72352 702800
rect 72652 702500 72852 702800
rect 73152 702500 73194 702800
rect 68194 702300 73194 702500
rect 120194 703800 125194 704800
rect 120194 703500 120352 703800
rect 120652 703500 120852 703800
rect 121152 703500 121352 703800
rect 121652 703500 121852 703800
rect 122152 703500 122352 703800
rect 122652 703500 122852 703800
rect 123152 703500 123352 703800
rect 123652 703500 123852 703800
rect 124152 703500 124352 703800
rect 124652 703500 124852 703800
rect 125152 703500 125194 703800
rect 120194 703300 125194 703500
rect 120194 703000 120352 703300
rect 120652 703000 120852 703300
rect 121152 703000 121352 703300
rect 121652 703000 121852 703300
rect 122152 703000 122352 703300
rect 122652 703000 122852 703300
rect 123152 703000 123352 703300
rect 123652 703000 123852 703300
rect 124152 703000 124352 703300
rect 124652 703000 124852 703300
rect 125152 703000 125194 703300
rect 120194 702800 125194 703000
rect 120194 702500 120352 702800
rect 120652 702500 120852 702800
rect 121152 702500 121352 702800
rect 121652 702500 121852 702800
rect 122152 702500 122352 702800
rect 122652 702500 122852 702800
rect 123152 702500 123352 702800
rect 123652 702500 123852 702800
rect 124152 702500 124352 702800
rect 124652 702500 124852 702800
rect 125152 702500 125194 702800
rect 120194 702300 125194 702500
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703110 418394 704800
rect 413394 703040 415760 703110
rect 415830 703040 415850 703110
rect 415920 703040 415940 703110
rect 416010 703040 416030 703110
rect 416100 703040 416120 703110
rect 416190 703040 418394 703110
rect 413394 703020 418394 703040
rect 413394 702950 415760 703020
rect 415830 702950 415850 703020
rect 415920 702950 415940 703020
rect 416010 702950 416030 703020
rect 416100 702950 416120 703020
rect 416190 702950 418394 703020
rect 413394 702930 418394 702950
rect 413394 702860 415760 702930
rect 415830 702860 415850 702930
rect 415920 702860 415940 702930
rect 416010 702860 416030 702930
rect 416100 702860 416120 702930
rect 416190 702860 418394 702930
rect 413394 702840 418394 702860
rect 413394 702770 415760 702840
rect 415830 702770 415850 702840
rect 415920 702770 415940 702840
rect 416010 702770 416030 702840
rect 416100 702770 416120 702840
rect 416190 702770 418394 702840
rect 413394 702750 418394 702770
rect 413394 702680 415760 702750
rect 415830 702680 415850 702750
rect 415920 702680 415940 702750
rect 416010 702680 416030 702750
rect 416100 702680 416120 702750
rect 416190 702680 418394 702750
rect 413394 702300 418394 702680
rect 465394 703110 470394 704800
rect 465394 703040 467010 703110
rect 467080 703040 467100 703110
rect 467170 703040 467190 703110
rect 467260 703040 467280 703110
rect 467350 703040 467370 703110
rect 467440 703040 470394 703110
rect 465394 703020 470394 703040
rect 465394 702950 467010 703020
rect 467080 702950 467100 703020
rect 467170 702950 467190 703020
rect 467260 702950 467280 703020
rect 467350 702950 467370 703020
rect 467440 702950 470394 703020
rect 465394 702930 470394 702950
rect 465394 702860 467010 702930
rect 467080 702860 467100 702930
rect 467170 702860 467190 702930
rect 467260 702860 467280 702930
rect 467350 702860 467370 702930
rect 467440 702860 470394 702930
rect 465394 702840 470394 702860
rect 465394 702770 467010 702840
rect 467080 702770 467100 702840
rect 467170 702770 467190 702840
rect 467260 702770 467280 702840
rect 467350 702770 467370 702840
rect 467440 702770 470394 702840
rect 465394 702750 470394 702770
rect 465394 702680 467010 702750
rect 467080 702680 467100 702750
rect 467170 702680 467190 702750
rect 467260 702680 467280 702750
rect 467350 702680 467370 702750
rect 467440 702680 470394 702750
rect 465394 702300 470394 702680
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 703110 571594 704800
rect 566594 703040 569140 703110
rect 569210 703040 569230 703110
rect 569300 703040 569320 703110
rect 569390 703040 569410 703110
rect 569480 703040 569500 703110
rect 569570 703040 571594 703110
rect 566594 703020 571594 703040
rect 566594 702950 569140 703020
rect 569210 702950 569230 703020
rect 569300 702950 569320 703020
rect 569390 702950 569410 703020
rect 569480 702950 569500 703020
rect 569570 702950 571594 703020
rect 566594 702930 571594 702950
rect 566594 702860 569140 702930
rect 569210 702860 569230 702930
rect 569300 702860 569320 702930
rect 569390 702860 569410 702930
rect 569480 702860 569500 702930
rect 569570 702860 571594 702930
rect 566594 702840 571594 702860
rect 566594 702770 569140 702840
rect 569210 702770 569230 702840
rect 569300 702770 569320 702840
rect 569390 702770 569410 702840
rect 569480 702770 569500 702840
rect 569570 702770 571594 702840
rect 566594 702750 571594 702770
rect 566594 702680 569140 702750
rect 569210 702680 569230 702750
rect 569300 702680 569320 702750
rect 569390 702680 569410 702750
rect 569480 702680 569500 702750
rect 569570 702680 571594 702750
rect 566594 702300 571594 702680
rect -800 683630 1700 685242
rect -800 683560 350 683630
rect 420 683560 440 683630
rect 510 683560 530 683630
rect 600 683560 620 683630
rect 690 683560 710 683630
rect 780 683560 800 683630
rect 870 683560 890 683630
rect 960 683560 980 683630
rect 1050 683560 1070 683630
rect 1140 683560 1160 683630
rect 1230 683560 1250 683630
rect 1320 683560 1340 683630
rect 1410 683560 1430 683630
rect 1500 683560 1520 683630
rect 1590 683560 1610 683630
rect 1680 683560 1700 683630
rect -800 683540 1700 683560
rect -800 683470 350 683540
rect 420 683470 440 683540
rect 510 683470 530 683540
rect 600 683470 620 683540
rect 690 683470 710 683540
rect 780 683470 800 683540
rect 870 683470 890 683540
rect 960 683470 980 683540
rect 1050 683470 1070 683540
rect 1140 683470 1160 683540
rect 1230 683470 1250 683540
rect 1320 683470 1340 683540
rect 1410 683470 1430 683540
rect 1500 683470 1520 683540
rect 1590 683470 1610 683540
rect 1680 683470 1700 683540
rect -800 683450 1700 683470
rect -800 683380 350 683450
rect 420 683380 440 683450
rect 510 683380 530 683450
rect 600 683380 620 683450
rect 690 683380 710 683450
rect 780 683380 800 683450
rect 870 683380 890 683450
rect 960 683380 980 683450
rect 1050 683380 1070 683450
rect 1140 683380 1160 683450
rect 1230 683380 1250 683450
rect 1320 683380 1340 683450
rect 1410 683380 1430 683450
rect 1500 683380 1520 683450
rect 1590 683380 1610 683450
rect 1680 683380 1700 683450
rect -800 683360 1700 683380
rect -800 683290 350 683360
rect 420 683290 440 683360
rect 510 683290 530 683360
rect 600 683290 620 683360
rect 690 683290 710 683360
rect 780 683290 800 683360
rect 870 683290 890 683360
rect 960 683290 980 683360
rect 1050 683290 1070 683360
rect 1140 683290 1160 683360
rect 1230 683290 1250 683360
rect 1320 683290 1340 683360
rect 1410 683290 1430 683360
rect 1500 683290 1520 683360
rect 1590 683290 1610 683360
rect 1680 683290 1700 683360
rect -800 683270 1700 683290
rect -800 683200 350 683270
rect 420 683200 440 683270
rect 510 683200 530 683270
rect 600 683200 620 683270
rect 690 683200 710 683270
rect 780 683200 800 683270
rect 870 683200 890 683270
rect 960 683200 980 683270
rect 1050 683200 1070 683270
rect 1140 683200 1160 683270
rect 1230 683200 1250 683270
rect 1320 683200 1340 683270
rect 1410 683200 1430 683270
rect 1500 683200 1520 683270
rect 1590 683200 1610 683270
rect 1680 683200 1700 683270
rect -800 683180 1700 683200
rect -800 683110 350 683180
rect 420 683110 440 683180
rect 510 683110 530 683180
rect 600 683110 620 683180
rect 690 683110 710 683180
rect 780 683110 800 683180
rect 870 683110 890 683180
rect 960 683110 980 683180
rect 1050 683110 1070 683180
rect 1140 683110 1160 683180
rect 1230 683110 1250 683180
rect 1320 683110 1340 683180
rect 1410 683110 1430 683180
rect 1500 683110 1520 683180
rect 1590 683110 1610 683180
rect 1680 683110 1700 683180
rect -800 683090 1700 683110
rect -800 683020 350 683090
rect 420 683020 440 683090
rect 510 683020 530 683090
rect 600 683020 620 683090
rect 690 683020 710 683090
rect 780 683020 800 683090
rect 870 683020 890 683090
rect 960 683020 980 683090
rect 1050 683020 1070 683090
rect 1140 683020 1160 683090
rect 1230 683020 1250 683090
rect 1320 683020 1340 683090
rect 1410 683020 1430 683090
rect 1500 683020 1520 683090
rect 1590 683020 1610 683090
rect 1680 683020 1700 683090
rect -800 683000 1700 683020
rect -800 682930 350 683000
rect 420 682930 440 683000
rect 510 682930 530 683000
rect 600 682930 620 683000
rect 690 682930 710 683000
rect 780 682930 800 683000
rect 870 682930 890 683000
rect 960 682930 980 683000
rect 1050 682930 1070 683000
rect 1140 682930 1160 683000
rect 1230 682930 1250 683000
rect 1320 682930 1340 683000
rect 1410 682930 1430 683000
rect 1500 682930 1520 683000
rect 1590 682930 1610 683000
rect 1680 682930 1700 683000
rect -800 682910 1700 682930
rect -800 682840 350 682910
rect 420 682840 440 682910
rect 510 682840 530 682910
rect 600 682840 620 682910
rect 690 682840 710 682910
rect 780 682840 800 682910
rect 870 682840 890 682910
rect 960 682840 980 682910
rect 1050 682840 1070 682910
rect 1140 682840 1160 682910
rect 1230 682840 1250 682910
rect 1320 682840 1340 682910
rect 1410 682840 1430 682910
rect 1500 682840 1520 682910
rect 1590 682840 1610 682910
rect 1680 682840 1700 682910
rect -800 682820 1700 682840
rect -800 682750 350 682820
rect 420 682750 440 682820
rect 510 682750 530 682820
rect 600 682750 620 682820
rect 690 682750 710 682820
rect 780 682750 800 682820
rect 870 682750 890 682820
rect 960 682750 980 682820
rect 1050 682750 1070 682820
rect 1140 682750 1160 682820
rect 1230 682750 1250 682820
rect 1320 682750 1340 682820
rect 1410 682750 1430 682820
rect 1500 682750 1520 682820
rect 1590 682750 1610 682820
rect 1680 682750 1700 682820
rect -800 682730 1700 682750
rect -800 682660 350 682730
rect 420 682660 440 682730
rect 510 682660 530 682730
rect 600 682660 620 682730
rect 690 682660 710 682730
rect 780 682660 800 682730
rect 870 682660 890 682730
rect 960 682660 980 682730
rect 1050 682660 1070 682730
rect 1140 682660 1160 682730
rect 1230 682660 1250 682730
rect 1320 682660 1340 682730
rect 1410 682660 1430 682730
rect 1500 682660 1520 682730
rect 1590 682660 1610 682730
rect 1680 682660 1700 682730
rect -800 682640 1700 682660
rect -800 682570 350 682640
rect 420 682570 440 682640
rect 510 682570 530 682640
rect 600 682570 620 682640
rect 690 682570 710 682640
rect 780 682570 800 682640
rect 870 682570 890 682640
rect 960 682570 980 682640
rect 1050 682570 1070 682640
rect 1140 682570 1160 682640
rect 1230 682570 1250 682640
rect 1320 682570 1340 682640
rect 1410 682570 1430 682640
rect 1500 682570 1520 682640
rect 1590 682570 1610 682640
rect 1680 682570 1700 682640
rect -800 682550 1700 682570
rect -800 682480 350 682550
rect 420 682480 440 682550
rect 510 682480 530 682550
rect 600 682480 620 682550
rect 690 682480 710 682550
rect 780 682480 800 682550
rect 870 682480 890 682550
rect 960 682480 980 682550
rect 1050 682480 1070 682550
rect 1140 682480 1160 682550
rect 1230 682480 1250 682550
rect 1320 682480 1340 682550
rect 1410 682480 1430 682550
rect 1500 682480 1520 682550
rect 1590 682480 1610 682550
rect 1680 682480 1700 682550
rect -800 682460 1700 682480
rect -800 682390 350 682460
rect 420 682390 440 682460
rect 510 682390 530 682460
rect 600 682390 620 682460
rect 690 682390 710 682460
rect 780 682390 800 682460
rect 870 682390 890 682460
rect 960 682390 980 682460
rect 1050 682390 1070 682460
rect 1140 682390 1160 682460
rect 1230 682390 1250 682460
rect 1320 682390 1340 682460
rect 1410 682390 1430 682460
rect 1500 682390 1520 682460
rect 1590 682390 1610 682460
rect 1680 682390 1700 682460
rect -800 682370 1700 682390
rect -800 682300 350 682370
rect 420 682300 440 682370
rect 510 682300 530 682370
rect 600 682300 620 682370
rect 690 682300 710 682370
rect 780 682300 800 682370
rect 870 682300 890 682370
rect 960 682300 980 682370
rect 1050 682300 1070 682370
rect 1140 682300 1160 682370
rect 1230 682300 1250 682370
rect 1320 682300 1340 682370
rect 1410 682300 1430 682370
rect 1500 682300 1520 682370
rect 1590 682300 1610 682370
rect 1680 682300 1700 682370
rect -800 682280 1700 682300
rect -800 682210 350 682280
rect 420 682210 440 682280
rect 510 682210 530 682280
rect 600 682210 620 682280
rect 690 682210 710 682280
rect 780 682210 800 682280
rect 870 682210 890 682280
rect 960 682210 980 682280
rect 1050 682210 1070 682280
rect 1140 682210 1160 682280
rect 1230 682210 1250 682280
rect 1320 682210 1340 682280
rect 1410 682210 1430 682280
rect 1500 682210 1520 682280
rect 1590 682210 1610 682280
rect 1680 682210 1700 682280
rect -800 682190 1700 682210
rect -800 682120 350 682190
rect 420 682120 440 682190
rect 510 682120 530 682190
rect 600 682120 620 682190
rect 690 682120 710 682190
rect 780 682120 800 682190
rect 870 682120 890 682190
rect 960 682120 980 682190
rect 1050 682120 1070 682190
rect 1140 682120 1160 682190
rect 1230 682120 1250 682190
rect 1320 682120 1340 682190
rect 1410 682120 1430 682190
rect 1500 682120 1520 682190
rect 1590 682120 1610 682190
rect 1680 682120 1700 682190
rect -800 682100 1700 682120
rect -800 682030 350 682100
rect 420 682030 440 682100
rect 510 682030 530 682100
rect 600 682030 620 682100
rect 690 682030 710 682100
rect 780 682030 800 682100
rect 870 682030 890 682100
rect 960 682030 980 682100
rect 1050 682030 1070 682100
rect 1140 682030 1160 682100
rect 1230 682030 1250 682100
rect 1320 682030 1340 682100
rect 1410 682030 1430 682100
rect 1500 682030 1520 682100
rect 1590 682030 1610 682100
rect 1680 682030 1700 682100
rect -800 682010 1700 682030
rect -800 681940 350 682010
rect 420 681940 440 682010
rect 510 681940 530 682010
rect 600 681940 620 682010
rect 690 681940 710 682010
rect 780 681940 800 682010
rect 870 681940 890 682010
rect 960 681940 980 682010
rect 1050 681940 1070 682010
rect 1140 681940 1160 682010
rect 1230 681940 1250 682010
rect 1320 681940 1340 682010
rect 1410 681940 1430 682010
rect 1500 681940 1520 682010
rect 1590 681940 1610 682010
rect 1680 681940 1700 682010
rect -800 681920 1700 681940
rect -800 681850 350 681920
rect 420 681850 440 681920
rect 510 681850 530 681920
rect 600 681850 620 681920
rect 690 681850 710 681920
rect 780 681850 800 681920
rect 870 681850 890 681920
rect 960 681850 980 681920
rect 1050 681850 1070 681920
rect 1140 681850 1160 681920
rect 1230 681850 1250 681920
rect 1320 681850 1340 681920
rect 1410 681850 1430 681920
rect 1500 681850 1520 681920
rect 1590 681850 1610 681920
rect 1680 681850 1700 681920
rect -800 681830 1700 681850
rect -800 681760 350 681830
rect 420 681760 440 681830
rect 510 681760 530 681830
rect 600 681760 620 681830
rect 690 681760 710 681830
rect 780 681760 800 681830
rect 870 681760 890 681830
rect 960 681760 980 681830
rect 1050 681760 1070 681830
rect 1140 681760 1160 681830
rect 1230 681760 1250 681830
rect 1320 681760 1340 681830
rect 1410 681760 1430 681830
rect 1500 681760 1520 681830
rect 1590 681760 1610 681830
rect 1680 681760 1700 681830
rect -800 681740 1700 681760
rect -800 681670 350 681740
rect 420 681670 440 681740
rect 510 681670 530 681740
rect 600 681670 620 681740
rect 690 681670 710 681740
rect 780 681670 800 681740
rect 870 681670 890 681740
rect 960 681670 980 681740
rect 1050 681670 1070 681740
rect 1140 681670 1160 681740
rect 1230 681670 1250 681740
rect 1320 681670 1340 681740
rect 1410 681670 1430 681740
rect 1500 681670 1520 681740
rect 1590 681670 1610 681740
rect 1680 681670 1700 681740
rect -800 680242 1700 681670
rect 582300 681110 584800 682984
rect 582300 681040 582680 681110
rect 582750 681040 582770 681110
rect 582840 681040 582860 681110
rect 582930 681040 582950 681110
rect 583020 681040 583040 681110
rect 583110 681040 584800 681110
rect 582300 681020 584800 681040
rect 582300 680950 582680 681020
rect 582750 680950 582770 681020
rect 582840 680950 582860 681020
rect 582930 680950 582950 681020
rect 583020 680950 583040 681020
rect 583110 680950 584800 681020
rect 582300 680930 584800 680950
rect 582300 680860 582680 680930
rect 582750 680860 582770 680930
rect 582840 680860 582860 680930
rect 582930 680860 582950 680930
rect 583020 680860 583040 680930
rect 583110 680860 584800 680930
rect 582300 680840 584800 680860
rect 582300 680770 582680 680840
rect 582750 680770 582770 680840
rect 582840 680770 582860 680840
rect 582930 680770 582950 680840
rect 583020 680770 583040 680840
rect 583110 680770 584800 680840
rect 582300 680750 584800 680770
rect 582300 680680 582680 680750
rect 582750 680680 582770 680750
rect 582840 680680 582860 680750
rect 582930 680680 582950 680750
rect 583020 680680 583040 680750
rect 583110 680680 584800 680750
rect 582300 677984 584800 680680
rect -800 643842 1660 648642
rect 582340 639784 584800 644584
rect -800 633842 1660 638642
rect 94254 638170 94574 638390
rect 94254 638100 94280 638170
rect 94350 638100 94380 638170
rect 94450 638100 94480 638170
rect 94550 638100 94574 638170
rect 94254 638080 94574 638100
rect 94254 638010 94280 638080
rect 94350 638010 94380 638080
rect 94450 638010 94480 638080
rect 94550 638010 94574 638080
rect 94254 637980 94574 638010
rect 98814 638170 99134 638390
rect 98814 638100 98838 638170
rect 98908 638100 98938 638170
rect 99008 638100 99038 638170
rect 99108 638100 99134 638170
rect 98814 638080 99134 638100
rect 98814 638010 98838 638080
rect 98908 638010 98938 638080
rect 99008 638010 99038 638080
rect 99108 638010 99134 638080
rect 98814 637980 99134 638010
rect 582340 629784 584800 634584
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 17270 703580 17340 703650
rect 17360 703580 17430 703650
rect 17450 703580 17520 703650
rect 17540 703580 17610 703650
rect 17630 703580 17700 703650
rect 17720 703580 17790 703650
rect 17810 703580 17880 703650
rect 17900 703580 17970 703650
rect 17990 703580 18060 703650
rect 18080 703580 18150 703650
rect 18170 703580 18240 703650
rect 18260 703580 18330 703650
rect 18350 703580 18420 703650
rect 18440 703580 18510 703650
rect 18530 703580 18600 703650
rect 18620 703580 18690 703650
rect 18710 703580 18780 703650
rect 18800 703580 18870 703650
rect 18890 703580 18960 703650
rect 18980 703580 19050 703650
rect 19070 703580 19140 703650
rect 19160 703580 19230 703650
rect 17270 703490 17340 703560
rect 17360 703490 17430 703560
rect 17450 703490 17520 703560
rect 17540 703490 17610 703560
rect 17630 703490 17700 703560
rect 17720 703490 17790 703560
rect 17810 703490 17880 703560
rect 17900 703490 17970 703560
rect 17990 703490 18060 703560
rect 18080 703490 18150 703560
rect 18170 703490 18240 703560
rect 18260 703490 18330 703560
rect 18350 703490 18420 703560
rect 18440 703490 18510 703560
rect 18530 703490 18600 703560
rect 18620 703490 18690 703560
rect 18710 703490 18780 703560
rect 18800 703490 18870 703560
rect 18890 703490 18960 703560
rect 18980 703490 19050 703560
rect 19070 703490 19140 703560
rect 19160 703490 19230 703560
rect 17270 703400 17340 703470
rect 17360 703400 17430 703470
rect 17450 703400 17520 703470
rect 17540 703400 17610 703470
rect 17630 703400 17700 703470
rect 17720 703400 17790 703470
rect 17810 703400 17880 703470
rect 17900 703400 17970 703470
rect 17990 703400 18060 703470
rect 18080 703400 18150 703470
rect 18170 703400 18240 703470
rect 18260 703400 18330 703470
rect 18350 703400 18420 703470
rect 18440 703400 18510 703470
rect 18530 703400 18600 703470
rect 18620 703400 18690 703470
rect 18710 703400 18780 703470
rect 18800 703400 18870 703470
rect 18890 703400 18960 703470
rect 18980 703400 19050 703470
rect 19070 703400 19140 703470
rect 19160 703400 19230 703470
rect 17270 703310 17340 703380
rect 17360 703310 17430 703380
rect 17450 703310 17520 703380
rect 17540 703310 17610 703380
rect 17630 703310 17700 703380
rect 17720 703310 17790 703380
rect 17810 703310 17880 703380
rect 17900 703310 17970 703380
rect 17990 703310 18060 703380
rect 18080 703310 18150 703380
rect 18170 703310 18240 703380
rect 18260 703310 18330 703380
rect 18350 703310 18420 703380
rect 18440 703310 18510 703380
rect 18530 703310 18600 703380
rect 18620 703310 18690 703380
rect 18710 703310 18780 703380
rect 18800 703310 18870 703380
rect 18890 703310 18960 703380
rect 18980 703310 19050 703380
rect 19070 703310 19140 703380
rect 19160 703310 19230 703380
rect 17270 703220 17340 703290
rect 17360 703220 17430 703290
rect 17450 703220 17520 703290
rect 17540 703220 17610 703290
rect 17630 703220 17700 703290
rect 17720 703220 17790 703290
rect 17810 703220 17880 703290
rect 17900 703220 17970 703290
rect 17990 703220 18060 703290
rect 18080 703220 18150 703290
rect 18170 703220 18240 703290
rect 18260 703220 18330 703290
rect 18350 703220 18420 703290
rect 18440 703220 18510 703290
rect 18530 703220 18600 703290
rect 18620 703220 18690 703290
rect 18710 703220 18780 703290
rect 18800 703220 18870 703290
rect 18890 703220 18960 703290
rect 18980 703220 19050 703290
rect 19070 703220 19140 703290
rect 19160 703220 19230 703290
rect 17270 703130 17340 703200
rect 17360 703130 17430 703200
rect 17450 703130 17520 703200
rect 17540 703130 17610 703200
rect 17630 703130 17700 703200
rect 17720 703130 17790 703200
rect 17810 703130 17880 703200
rect 17900 703130 17970 703200
rect 17990 703130 18060 703200
rect 18080 703130 18150 703200
rect 18170 703130 18240 703200
rect 18260 703130 18330 703200
rect 18350 703130 18420 703200
rect 18440 703130 18510 703200
rect 18530 703130 18600 703200
rect 18620 703130 18690 703200
rect 18710 703130 18780 703200
rect 18800 703130 18870 703200
rect 18890 703130 18960 703200
rect 18980 703130 19050 703200
rect 19070 703130 19140 703200
rect 19160 703130 19230 703200
rect 17270 703040 17340 703110
rect 17360 703040 17430 703110
rect 17450 703040 17520 703110
rect 17540 703040 17610 703110
rect 17630 703040 17700 703110
rect 17720 703040 17790 703110
rect 17810 703040 17880 703110
rect 17900 703040 17970 703110
rect 17990 703040 18060 703110
rect 18080 703040 18150 703110
rect 18170 703040 18240 703110
rect 18260 703040 18330 703110
rect 18350 703040 18420 703110
rect 18440 703040 18510 703110
rect 18530 703040 18600 703110
rect 18620 703040 18690 703110
rect 18710 703040 18780 703110
rect 18800 703040 18870 703110
rect 18890 703040 18960 703110
rect 18980 703040 19050 703110
rect 19070 703040 19140 703110
rect 19160 703040 19230 703110
rect 17270 702950 17340 703020
rect 17360 702950 17430 703020
rect 17450 702950 17520 703020
rect 17540 702950 17610 703020
rect 17630 702950 17700 703020
rect 17720 702950 17790 703020
rect 17810 702950 17880 703020
rect 17900 702950 17970 703020
rect 17990 702950 18060 703020
rect 18080 702950 18150 703020
rect 18170 702950 18240 703020
rect 18260 702950 18330 703020
rect 18350 702950 18420 703020
rect 18440 702950 18510 703020
rect 18530 702950 18600 703020
rect 18620 702950 18690 703020
rect 18710 702950 18780 703020
rect 18800 702950 18870 703020
rect 18890 702950 18960 703020
rect 18980 702950 19050 703020
rect 19070 702950 19140 703020
rect 19160 702950 19230 703020
rect 17270 702860 17340 702930
rect 17360 702860 17430 702930
rect 17450 702860 17520 702930
rect 17540 702860 17610 702930
rect 17630 702860 17700 702930
rect 17720 702860 17790 702930
rect 17810 702860 17880 702930
rect 17900 702860 17970 702930
rect 17990 702860 18060 702930
rect 18080 702860 18150 702930
rect 18170 702860 18240 702930
rect 18260 702860 18330 702930
rect 18350 702860 18420 702930
rect 18440 702860 18510 702930
rect 18530 702860 18600 702930
rect 18620 702860 18690 702930
rect 18710 702860 18780 702930
rect 18800 702860 18870 702930
rect 18890 702860 18960 702930
rect 18980 702860 19050 702930
rect 19070 702860 19140 702930
rect 19160 702860 19230 702930
rect 17270 702770 17340 702840
rect 17360 702770 17430 702840
rect 17450 702770 17520 702840
rect 17540 702770 17610 702840
rect 17630 702770 17700 702840
rect 17720 702770 17790 702840
rect 17810 702770 17880 702840
rect 17900 702770 17970 702840
rect 17990 702770 18060 702840
rect 18080 702770 18150 702840
rect 18170 702770 18240 702840
rect 18260 702770 18330 702840
rect 18350 702770 18420 702840
rect 18440 702770 18510 702840
rect 18530 702770 18600 702840
rect 18620 702770 18690 702840
rect 18710 702770 18780 702840
rect 18800 702770 18870 702840
rect 18890 702770 18960 702840
rect 18980 702770 19050 702840
rect 19070 702770 19140 702840
rect 19160 702770 19230 702840
rect 17270 702680 17340 702750
rect 17360 702680 17430 702750
rect 17450 702680 17520 702750
rect 17540 702680 17610 702750
rect 17630 702680 17700 702750
rect 17720 702680 17790 702750
rect 17810 702680 17880 702750
rect 17900 702680 17970 702750
rect 17990 702680 18060 702750
rect 18080 702680 18150 702750
rect 18170 702680 18240 702750
rect 18260 702680 18330 702750
rect 18350 702680 18420 702750
rect 18440 702680 18510 702750
rect 18530 702680 18600 702750
rect 18620 702680 18690 702750
rect 18710 702680 18780 702750
rect 18800 702680 18870 702750
rect 18890 702680 18960 702750
rect 18980 702680 19050 702750
rect 19070 702680 19140 702750
rect 19160 702680 19230 702750
rect 17270 702590 17340 702660
rect 17360 702590 17430 702660
rect 17450 702590 17520 702660
rect 17540 702590 17610 702660
rect 17630 702590 17700 702660
rect 17720 702590 17790 702660
rect 17810 702590 17880 702660
rect 17900 702590 17970 702660
rect 17990 702590 18060 702660
rect 18080 702590 18150 702660
rect 18170 702590 18240 702660
rect 18260 702590 18330 702660
rect 18350 702590 18420 702660
rect 18440 702590 18510 702660
rect 18530 702590 18600 702660
rect 18620 702590 18690 702660
rect 18710 702590 18780 702660
rect 18800 702590 18870 702660
rect 18890 702590 18960 702660
rect 18980 702590 19050 702660
rect 19070 702590 19140 702660
rect 19160 702590 19230 702660
rect 17270 702500 17340 702570
rect 17360 702500 17430 702570
rect 17450 702500 17520 702570
rect 17540 702500 17610 702570
rect 17630 702500 17700 702570
rect 17720 702500 17790 702570
rect 17810 702500 17880 702570
rect 17900 702500 17970 702570
rect 17990 702500 18060 702570
rect 18080 702500 18150 702570
rect 18170 702500 18240 702570
rect 18260 702500 18330 702570
rect 18350 702500 18420 702570
rect 18440 702500 18510 702570
rect 18530 702500 18600 702570
rect 18620 702500 18690 702570
rect 18710 702500 18780 702570
rect 18800 702500 18870 702570
rect 18890 702500 18960 702570
rect 18980 702500 19050 702570
rect 19070 702500 19140 702570
rect 19160 702500 19230 702570
rect 17270 702410 17340 702480
rect 17360 702410 17430 702480
rect 17450 702410 17520 702480
rect 17540 702410 17610 702480
rect 17630 702410 17700 702480
rect 17720 702410 17790 702480
rect 17810 702410 17880 702480
rect 17900 702410 17970 702480
rect 17990 702410 18060 702480
rect 18080 702410 18150 702480
rect 18170 702410 18240 702480
rect 18260 702410 18330 702480
rect 18350 702410 18420 702480
rect 18440 702410 18510 702480
rect 18530 702410 18600 702480
rect 18620 702410 18690 702480
rect 18710 702410 18780 702480
rect 18800 702410 18870 702480
rect 18890 702410 18960 702480
rect 18980 702410 19050 702480
rect 19070 702410 19140 702480
rect 19160 702410 19230 702480
rect 17270 702320 17340 702390
rect 17360 702320 17430 702390
rect 17450 702320 17520 702390
rect 17540 702320 17610 702390
rect 17630 702320 17700 702390
rect 17720 702320 17790 702390
rect 17810 702320 17880 702390
rect 17900 702320 17970 702390
rect 17990 702320 18060 702390
rect 18080 702320 18150 702390
rect 18170 702320 18240 702390
rect 18260 702320 18330 702390
rect 18350 702320 18420 702390
rect 18440 702320 18510 702390
rect 18530 702320 18600 702390
rect 18620 702320 18690 702390
rect 18710 702320 18780 702390
rect 18800 702320 18870 702390
rect 18890 702320 18960 702390
rect 18980 702320 19050 702390
rect 19070 702320 19140 702390
rect 19160 702320 19230 702390
rect 68352 703500 68652 703800
rect 68852 703500 69152 703800
rect 69352 703500 69652 703800
rect 69852 703500 70152 703800
rect 70352 703500 70652 703800
rect 70852 703500 71152 703800
rect 71352 703500 71652 703800
rect 71852 703500 72152 703800
rect 72352 703500 72652 703800
rect 72852 703500 73152 703800
rect 68352 703000 68652 703300
rect 68852 703000 69152 703300
rect 69352 703000 69652 703300
rect 69852 703000 70152 703300
rect 70352 703000 70652 703300
rect 70852 703000 71152 703300
rect 71352 703000 71652 703300
rect 71852 703000 72152 703300
rect 72352 703000 72652 703300
rect 72852 703000 73152 703300
rect 68352 702500 68652 702800
rect 68852 702500 69152 702800
rect 69352 702500 69652 702800
rect 69852 702500 70152 702800
rect 70352 702500 70652 702800
rect 70852 702500 71152 702800
rect 71352 702500 71652 702800
rect 71852 702500 72152 702800
rect 72352 702500 72652 702800
rect 72852 702500 73152 702800
rect 120352 703500 120652 703800
rect 120852 703500 121152 703800
rect 121352 703500 121652 703800
rect 121852 703500 122152 703800
rect 122352 703500 122652 703800
rect 122852 703500 123152 703800
rect 123352 703500 123652 703800
rect 123852 703500 124152 703800
rect 124352 703500 124652 703800
rect 124852 703500 125152 703800
rect 120352 703000 120652 703300
rect 120852 703000 121152 703300
rect 121352 703000 121652 703300
rect 121852 703000 122152 703300
rect 122352 703000 122652 703300
rect 122852 703000 123152 703300
rect 123352 703000 123652 703300
rect 123852 703000 124152 703300
rect 124352 703000 124652 703300
rect 124852 703000 125152 703300
rect 120352 702500 120652 702800
rect 120852 702500 121152 702800
rect 121352 702500 121652 702800
rect 121852 702500 122152 702800
rect 122352 702500 122652 702800
rect 122852 702500 123152 702800
rect 123352 702500 123652 702800
rect 123852 702500 124152 702800
rect 124352 702500 124652 702800
rect 124852 702500 125152 702800
rect 415760 703040 415830 703110
rect 415850 703040 415920 703110
rect 415940 703040 416010 703110
rect 416030 703040 416100 703110
rect 416120 703040 416190 703110
rect 415760 702950 415830 703020
rect 415850 702950 415920 703020
rect 415940 702950 416010 703020
rect 416030 702950 416100 703020
rect 416120 702950 416190 703020
rect 415760 702860 415830 702930
rect 415850 702860 415920 702930
rect 415940 702860 416010 702930
rect 416030 702860 416100 702930
rect 416120 702860 416190 702930
rect 415760 702770 415830 702840
rect 415850 702770 415920 702840
rect 415940 702770 416010 702840
rect 416030 702770 416100 702840
rect 416120 702770 416190 702840
rect 415760 702680 415830 702750
rect 415850 702680 415920 702750
rect 415940 702680 416010 702750
rect 416030 702680 416100 702750
rect 416120 702680 416190 702750
rect 467010 703040 467080 703110
rect 467100 703040 467170 703110
rect 467190 703040 467260 703110
rect 467280 703040 467350 703110
rect 467370 703040 467440 703110
rect 467010 702950 467080 703020
rect 467100 702950 467170 703020
rect 467190 702950 467260 703020
rect 467280 702950 467350 703020
rect 467370 702950 467440 703020
rect 467010 702860 467080 702930
rect 467100 702860 467170 702930
rect 467190 702860 467260 702930
rect 467280 702860 467350 702930
rect 467370 702860 467440 702930
rect 467010 702770 467080 702840
rect 467100 702770 467170 702840
rect 467190 702770 467260 702840
rect 467280 702770 467350 702840
rect 467370 702770 467440 702840
rect 467010 702680 467080 702750
rect 467100 702680 467170 702750
rect 467190 702680 467260 702750
rect 467280 702680 467350 702750
rect 467370 702680 467440 702750
rect 569140 703040 569210 703110
rect 569230 703040 569300 703110
rect 569320 703040 569390 703110
rect 569410 703040 569480 703110
rect 569500 703040 569570 703110
rect 569140 702950 569210 703020
rect 569230 702950 569300 703020
rect 569320 702950 569390 703020
rect 569410 702950 569480 703020
rect 569500 702950 569570 703020
rect 569140 702860 569210 702930
rect 569230 702860 569300 702930
rect 569320 702860 569390 702930
rect 569410 702860 569480 702930
rect 569500 702860 569570 702930
rect 569140 702770 569210 702840
rect 569230 702770 569300 702840
rect 569320 702770 569390 702840
rect 569410 702770 569480 702840
rect 569500 702770 569570 702840
rect 569140 702680 569210 702750
rect 569230 702680 569300 702750
rect 569320 702680 569390 702750
rect 569410 702680 569480 702750
rect 569500 702680 569570 702750
rect 350 683560 420 683630
rect 440 683560 510 683630
rect 530 683560 600 683630
rect 620 683560 690 683630
rect 710 683560 780 683630
rect 800 683560 870 683630
rect 890 683560 960 683630
rect 980 683560 1050 683630
rect 1070 683560 1140 683630
rect 1160 683560 1230 683630
rect 1250 683560 1320 683630
rect 1340 683560 1410 683630
rect 1430 683560 1500 683630
rect 1520 683560 1590 683630
rect 1610 683560 1680 683630
rect 350 683470 420 683540
rect 440 683470 510 683540
rect 530 683470 600 683540
rect 620 683470 690 683540
rect 710 683470 780 683540
rect 800 683470 870 683540
rect 890 683470 960 683540
rect 980 683470 1050 683540
rect 1070 683470 1140 683540
rect 1160 683470 1230 683540
rect 1250 683470 1320 683540
rect 1340 683470 1410 683540
rect 1430 683470 1500 683540
rect 1520 683470 1590 683540
rect 1610 683470 1680 683540
rect 350 683380 420 683450
rect 440 683380 510 683450
rect 530 683380 600 683450
rect 620 683380 690 683450
rect 710 683380 780 683450
rect 800 683380 870 683450
rect 890 683380 960 683450
rect 980 683380 1050 683450
rect 1070 683380 1140 683450
rect 1160 683380 1230 683450
rect 1250 683380 1320 683450
rect 1340 683380 1410 683450
rect 1430 683380 1500 683450
rect 1520 683380 1590 683450
rect 1610 683380 1680 683450
rect 350 683290 420 683360
rect 440 683290 510 683360
rect 530 683290 600 683360
rect 620 683290 690 683360
rect 710 683290 780 683360
rect 800 683290 870 683360
rect 890 683290 960 683360
rect 980 683290 1050 683360
rect 1070 683290 1140 683360
rect 1160 683290 1230 683360
rect 1250 683290 1320 683360
rect 1340 683290 1410 683360
rect 1430 683290 1500 683360
rect 1520 683290 1590 683360
rect 1610 683290 1680 683360
rect 350 683200 420 683270
rect 440 683200 510 683270
rect 530 683200 600 683270
rect 620 683200 690 683270
rect 710 683200 780 683270
rect 800 683200 870 683270
rect 890 683200 960 683270
rect 980 683200 1050 683270
rect 1070 683200 1140 683270
rect 1160 683200 1230 683270
rect 1250 683200 1320 683270
rect 1340 683200 1410 683270
rect 1430 683200 1500 683270
rect 1520 683200 1590 683270
rect 1610 683200 1680 683270
rect 350 683110 420 683180
rect 440 683110 510 683180
rect 530 683110 600 683180
rect 620 683110 690 683180
rect 710 683110 780 683180
rect 800 683110 870 683180
rect 890 683110 960 683180
rect 980 683110 1050 683180
rect 1070 683110 1140 683180
rect 1160 683110 1230 683180
rect 1250 683110 1320 683180
rect 1340 683110 1410 683180
rect 1430 683110 1500 683180
rect 1520 683110 1590 683180
rect 1610 683110 1680 683180
rect 350 683020 420 683090
rect 440 683020 510 683090
rect 530 683020 600 683090
rect 620 683020 690 683090
rect 710 683020 780 683090
rect 800 683020 870 683090
rect 890 683020 960 683090
rect 980 683020 1050 683090
rect 1070 683020 1140 683090
rect 1160 683020 1230 683090
rect 1250 683020 1320 683090
rect 1340 683020 1410 683090
rect 1430 683020 1500 683090
rect 1520 683020 1590 683090
rect 1610 683020 1680 683090
rect 350 682930 420 683000
rect 440 682930 510 683000
rect 530 682930 600 683000
rect 620 682930 690 683000
rect 710 682930 780 683000
rect 800 682930 870 683000
rect 890 682930 960 683000
rect 980 682930 1050 683000
rect 1070 682930 1140 683000
rect 1160 682930 1230 683000
rect 1250 682930 1320 683000
rect 1340 682930 1410 683000
rect 1430 682930 1500 683000
rect 1520 682930 1590 683000
rect 1610 682930 1680 683000
rect 350 682840 420 682910
rect 440 682840 510 682910
rect 530 682840 600 682910
rect 620 682840 690 682910
rect 710 682840 780 682910
rect 800 682840 870 682910
rect 890 682840 960 682910
rect 980 682840 1050 682910
rect 1070 682840 1140 682910
rect 1160 682840 1230 682910
rect 1250 682840 1320 682910
rect 1340 682840 1410 682910
rect 1430 682840 1500 682910
rect 1520 682840 1590 682910
rect 1610 682840 1680 682910
rect 350 682750 420 682820
rect 440 682750 510 682820
rect 530 682750 600 682820
rect 620 682750 690 682820
rect 710 682750 780 682820
rect 800 682750 870 682820
rect 890 682750 960 682820
rect 980 682750 1050 682820
rect 1070 682750 1140 682820
rect 1160 682750 1230 682820
rect 1250 682750 1320 682820
rect 1340 682750 1410 682820
rect 1430 682750 1500 682820
rect 1520 682750 1590 682820
rect 1610 682750 1680 682820
rect 350 682660 420 682730
rect 440 682660 510 682730
rect 530 682660 600 682730
rect 620 682660 690 682730
rect 710 682660 780 682730
rect 800 682660 870 682730
rect 890 682660 960 682730
rect 980 682660 1050 682730
rect 1070 682660 1140 682730
rect 1160 682660 1230 682730
rect 1250 682660 1320 682730
rect 1340 682660 1410 682730
rect 1430 682660 1500 682730
rect 1520 682660 1590 682730
rect 1610 682660 1680 682730
rect 350 682570 420 682640
rect 440 682570 510 682640
rect 530 682570 600 682640
rect 620 682570 690 682640
rect 710 682570 780 682640
rect 800 682570 870 682640
rect 890 682570 960 682640
rect 980 682570 1050 682640
rect 1070 682570 1140 682640
rect 1160 682570 1230 682640
rect 1250 682570 1320 682640
rect 1340 682570 1410 682640
rect 1430 682570 1500 682640
rect 1520 682570 1590 682640
rect 1610 682570 1680 682640
rect 350 682480 420 682550
rect 440 682480 510 682550
rect 530 682480 600 682550
rect 620 682480 690 682550
rect 710 682480 780 682550
rect 800 682480 870 682550
rect 890 682480 960 682550
rect 980 682480 1050 682550
rect 1070 682480 1140 682550
rect 1160 682480 1230 682550
rect 1250 682480 1320 682550
rect 1340 682480 1410 682550
rect 1430 682480 1500 682550
rect 1520 682480 1590 682550
rect 1610 682480 1680 682550
rect 350 682390 420 682460
rect 440 682390 510 682460
rect 530 682390 600 682460
rect 620 682390 690 682460
rect 710 682390 780 682460
rect 800 682390 870 682460
rect 890 682390 960 682460
rect 980 682390 1050 682460
rect 1070 682390 1140 682460
rect 1160 682390 1230 682460
rect 1250 682390 1320 682460
rect 1340 682390 1410 682460
rect 1430 682390 1500 682460
rect 1520 682390 1590 682460
rect 1610 682390 1680 682460
rect 350 682300 420 682370
rect 440 682300 510 682370
rect 530 682300 600 682370
rect 620 682300 690 682370
rect 710 682300 780 682370
rect 800 682300 870 682370
rect 890 682300 960 682370
rect 980 682300 1050 682370
rect 1070 682300 1140 682370
rect 1160 682300 1230 682370
rect 1250 682300 1320 682370
rect 1340 682300 1410 682370
rect 1430 682300 1500 682370
rect 1520 682300 1590 682370
rect 1610 682300 1680 682370
rect 350 682210 420 682280
rect 440 682210 510 682280
rect 530 682210 600 682280
rect 620 682210 690 682280
rect 710 682210 780 682280
rect 800 682210 870 682280
rect 890 682210 960 682280
rect 980 682210 1050 682280
rect 1070 682210 1140 682280
rect 1160 682210 1230 682280
rect 1250 682210 1320 682280
rect 1340 682210 1410 682280
rect 1430 682210 1500 682280
rect 1520 682210 1590 682280
rect 1610 682210 1680 682280
rect 350 682120 420 682190
rect 440 682120 510 682190
rect 530 682120 600 682190
rect 620 682120 690 682190
rect 710 682120 780 682190
rect 800 682120 870 682190
rect 890 682120 960 682190
rect 980 682120 1050 682190
rect 1070 682120 1140 682190
rect 1160 682120 1230 682190
rect 1250 682120 1320 682190
rect 1340 682120 1410 682190
rect 1430 682120 1500 682190
rect 1520 682120 1590 682190
rect 1610 682120 1680 682190
rect 350 682030 420 682100
rect 440 682030 510 682100
rect 530 682030 600 682100
rect 620 682030 690 682100
rect 710 682030 780 682100
rect 800 682030 870 682100
rect 890 682030 960 682100
rect 980 682030 1050 682100
rect 1070 682030 1140 682100
rect 1160 682030 1230 682100
rect 1250 682030 1320 682100
rect 1340 682030 1410 682100
rect 1430 682030 1500 682100
rect 1520 682030 1590 682100
rect 1610 682030 1680 682100
rect 350 681940 420 682010
rect 440 681940 510 682010
rect 530 681940 600 682010
rect 620 681940 690 682010
rect 710 681940 780 682010
rect 800 681940 870 682010
rect 890 681940 960 682010
rect 980 681940 1050 682010
rect 1070 681940 1140 682010
rect 1160 681940 1230 682010
rect 1250 681940 1320 682010
rect 1340 681940 1410 682010
rect 1430 681940 1500 682010
rect 1520 681940 1590 682010
rect 1610 681940 1680 682010
rect 350 681850 420 681920
rect 440 681850 510 681920
rect 530 681850 600 681920
rect 620 681850 690 681920
rect 710 681850 780 681920
rect 800 681850 870 681920
rect 890 681850 960 681920
rect 980 681850 1050 681920
rect 1070 681850 1140 681920
rect 1160 681850 1230 681920
rect 1250 681850 1320 681920
rect 1340 681850 1410 681920
rect 1430 681850 1500 681920
rect 1520 681850 1590 681920
rect 1610 681850 1680 681920
rect 350 681760 420 681830
rect 440 681760 510 681830
rect 530 681760 600 681830
rect 620 681760 690 681830
rect 710 681760 780 681830
rect 800 681760 870 681830
rect 890 681760 960 681830
rect 980 681760 1050 681830
rect 1070 681760 1140 681830
rect 1160 681760 1230 681830
rect 1250 681760 1320 681830
rect 1340 681760 1410 681830
rect 1430 681760 1500 681830
rect 1520 681760 1590 681830
rect 1610 681760 1680 681830
rect 350 681670 420 681740
rect 440 681670 510 681740
rect 530 681670 600 681740
rect 620 681670 690 681740
rect 710 681670 780 681740
rect 800 681670 870 681740
rect 890 681670 960 681740
rect 980 681670 1050 681740
rect 1070 681670 1140 681740
rect 1160 681670 1230 681740
rect 1250 681670 1320 681740
rect 1340 681670 1410 681740
rect 1430 681670 1500 681740
rect 1520 681670 1590 681740
rect 1610 681670 1680 681740
rect 582680 681040 582750 681110
rect 582770 681040 582840 681110
rect 582860 681040 582930 681110
rect 582950 681040 583020 681110
rect 583040 681040 583110 681110
rect 582680 680950 582750 681020
rect 582770 680950 582840 681020
rect 582860 680950 582930 681020
rect 582950 680950 583020 681020
rect 583040 680950 583110 681020
rect 582680 680860 582750 680930
rect 582770 680860 582840 680930
rect 582860 680860 582930 680930
rect 582950 680860 583020 680930
rect 583040 680860 583110 680930
rect 582680 680770 582750 680840
rect 582770 680770 582840 680840
rect 582860 680770 582930 680840
rect 582950 680770 583020 680840
rect 583040 680770 583110 680840
rect 582680 680680 582750 680750
rect 582770 680680 582840 680750
rect 582860 680680 582930 680750
rect 582950 680680 583020 680750
rect 583040 680680 583110 680750
rect 94280 638100 94350 638170
rect 94380 638100 94450 638170
rect 94480 638100 94550 638170
rect 94280 638010 94350 638080
rect 94380 638010 94450 638080
rect 94480 638010 94550 638080
rect 98838 638100 98908 638170
rect 98938 638100 99008 638170
rect 99038 638100 99108 638170
rect 98838 638010 98908 638080
rect 98938 638010 99008 638080
rect 99038 638010 99108 638080
<< metal4 >>
rect 68194 703800 73194 704000
rect 17246 703650 19246 703652
rect 17246 703580 17270 703650
rect 17340 703580 17360 703650
rect 17430 703580 17450 703650
rect 17520 703580 17540 703650
rect 17610 703580 17630 703650
rect 17700 703580 17720 703650
rect 17790 703580 17810 703650
rect 17880 703580 17900 703650
rect 17970 703580 17990 703650
rect 18060 703580 18080 703650
rect 18150 703580 18170 703650
rect 18240 703580 18260 703650
rect 18330 703580 18350 703650
rect 18420 703580 18440 703650
rect 18510 703580 18530 703650
rect 18600 703580 18620 703650
rect 18690 703580 18710 703650
rect 18780 703580 18800 703650
rect 18870 703580 18890 703650
rect 18960 703580 18980 703650
rect 19050 703580 19070 703650
rect 19140 703580 19160 703650
rect 19230 703580 19246 703650
rect 17246 703560 19246 703580
rect 17246 703490 17270 703560
rect 17340 703490 17360 703560
rect 17430 703490 17450 703560
rect 17520 703490 17540 703560
rect 17610 703490 17630 703560
rect 17700 703490 17720 703560
rect 17790 703490 17810 703560
rect 17880 703490 17900 703560
rect 17970 703490 17990 703560
rect 18060 703490 18080 703560
rect 18150 703490 18170 703560
rect 18240 703490 18260 703560
rect 18330 703490 18350 703560
rect 18420 703490 18440 703560
rect 18510 703490 18530 703560
rect 18600 703490 18620 703560
rect 18690 703490 18710 703560
rect 18780 703490 18800 703560
rect 18870 703490 18890 703560
rect 18960 703490 18980 703560
rect 19050 703490 19070 703560
rect 19140 703490 19160 703560
rect 19230 703490 19246 703560
rect 17246 703470 19246 703490
rect 17246 703400 17270 703470
rect 17340 703400 17360 703470
rect 17430 703400 17450 703470
rect 17520 703400 17540 703470
rect 17610 703400 17630 703470
rect 17700 703400 17720 703470
rect 17790 703400 17810 703470
rect 17880 703400 17900 703470
rect 17970 703400 17990 703470
rect 18060 703400 18080 703470
rect 18150 703400 18170 703470
rect 18240 703400 18260 703470
rect 18330 703400 18350 703470
rect 18420 703400 18440 703470
rect 18510 703400 18530 703470
rect 18600 703400 18620 703470
rect 18690 703400 18710 703470
rect 18780 703400 18800 703470
rect 18870 703400 18890 703470
rect 18960 703400 18980 703470
rect 19050 703400 19070 703470
rect 19140 703400 19160 703470
rect 19230 703400 19246 703470
rect 17246 703380 19246 703400
rect 17246 703310 17270 703380
rect 17340 703310 17360 703380
rect 17430 703310 17450 703380
rect 17520 703310 17540 703380
rect 17610 703310 17630 703380
rect 17700 703310 17720 703380
rect 17790 703310 17810 703380
rect 17880 703310 17900 703380
rect 17970 703310 17990 703380
rect 18060 703310 18080 703380
rect 18150 703310 18170 703380
rect 18240 703310 18260 703380
rect 18330 703310 18350 703380
rect 18420 703310 18440 703380
rect 18510 703310 18530 703380
rect 18600 703310 18620 703380
rect 18690 703310 18710 703380
rect 18780 703310 18800 703380
rect 18870 703310 18890 703380
rect 18960 703310 18980 703380
rect 19050 703310 19070 703380
rect 19140 703310 19160 703380
rect 19230 703310 19246 703380
rect 17246 703290 19246 703310
rect 17246 703220 17270 703290
rect 17340 703220 17360 703290
rect 17430 703220 17450 703290
rect 17520 703220 17540 703290
rect 17610 703220 17630 703290
rect 17700 703220 17720 703290
rect 17790 703220 17810 703290
rect 17880 703220 17900 703290
rect 17970 703220 17990 703290
rect 18060 703220 18080 703290
rect 18150 703220 18170 703290
rect 18240 703220 18260 703290
rect 18330 703220 18350 703290
rect 18420 703220 18440 703290
rect 18510 703220 18530 703290
rect 18600 703220 18620 703290
rect 18690 703220 18710 703290
rect 18780 703220 18800 703290
rect 18870 703220 18890 703290
rect 18960 703220 18980 703290
rect 19050 703220 19070 703290
rect 19140 703220 19160 703290
rect 19230 703220 19246 703290
rect 17246 703200 19246 703220
rect 17246 703130 17270 703200
rect 17340 703130 17360 703200
rect 17430 703130 17450 703200
rect 17520 703130 17540 703200
rect 17610 703130 17630 703200
rect 17700 703130 17720 703200
rect 17790 703130 17810 703200
rect 17880 703130 17900 703200
rect 17970 703130 17990 703200
rect 18060 703130 18080 703200
rect 18150 703130 18170 703200
rect 18240 703130 18260 703200
rect 18330 703130 18350 703200
rect 18420 703130 18440 703200
rect 18510 703130 18530 703200
rect 18600 703130 18620 703200
rect 18690 703130 18710 703200
rect 18780 703130 18800 703200
rect 18870 703130 18890 703200
rect 18960 703130 18980 703200
rect 19050 703130 19070 703200
rect 19140 703130 19160 703200
rect 19230 703130 19246 703200
rect 17246 703110 19246 703130
rect 17246 703040 17270 703110
rect 17340 703040 17360 703110
rect 17430 703040 17450 703110
rect 17520 703040 17540 703110
rect 17610 703040 17630 703110
rect 17700 703040 17720 703110
rect 17790 703040 17810 703110
rect 17880 703040 17900 703110
rect 17970 703040 17990 703110
rect 18060 703040 18080 703110
rect 18150 703040 18170 703110
rect 18240 703040 18260 703110
rect 18330 703040 18350 703110
rect 18420 703040 18440 703110
rect 18510 703040 18530 703110
rect 18600 703040 18620 703110
rect 18690 703040 18710 703110
rect 18780 703040 18800 703110
rect 18870 703040 18890 703110
rect 18960 703040 18980 703110
rect 19050 703040 19070 703110
rect 19140 703040 19160 703110
rect 19230 703040 19246 703110
rect 17246 703020 19246 703040
rect 17246 702950 17270 703020
rect 17340 702950 17360 703020
rect 17430 702950 17450 703020
rect 17520 702950 17540 703020
rect 17610 702950 17630 703020
rect 17700 702950 17720 703020
rect 17790 702950 17810 703020
rect 17880 702950 17900 703020
rect 17970 702950 17990 703020
rect 18060 702950 18080 703020
rect 18150 702950 18170 703020
rect 18240 702950 18260 703020
rect 18330 702950 18350 703020
rect 18420 702950 18440 703020
rect 18510 702950 18530 703020
rect 18600 702950 18620 703020
rect 18690 702950 18710 703020
rect 18780 702950 18800 703020
rect 18870 702950 18890 703020
rect 18960 702950 18980 703020
rect 19050 702950 19070 703020
rect 19140 702950 19160 703020
rect 19230 702950 19246 703020
rect 17246 702930 19246 702950
rect 17246 702860 17270 702930
rect 17340 702860 17360 702930
rect 17430 702860 17450 702930
rect 17520 702860 17540 702930
rect 17610 702860 17630 702930
rect 17700 702860 17720 702930
rect 17790 702860 17810 702930
rect 17880 702860 17900 702930
rect 17970 702860 17990 702930
rect 18060 702860 18080 702930
rect 18150 702860 18170 702930
rect 18240 702860 18260 702930
rect 18330 702860 18350 702930
rect 18420 702860 18440 702930
rect 18510 702860 18530 702930
rect 18600 702860 18620 702930
rect 18690 702860 18710 702930
rect 18780 702860 18800 702930
rect 18870 702860 18890 702930
rect 18960 702860 18980 702930
rect 19050 702860 19070 702930
rect 19140 702860 19160 702930
rect 19230 702860 19246 702930
rect 17246 702840 19246 702860
rect 17246 702770 17270 702840
rect 17340 702770 17360 702840
rect 17430 702770 17450 702840
rect 17520 702770 17540 702840
rect 17610 702770 17630 702840
rect 17700 702770 17720 702840
rect 17790 702770 17810 702840
rect 17880 702770 17900 702840
rect 17970 702770 17990 702840
rect 18060 702770 18080 702840
rect 18150 702770 18170 702840
rect 18240 702770 18260 702840
rect 18330 702770 18350 702840
rect 18420 702770 18440 702840
rect 18510 702770 18530 702840
rect 18600 702770 18620 702840
rect 18690 702770 18710 702840
rect 18780 702770 18800 702840
rect 18870 702770 18890 702840
rect 18960 702770 18980 702840
rect 19050 702770 19070 702840
rect 19140 702770 19160 702840
rect 19230 702770 19246 702840
rect 17246 702750 19246 702770
rect 17246 702680 17270 702750
rect 17340 702680 17360 702750
rect 17430 702680 17450 702750
rect 17520 702680 17540 702750
rect 17610 702680 17630 702750
rect 17700 702680 17720 702750
rect 17790 702680 17810 702750
rect 17880 702680 17900 702750
rect 17970 702680 17990 702750
rect 18060 702680 18080 702750
rect 18150 702680 18170 702750
rect 18240 702680 18260 702750
rect 18330 702680 18350 702750
rect 18420 702680 18440 702750
rect 18510 702680 18530 702750
rect 18600 702680 18620 702750
rect 18690 702680 18710 702750
rect 18780 702680 18800 702750
rect 18870 702680 18890 702750
rect 18960 702680 18980 702750
rect 19050 702680 19070 702750
rect 19140 702680 19160 702750
rect 19230 702680 19246 702750
rect 17246 702660 19246 702680
rect 17246 702590 17270 702660
rect 17340 702590 17360 702660
rect 17430 702590 17450 702660
rect 17520 702590 17540 702660
rect 17610 702590 17630 702660
rect 17700 702590 17720 702660
rect 17790 702590 17810 702660
rect 17880 702590 17900 702660
rect 17970 702590 17990 702660
rect 18060 702590 18080 702660
rect 18150 702590 18170 702660
rect 18240 702590 18260 702660
rect 18330 702590 18350 702660
rect 18420 702590 18440 702660
rect 18510 702590 18530 702660
rect 18600 702590 18620 702660
rect 18690 702590 18710 702660
rect 18780 702590 18800 702660
rect 18870 702590 18890 702660
rect 18960 702590 18980 702660
rect 19050 702590 19070 702660
rect 19140 702590 19160 702660
rect 19230 702590 19246 702660
rect 17246 702570 19246 702590
rect 17246 702500 17270 702570
rect 17340 702500 17360 702570
rect 17430 702500 17450 702570
rect 17520 702500 17540 702570
rect 17610 702500 17630 702570
rect 17700 702500 17720 702570
rect 17790 702500 17810 702570
rect 17880 702500 17900 702570
rect 17970 702500 17990 702570
rect 18060 702500 18080 702570
rect 18150 702500 18170 702570
rect 18240 702500 18260 702570
rect 18330 702500 18350 702570
rect 18420 702500 18440 702570
rect 18510 702500 18530 702570
rect 18600 702500 18620 702570
rect 18690 702500 18710 702570
rect 18780 702500 18800 702570
rect 18870 702500 18890 702570
rect 18960 702500 18980 702570
rect 19050 702500 19070 702570
rect 19140 702500 19160 702570
rect 19230 702500 19246 702570
rect 17246 702480 19246 702500
rect 17246 702410 17270 702480
rect 17340 702410 17360 702480
rect 17430 702410 17450 702480
rect 17520 702410 17540 702480
rect 17610 702410 17630 702480
rect 17700 702410 17720 702480
rect 17790 702410 17810 702480
rect 17880 702410 17900 702480
rect 17970 702410 17990 702480
rect 18060 702410 18080 702480
rect 18150 702410 18170 702480
rect 18240 702410 18260 702480
rect 18330 702410 18350 702480
rect 18420 702410 18440 702480
rect 18510 702410 18530 702480
rect 18600 702410 18620 702480
rect 18690 702410 18710 702480
rect 18780 702410 18800 702480
rect 18870 702410 18890 702480
rect 18960 702410 18980 702480
rect 19050 702410 19070 702480
rect 19140 702410 19160 702480
rect 19230 702410 19246 702480
rect 17246 702390 19246 702410
rect 17246 702320 17270 702390
rect 17340 702320 17360 702390
rect 17430 702320 17450 702390
rect 17520 702320 17540 702390
rect 17610 702320 17630 702390
rect 17700 702320 17720 702390
rect 17790 702320 17810 702390
rect 17880 702320 17900 702390
rect 17970 702320 17990 702390
rect 18060 702320 18080 702390
rect 18150 702320 18170 702390
rect 18240 702320 18260 702390
rect 18330 702320 18350 702390
rect 18420 702320 18440 702390
rect 18510 702320 18530 702390
rect 18600 702320 18620 702390
rect 18690 702320 18710 702390
rect 18780 702320 18800 702390
rect 18870 702320 18890 702390
rect 18960 702320 18980 702390
rect 19050 702320 19070 702390
rect 19140 702320 19160 702390
rect 19230 702320 19246 702390
rect 17246 697254 19246 702320
rect 68194 703500 68352 703800
rect 68652 703500 68852 703800
rect 69152 703500 69352 703800
rect 69652 703500 69852 703800
rect 70152 703500 70352 703800
rect 70652 703500 70852 703800
rect 71152 703500 71352 703800
rect 71652 703500 71852 703800
rect 72152 703500 72352 703800
rect 72652 703500 72852 703800
rect 73152 703500 73194 703800
rect 68194 703300 73194 703500
rect 68194 703000 68352 703300
rect 68652 703000 68852 703300
rect 69152 703000 69352 703300
rect 69652 703000 69852 703300
rect 70152 703000 70352 703300
rect 70652 703000 70852 703300
rect 71152 703000 71352 703300
rect 71652 703000 71852 703300
rect 72152 703000 72352 703300
rect 72652 703000 72852 703300
rect 73152 703000 73194 703300
rect 68194 702800 73194 703000
rect 68194 702500 68352 702800
rect 68652 702500 68852 702800
rect 69152 702500 69352 702800
rect 69652 702500 69852 702800
rect 70152 702500 70352 702800
rect 70652 702500 70852 702800
rect 71152 702500 71352 702800
rect 71652 702500 71852 702800
rect 72152 702500 72352 702800
rect 72652 702500 72852 702800
rect 73152 702500 73194 702800
rect 68194 702300 73194 702500
rect 120194 703800 125194 704000
rect 120194 703500 120352 703800
rect 120652 703500 120852 703800
rect 121152 703500 121352 703800
rect 121652 703500 121852 703800
rect 122152 703500 122352 703800
rect 122652 703500 122852 703800
rect 123152 703500 123352 703800
rect 123652 703500 123852 703800
rect 124152 703500 124352 703800
rect 124652 703500 124852 703800
rect 125152 703500 125194 703800
rect 120194 703300 125194 703500
rect 120194 703000 120352 703300
rect 120652 703000 120852 703300
rect 121152 703000 121352 703300
rect 121652 703000 121852 703300
rect 122152 703000 122352 703300
rect 122652 703000 122852 703300
rect 123152 703000 123352 703300
rect 123652 703000 123852 703300
rect 124152 703000 124352 703300
rect 124652 703000 124852 703300
rect 125152 703000 125194 703300
rect 120194 702800 125194 703000
rect 120194 702500 120352 702800
rect 120652 702500 120852 702800
rect 121152 702500 121352 702800
rect 121652 702500 121852 702800
rect 122152 702500 122352 702800
rect 122652 702500 122852 702800
rect 123152 702500 123352 702800
rect 123652 702500 123852 702800
rect 124152 702500 124352 702800
rect 124652 702500 124852 702800
rect 125152 702500 125194 702800
rect 120194 702300 125194 702500
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 415740 703110 416220 703170
rect 415740 703040 415760 703110
rect 415830 703040 415850 703110
rect 415920 703040 415940 703110
rect 416010 703040 416030 703110
rect 416100 703040 416120 703110
rect 416190 703040 416220 703110
rect 415740 703020 416220 703040
rect 415740 702950 415760 703020
rect 415830 702950 415850 703020
rect 415920 702950 415940 703020
rect 416010 702950 416030 703020
rect 416100 702950 416120 703020
rect 416190 702950 416220 703020
rect 415740 702930 416220 702950
rect 415740 702860 415760 702930
rect 415830 702860 415850 702930
rect 415920 702860 415940 702930
rect 416010 702860 416030 702930
rect 416100 702860 416120 702930
rect 416190 702860 416220 702930
rect 415740 702840 416220 702860
rect 415740 702770 415760 702840
rect 415830 702770 415850 702840
rect 415920 702770 415940 702840
rect 416010 702770 416030 702840
rect 416100 702770 416120 702840
rect 416190 702770 416220 702840
rect 415740 702750 416220 702770
rect 415740 702680 415760 702750
rect 415830 702680 415850 702750
rect 415920 702680 415940 702750
rect 416010 702680 416030 702750
rect 416100 702680 416120 702750
rect 416190 702680 416220 702750
rect 321017 701268 321497 702300
rect 415740 701268 416220 702680
rect 466990 703110 467470 703170
rect 466990 703040 467010 703110
rect 467080 703040 467100 703110
rect 467170 703040 467190 703110
rect 467260 703040 467280 703110
rect 467350 703040 467370 703110
rect 467440 703040 467470 703110
rect 466990 703020 467470 703040
rect 466990 702950 467010 703020
rect 467080 702950 467100 703020
rect 467170 702950 467190 703020
rect 467260 702950 467280 703020
rect 467350 702950 467370 703020
rect 467440 702950 467470 703020
rect 466990 702930 467470 702950
rect 466990 702860 467010 702930
rect 467080 702860 467100 702930
rect 467170 702860 467190 702930
rect 467260 702860 467280 702930
rect 467350 702860 467370 702930
rect 467440 702860 467470 702930
rect 466990 702840 467470 702860
rect 466990 702770 467010 702840
rect 467080 702770 467100 702840
rect 467170 702770 467190 702840
rect 467260 702770 467280 702840
rect 467350 702770 467370 702840
rect 467440 702770 467470 702840
rect 466990 702750 467470 702770
rect 466990 702680 467010 702750
rect 467080 702680 467100 702750
rect 467170 702680 467190 702750
rect 467260 702680 467280 702750
rect 467350 702680 467370 702750
rect 467440 702680 467470 702750
rect 466990 701268 467470 702680
rect 569120 703110 569600 703170
rect 569120 703040 569140 703110
rect 569210 703040 569230 703110
rect 569300 703040 569320 703110
rect 569390 703040 569410 703110
rect 569480 703040 569500 703110
rect 569570 703040 569600 703110
rect 569120 703020 569600 703040
rect 569120 702950 569140 703020
rect 569210 702950 569230 703020
rect 569300 702950 569320 703020
rect 569390 702950 569410 703020
rect 569480 702950 569500 703020
rect 569570 702950 569600 703020
rect 569120 702930 569600 702950
rect 569120 702860 569140 702930
rect 569210 702860 569230 702930
rect 569300 702860 569320 702930
rect 569390 702860 569410 702930
rect 569480 702860 569500 702930
rect 569570 702860 569600 702930
rect 569120 702840 569600 702860
rect 569120 702770 569140 702840
rect 569210 702770 569230 702840
rect 569300 702770 569320 702840
rect 569390 702770 569410 702840
rect 569480 702770 569500 702840
rect 569570 702770 569600 702840
rect 569120 702750 569600 702770
rect 569120 702680 569140 702750
rect 569210 702680 569230 702750
rect 569300 702680 569320 702750
rect 569390 702680 569410 702750
rect 569480 702680 569500 702750
rect 569570 702680 569600 702750
rect 569120 701268 569600 702680
rect 131494 684668 146744 685148
rect 272 683630 4312 683653
rect 272 683560 350 683630
rect 420 683560 440 683630
rect 510 683560 530 683630
rect 600 683560 620 683630
rect 690 683560 710 683630
rect 780 683560 800 683630
rect 870 683560 890 683630
rect 960 683560 980 683630
rect 1050 683560 1070 683630
rect 1140 683560 1160 683630
rect 1230 683560 1250 683630
rect 1320 683560 1340 683630
rect 1410 683560 1430 683630
rect 1500 683560 1520 683630
rect 1590 683560 1610 683630
rect 1680 683560 4312 683630
rect 272 683540 4312 683560
rect 272 683470 350 683540
rect 420 683470 440 683540
rect 510 683470 530 683540
rect 600 683470 620 683540
rect 690 683470 710 683540
rect 780 683470 800 683540
rect 870 683470 890 683540
rect 960 683470 980 683540
rect 1050 683470 1070 683540
rect 1140 683470 1160 683540
rect 1230 683470 1250 683540
rect 1320 683470 1340 683540
rect 1410 683470 1430 683540
rect 1500 683470 1520 683540
rect 1590 683470 1610 683540
rect 1680 683470 4312 683540
rect 272 683450 4312 683470
rect 272 683380 350 683450
rect 420 683380 440 683450
rect 510 683380 530 683450
rect 600 683380 620 683450
rect 690 683380 710 683450
rect 780 683380 800 683450
rect 870 683380 890 683450
rect 960 683380 980 683450
rect 1050 683380 1070 683450
rect 1140 683380 1160 683450
rect 1230 683380 1250 683450
rect 1320 683380 1340 683450
rect 1410 683380 1430 683450
rect 1500 683380 1520 683450
rect 1590 683380 1610 683450
rect 1680 683380 4312 683450
rect 272 683360 4312 683380
rect 272 683290 350 683360
rect 420 683290 440 683360
rect 510 683290 530 683360
rect 600 683290 620 683360
rect 690 683290 710 683360
rect 780 683290 800 683360
rect 870 683290 890 683360
rect 960 683290 980 683360
rect 1050 683290 1070 683360
rect 1140 683290 1160 683360
rect 1230 683290 1250 683360
rect 1320 683290 1340 683360
rect 1410 683290 1430 683360
rect 1500 683290 1520 683360
rect 1590 683290 1610 683360
rect 1680 683290 4312 683360
rect 272 683270 4312 683290
rect 272 683200 350 683270
rect 420 683200 440 683270
rect 510 683200 530 683270
rect 600 683200 620 683270
rect 690 683200 710 683270
rect 780 683200 800 683270
rect 870 683200 890 683270
rect 960 683200 980 683270
rect 1050 683200 1070 683270
rect 1140 683200 1160 683270
rect 1230 683200 1250 683270
rect 1320 683200 1340 683270
rect 1410 683200 1430 683270
rect 1500 683200 1520 683270
rect 1590 683200 1610 683270
rect 1680 683200 4312 683270
rect 272 683180 4312 683200
rect 272 683110 350 683180
rect 420 683110 440 683180
rect 510 683110 530 683180
rect 600 683110 620 683180
rect 690 683110 710 683180
rect 780 683110 800 683180
rect 870 683110 890 683180
rect 960 683110 980 683180
rect 1050 683110 1070 683180
rect 1140 683110 1160 683180
rect 1230 683110 1250 683180
rect 1320 683110 1340 683180
rect 1410 683110 1430 683180
rect 1500 683110 1520 683180
rect 1590 683110 1610 683180
rect 1680 683110 4312 683180
rect 272 683090 4312 683110
rect 272 683020 350 683090
rect 420 683020 440 683090
rect 510 683020 530 683090
rect 600 683020 620 683090
rect 690 683020 710 683090
rect 780 683020 800 683090
rect 870 683020 890 683090
rect 960 683020 980 683090
rect 1050 683020 1070 683090
rect 1140 683020 1160 683090
rect 1230 683020 1250 683090
rect 1320 683020 1340 683090
rect 1410 683020 1430 683090
rect 1500 683020 1520 683090
rect 1590 683020 1610 683090
rect 1680 683020 4312 683090
rect 272 683000 4312 683020
rect 272 682930 350 683000
rect 420 682930 440 683000
rect 510 682930 530 683000
rect 600 682930 620 683000
rect 690 682930 710 683000
rect 780 682930 800 683000
rect 870 682930 890 683000
rect 960 682930 980 683000
rect 1050 682930 1070 683000
rect 1140 682930 1160 683000
rect 1230 682930 1250 683000
rect 1320 682930 1340 683000
rect 1410 682930 1430 683000
rect 1500 682930 1520 683000
rect 1590 682930 1610 683000
rect 1680 682930 4312 683000
rect 272 682910 4312 682930
rect 272 682840 350 682910
rect 420 682840 440 682910
rect 510 682840 530 682910
rect 600 682840 620 682910
rect 690 682840 710 682910
rect 780 682840 800 682910
rect 870 682840 890 682910
rect 960 682840 980 682910
rect 1050 682840 1070 682910
rect 1140 682840 1160 682910
rect 1230 682840 1250 682910
rect 1320 682840 1340 682910
rect 1410 682840 1430 682910
rect 1500 682840 1520 682910
rect 1590 682840 1610 682910
rect 1680 682840 4312 682910
rect 272 682820 4312 682840
rect 272 682750 350 682820
rect 420 682750 440 682820
rect 510 682750 530 682820
rect 600 682750 620 682820
rect 690 682750 710 682820
rect 780 682750 800 682820
rect 870 682750 890 682820
rect 960 682750 980 682820
rect 1050 682750 1070 682820
rect 1140 682750 1160 682820
rect 1230 682750 1250 682820
rect 1320 682750 1340 682820
rect 1410 682750 1430 682820
rect 1500 682750 1520 682820
rect 1590 682750 1610 682820
rect 1680 682750 4312 682820
rect 272 682730 4312 682750
rect 272 682660 350 682730
rect 420 682660 440 682730
rect 510 682660 530 682730
rect 600 682660 620 682730
rect 690 682660 710 682730
rect 780 682660 800 682730
rect 870 682660 890 682730
rect 960 682660 980 682730
rect 1050 682660 1070 682730
rect 1140 682660 1160 682730
rect 1230 682660 1250 682730
rect 1320 682660 1340 682730
rect 1410 682660 1430 682730
rect 1500 682660 1520 682730
rect 1590 682660 1610 682730
rect 1680 682660 4312 682730
rect 272 682640 4312 682660
rect 272 682570 350 682640
rect 420 682570 440 682640
rect 510 682570 530 682640
rect 600 682570 620 682640
rect 690 682570 710 682640
rect 780 682570 800 682640
rect 870 682570 890 682640
rect 960 682570 980 682640
rect 1050 682570 1070 682640
rect 1140 682570 1160 682640
rect 1230 682570 1250 682640
rect 1320 682570 1340 682640
rect 1410 682570 1430 682640
rect 1500 682570 1520 682640
rect 1590 682570 1610 682640
rect 1680 682570 4312 682640
rect 272 682550 4312 682570
rect 272 682480 350 682550
rect 420 682480 440 682550
rect 510 682480 530 682550
rect 600 682480 620 682550
rect 690 682480 710 682550
rect 780 682480 800 682550
rect 870 682480 890 682550
rect 960 682480 980 682550
rect 1050 682480 1070 682550
rect 1140 682480 1160 682550
rect 1230 682480 1250 682550
rect 1320 682480 1340 682550
rect 1410 682480 1430 682550
rect 1500 682480 1520 682550
rect 1590 682480 1610 682550
rect 1680 682480 4312 682550
rect 272 682460 4312 682480
rect 272 682390 350 682460
rect 420 682390 440 682460
rect 510 682390 530 682460
rect 600 682390 620 682460
rect 690 682390 710 682460
rect 780 682390 800 682460
rect 870 682390 890 682460
rect 960 682390 980 682460
rect 1050 682390 1070 682460
rect 1140 682390 1160 682460
rect 1230 682390 1250 682460
rect 1320 682390 1340 682460
rect 1410 682390 1430 682460
rect 1500 682390 1520 682460
rect 1590 682390 1610 682460
rect 1680 682390 4312 682460
rect 272 682370 4312 682390
rect 272 682300 350 682370
rect 420 682300 440 682370
rect 510 682300 530 682370
rect 600 682300 620 682370
rect 690 682300 710 682370
rect 780 682300 800 682370
rect 870 682300 890 682370
rect 960 682300 980 682370
rect 1050 682300 1070 682370
rect 1140 682300 1160 682370
rect 1230 682300 1250 682370
rect 1320 682300 1340 682370
rect 1410 682300 1430 682370
rect 1500 682300 1520 682370
rect 1590 682300 1610 682370
rect 1680 682300 4312 682370
rect 272 682280 4312 682300
rect 272 682210 350 682280
rect 420 682210 440 682280
rect 510 682210 530 682280
rect 600 682210 620 682280
rect 690 682210 710 682280
rect 780 682210 800 682280
rect 870 682210 890 682280
rect 960 682210 980 682280
rect 1050 682210 1070 682280
rect 1140 682210 1160 682280
rect 1230 682210 1250 682280
rect 1320 682210 1340 682280
rect 1410 682210 1430 682280
rect 1500 682210 1520 682280
rect 1590 682210 1610 682280
rect 1680 682210 4312 682280
rect 272 682190 4312 682210
rect 272 682120 350 682190
rect 420 682120 440 682190
rect 510 682120 530 682190
rect 600 682120 620 682190
rect 690 682120 710 682190
rect 780 682120 800 682190
rect 870 682120 890 682190
rect 960 682120 980 682190
rect 1050 682120 1070 682190
rect 1140 682120 1160 682190
rect 1230 682120 1250 682190
rect 1320 682120 1340 682190
rect 1410 682120 1430 682190
rect 1500 682120 1520 682190
rect 1590 682120 1610 682190
rect 1680 682120 4312 682190
rect 272 682100 4312 682120
rect 272 682030 350 682100
rect 420 682030 440 682100
rect 510 682030 530 682100
rect 600 682030 620 682100
rect 690 682030 710 682100
rect 780 682030 800 682100
rect 870 682030 890 682100
rect 960 682030 980 682100
rect 1050 682030 1070 682100
rect 1140 682030 1160 682100
rect 1230 682030 1250 682100
rect 1320 682030 1340 682100
rect 1410 682030 1430 682100
rect 1500 682030 1520 682100
rect 1590 682030 1610 682100
rect 1680 682030 4312 682100
rect 272 682010 4312 682030
rect 272 681940 350 682010
rect 420 681940 440 682010
rect 510 681940 530 682010
rect 600 681940 620 682010
rect 690 681940 710 682010
rect 780 681940 800 682010
rect 870 681940 890 682010
rect 960 681940 980 682010
rect 1050 681940 1070 682010
rect 1140 681940 1160 682010
rect 1230 681940 1250 682010
rect 1320 681940 1340 682010
rect 1410 681940 1430 682010
rect 1500 681940 1520 682010
rect 1590 681940 1610 682010
rect 1680 681940 4312 682010
rect 272 681920 4312 681940
rect 272 681850 350 681920
rect 420 681850 440 681920
rect 510 681850 530 681920
rect 600 681850 620 681920
rect 690 681850 710 681920
rect 780 681850 800 681920
rect 870 681850 890 681920
rect 960 681850 980 681920
rect 1050 681850 1070 681920
rect 1140 681850 1160 681920
rect 1230 681850 1250 681920
rect 1320 681850 1340 681920
rect 1410 681850 1430 681920
rect 1500 681850 1520 681920
rect 1590 681850 1610 681920
rect 1680 681850 4312 681920
rect 272 681830 4312 681850
rect 272 681760 350 681830
rect 420 681760 440 681830
rect 510 681760 530 681830
rect 600 681760 620 681830
rect 690 681760 710 681830
rect 780 681760 800 681830
rect 870 681760 890 681830
rect 960 681760 980 681830
rect 1050 681760 1070 681830
rect 1140 681760 1160 681830
rect 1230 681760 1250 681830
rect 1320 681760 1340 681830
rect 1410 681760 1430 681830
rect 1500 681760 1520 681830
rect 1590 681760 1610 681830
rect 1680 681760 4312 681830
rect 272 681740 4312 681760
rect 272 681670 350 681740
rect 420 681670 440 681740
rect 510 681670 530 681740
rect 600 681670 620 681740
rect 690 681670 710 681740
rect 780 681670 800 681740
rect 870 681670 890 681740
rect 960 681670 980 681740
rect 1050 681670 1070 681740
rect 1140 681670 1160 681740
rect 1230 681670 1250 681740
rect 1320 681670 1340 681740
rect 1410 681670 1430 681740
rect 1500 681670 1520 681740
rect 1590 681670 1610 681740
rect 1680 681670 4312 681740
rect 272 681653 4312 681670
rect 131494 672350 131974 684668
rect 110364 671870 131974 672350
rect 132937 683454 146744 683931
rect 110364 670830 110524 671870
rect 132937 670640 133414 683454
rect 128410 670160 133414 670640
rect 134191 682386 146744 682866
rect 134191 651640 134671 682386
rect 120014 651320 134671 651640
rect 135741 680669 146744 681160
rect 580942 681130 581422 688518
rect 580942 681110 583170 681130
rect 580942 681040 582680 681110
rect 582750 681040 582770 681110
rect 582840 681040 582860 681110
rect 582930 681040 582950 681110
rect 583020 681040 583040 681110
rect 583110 681040 583170 681110
rect 580942 681020 583170 681040
rect 580942 680950 582680 681020
rect 582750 680950 582770 681020
rect 582840 680950 582860 681020
rect 582930 680950 582950 681020
rect 583020 680950 583040 681020
rect 583110 680950 583170 681020
rect 580942 680930 583170 680950
rect 580942 680860 582680 680930
rect 582750 680860 582770 680930
rect 582840 680860 582860 680930
rect 582930 680860 582950 680930
rect 583020 680860 583040 680930
rect 583110 680860 583170 680930
rect 580942 680840 583170 680860
rect 580942 680770 582680 680840
rect 582750 680770 582770 680840
rect 582840 680770 582860 680840
rect 582930 680770 582950 680840
rect 583020 680770 583040 680840
rect 583110 680770 583170 680840
rect 580942 680750 583170 680770
rect 580942 680680 582680 680750
rect 582750 680680 582770 680750
rect 582840 680680 582860 680750
rect 582930 680680 582950 680750
rect 583020 680680 583040 680750
rect 583110 680680 583170 680750
rect 135741 645780 136232 680669
rect 580942 680650 583170 680680
rect 119854 645460 136232 645780
rect 137524 678966 146744 679446
rect 137524 639921 138004 678966
rect 119500 639600 138004 639921
rect 93369 638170 95369 638207
rect 93369 638100 94280 638170
rect 94350 638100 94380 638170
rect 94450 638100 94480 638170
rect 94550 638100 95369 638170
rect 93369 638080 95369 638100
rect 93369 638010 94280 638080
rect 94350 638010 94380 638080
rect 94450 638010 94480 638080
rect 94550 638010 95369 638080
rect 93369 635957 95369 638010
rect 97956 638170 99956 638193
rect 97956 638100 98838 638170
rect 98908 638100 98938 638170
rect 99008 638100 99038 638170
rect 99108 638100 99956 638170
rect 97956 638080 99956 638100
rect 97956 638010 98838 638080
rect 98908 638010 98938 638080
rect 99008 638010 99038 638080
rect 99108 638010 99956 638080
rect 97956 635957 99956 638010
rect 213722 597445 218699 604249
rect 159903 592449 218699 597445
rect 159903 585564 164900 592449
rect 167020 585564 213234 585565
rect 213700 585564 218699 592449
rect 159903 583817 218699 585564
rect 159903 580569 218696 583817
rect 159903 576976 164900 580569
rect 213700 576976 218696 580569
rect 159903 571979 218696 576976
rect 159903 559151 164900 571979
rect 213700 559151 218696 571979
rect 154044 554151 218696 559151
<< metal5 >>
rect 165594 701000 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 3000 696000 581000 701000
rect 3000 651000 8000 696000
rect 11000 688000 573000 693000
rect 11000 651000 16000 688000
rect 568000 651000 573000 688000
rect 576000 651000 581000 696000
rect 154044 592379 156710 604249
rect 154044 587379 211748 592379
rect 154044 567737 156710 587379
rect 154044 562737 212204 567737
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use big_cap  big_cap_0
timestamp 1636526374
transform 1 0 105480 0 1 586857
box 60730 -31110 106740 14450
use top  top_0
timestamp 1636213485
transform 1 0 89244 0 1 662150
box -6530 -24030 39650 21850
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
