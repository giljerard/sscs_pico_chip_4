magic
tech sky130A
magscale 1 2
timestamp 1637624949
<< res1p41 >>
rect -143 -52 143 52
<< properties >>
string gencell sky130_fd_pr__res_high_po_1p41
string parameters w 1.410 l 0.50 m 1 nx 1 wmin 1.410 lmin 0.50 rho 319.8 val 140.621 dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 0 wmax 1.410 n_guard 0 hv_guard 0 vias 0 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
