magic
tech sky130A
timestamp 1636213402
<< nwell >>
rect -25 505 180 2030
<< nmos >>
rect -3485 -245 3615 -195
rect -3485 -345 3615 -295
rect -3485 -445 3615 -395
rect -3485 -545 3615 -495
rect -3485 -645 3615 -595
rect -3485 -745 3615 -695
rect -3485 -845 3615 -795
rect -3485 -945 3615 -895
rect -3485 -1045 3615 -995
rect -3485 -1145 3615 -1095
<< ndiff >>
rect -3485 -160 3615 -150
rect -3485 -180 -3470 -160
rect -3450 -180 -3430 -160
rect -3410 -180 -3390 -160
rect -3370 -180 -3350 -160
rect -3330 -180 -3310 -160
rect -3290 -180 -3270 -160
rect -3250 -180 -3230 -160
rect -3210 -180 -3190 -160
rect -3170 -180 -3150 -160
rect -3130 -180 -3110 -160
rect -3090 -180 -3070 -160
rect -3050 -180 -3030 -160
rect -3010 -180 -2990 -160
rect -2970 -180 -2950 -160
rect -2930 -180 -2910 -160
rect -2890 -180 -2870 -160
rect -2850 -180 -2830 -160
rect -2810 -180 -2790 -160
rect -2770 -180 -2750 -160
rect -2730 -180 -2710 -160
rect -2690 -180 -2670 -160
rect -2650 -180 -2630 -160
rect -2610 -180 -2590 -160
rect -2570 -180 -2550 -160
rect -2530 -180 -2510 -160
rect -2490 -180 -2470 -160
rect -2450 -180 -2430 -160
rect -2410 -180 -2390 -160
rect -2370 -180 -2350 -160
rect -2330 -180 -2310 -160
rect -2290 -180 -2270 -160
rect -2250 -180 -2230 -160
rect -2210 -180 -2190 -160
rect -2170 -180 -2150 -160
rect -2130 -180 -2110 -160
rect -2090 -180 -2070 -160
rect -2050 -180 -2030 -160
rect -2010 -180 -1990 -160
rect -1970 -180 -1950 -160
rect -1930 -180 -1910 -160
rect -1890 -180 -1870 -160
rect -1850 -180 -1830 -160
rect -1810 -180 -1790 -160
rect -1770 -180 -1750 -160
rect -1730 -180 -1710 -160
rect -1690 -180 -1670 -160
rect -1650 -180 -1630 -160
rect -1610 -180 -1590 -160
rect -1570 -180 -1550 -160
rect -1530 -180 -1510 -160
rect -1460 -180 -1440 -160
rect -1420 -180 -1400 -160
rect -1380 -180 -1360 -160
rect -1340 -180 -1320 -160
rect -1300 -180 -1280 -160
rect -1260 -180 -1240 -160
rect -1220 -180 -1200 -160
rect -1180 -180 -1160 -160
rect -1140 -180 -1120 -160
rect -1100 -180 -1080 -160
rect -1060 -180 -1040 -160
rect -1020 -180 -1000 -160
rect -980 -180 -960 -160
rect -940 -180 -920 -160
rect -900 -180 -880 -160
rect -860 -180 -840 -160
rect -820 -180 -800 -160
rect -780 -180 -760 -160
rect -740 -180 -720 -160
rect -700 -180 -680 -160
rect -660 -180 -640 -160
rect -620 -180 -600 -160
rect -580 -180 -560 -160
rect -540 -180 -520 -160
rect -500 -180 -480 -160
rect -460 -180 -440 -160
rect -420 -180 -400 -160
rect -380 -180 -360 -160
rect -340 -180 -320 -160
rect -300 -180 -280 -160
rect -260 -180 -230 -160
rect -210 -180 -190 -160
rect -170 -180 -150 -160
rect -130 -180 -110 -160
rect -90 -180 -70 -160
rect -50 -180 -30 -160
rect -10 -180 10 -160
rect 30 -180 50 -160
rect 80 -180 100 -160
rect 120 -180 140 -160
rect 160 -180 180 -160
rect 200 -180 220 -160
rect 240 -180 260 -160
rect 280 -180 300 -160
rect 320 -180 340 -160
rect 360 -180 390 -160
rect 410 -180 430 -160
rect 450 -180 470 -160
rect 490 -180 510 -160
rect 530 -180 550 -160
rect 570 -180 590 -160
rect 610 -180 630 -160
rect 650 -180 670 -160
rect 690 -180 710 -160
rect 730 -180 750 -160
rect 770 -180 790 -160
rect 810 -180 830 -160
rect 850 -180 870 -160
rect 890 -180 910 -160
rect 930 -180 950 -160
rect 970 -180 990 -160
rect 1010 -180 1030 -160
rect 1050 -180 1070 -160
rect 1090 -180 1110 -160
rect 1130 -180 1150 -160
rect 1170 -180 1190 -160
rect 1210 -180 1230 -160
rect 1250 -180 1270 -160
rect 1290 -180 1310 -160
rect 1330 -180 1350 -160
rect 1370 -180 1390 -160
rect 1410 -180 1430 -160
rect 1450 -180 1470 -160
rect 1490 -180 1510 -160
rect 1530 -180 1550 -160
rect 1570 -180 1590 -160
rect 1640 -180 1660 -160
rect 1680 -180 1700 -160
rect 1720 -180 1740 -160
rect 1760 -180 1780 -160
rect 1800 -180 1820 -160
rect 1840 -180 1860 -160
rect 1880 -180 1900 -160
rect 1920 -180 1940 -160
rect 1960 -180 1980 -160
rect 2000 -180 2020 -160
rect 2040 -180 2060 -160
rect 2080 -180 2100 -160
rect 2120 -180 2140 -160
rect 2160 -180 2180 -160
rect 2200 -180 2220 -160
rect 2240 -180 2260 -160
rect 2280 -180 2300 -160
rect 2320 -180 2340 -160
rect 2360 -180 2380 -160
rect 2400 -180 2420 -160
rect 2440 -180 2460 -160
rect 2480 -180 2500 -160
rect 2520 -180 2540 -160
rect 2560 -180 2580 -160
rect 2600 -180 2620 -160
rect 2640 -180 2660 -160
rect 2680 -180 2700 -160
rect 2720 -180 2740 -160
rect 2760 -180 2780 -160
rect 2800 -180 2820 -160
rect 2840 -180 2860 -160
rect 2880 -180 2900 -160
rect 2920 -180 2940 -160
rect 2960 -180 2980 -160
rect 3000 -180 3020 -160
rect 3040 -180 3060 -160
rect 3080 -180 3100 -160
rect 3120 -180 3140 -160
rect 3160 -180 3180 -160
rect 3200 -180 3220 -160
rect 3240 -180 3260 -160
rect 3280 -180 3300 -160
rect 3320 -180 3340 -160
rect 3360 -180 3380 -160
rect 3400 -180 3420 -160
rect 3440 -180 3460 -160
rect 3480 -180 3500 -160
rect 3520 -180 3540 -160
rect 3560 -180 3580 -160
rect 3600 -180 3615 -160
rect -3485 -195 3615 -180
rect -3485 -260 3615 -245
rect -3485 -280 -3470 -260
rect -3450 -280 -3430 -260
rect -3410 -280 -3390 -260
rect -3370 -280 -3350 -260
rect -3330 -280 -3310 -260
rect -3290 -280 -3270 -260
rect -3250 -280 -3230 -260
rect -3210 -280 -3190 -260
rect -3170 -280 -3150 -260
rect -3130 -280 -3110 -260
rect -3090 -280 -3070 -260
rect -3050 -280 -3030 -260
rect -3010 -280 -2990 -260
rect -2970 -280 -2950 -260
rect -2930 -280 -2910 -260
rect -2890 -280 -2870 -260
rect -2850 -280 -2830 -260
rect -2810 -280 -2790 -260
rect -2770 -280 -2750 -260
rect -2730 -280 -2710 -260
rect -2690 -280 -2670 -260
rect -2650 -280 -2630 -260
rect -2610 -280 -2590 -260
rect -2570 -280 -2550 -260
rect -2530 -280 -2510 -260
rect -2490 -280 -2470 -260
rect -2450 -280 -2430 -260
rect -2410 -280 -2390 -260
rect -2370 -280 -2350 -260
rect -2330 -280 -2310 -260
rect -2290 -280 -2270 -260
rect -2250 -280 -2230 -260
rect -2210 -280 -2190 -260
rect -2170 -280 -2150 -260
rect -2130 -280 -2110 -260
rect -2090 -280 -2070 -260
rect -2050 -280 -2030 -260
rect -2010 -280 -1990 -260
rect -1970 -280 -1950 -260
rect -1930 -280 -1910 -260
rect -1890 -280 -1870 -260
rect -1850 -280 -1830 -260
rect -1810 -280 -1790 -260
rect -1770 -280 -1750 -260
rect -1730 -280 -1710 -260
rect -1690 -280 -1670 -260
rect -1650 -280 -1630 -260
rect -1610 -280 -1590 -260
rect -1570 -280 -1550 -260
rect -1530 -280 -1510 -260
rect -1460 -280 -1440 -260
rect -1420 -280 -1400 -260
rect -1380 -280 -1360 -260
rect -1340 -280 -1320 -260
rect -1300 -280 -1280 -260
rect -1260 -280 -1240 -260
rect -1220 -280 -1200 -260
rect -1180 -280 -1160 -260
rect -1140 -280 -1120 -260
rect -1100 -280 -1080 -260
rect -1060 -280 -1040 -260
rect -1020 -280 -1000 -260
rect -980 -280 -960 -260
rect -940 -280 -920 -260
rect -900 -280 -880 -260
rect -860 -280 -840 -260
rect -820 -280 -800 -260
rect -780 -280 -760 -260
rect -740 -280 -720 -260
rect -700 -280 -680 -260
rect -660 -280 -640 -260
rect -620 -280 -600 -260
rect -580 -280 -560 -260
rect -540 -280 -520 -260
rect -500 -280 -480 -260
rect -460 -280 -440 -260
rect -420 -280 -400 -260
rect -380 -280 -360 -260
rect -340 -280 -320 -260
rect -300 -280 -280 -260
rect -260 -280 -230 -260
rect -210 -280 -190 -260
rect -170 -280 -150 -260
rect -130 -280 -110 -260
rect -90 -280 -70 -260
rect -50 -280 -30 -260
rect -10 -280 10 -260
rect 30 -280 50 -260
rect 80 -280 100 -260
rect 120 -280 140 -260
rect 160 -280 180 -260
rect 200 -280 220 -260
rect 240 -280 260 -260
rect 280 -280 300 -260
rect 320 -280 340 -260
rect 360 -280 390 -260
rect 410 -280 430 -260
rect 450 -280 470 -260
rect 490 -280 510 -260
rect 530 -280 550 -260
rect 570 -280 590 -260
rect 610 -280 630 -260
rect 650 -280 670 -260
rect 690 -280 710 -260
rect 730 -280 750 -260
rect 770 -280 790 -260
rect 810 -280 830 -260
rect 850 -280 870 -260
rect 890 -280 910 -260
rect 930 -280 950 -260
rect 970 -280 990 -260
rect 1010 -280 1030 -260
rect 1050 -280 1070 -260
rect 1090 -280 1110 -260
rect 1130 -280 1150 -260
rect 1170 -280 1190 -260
rect 1210 -280 1230 -260
rect 1250 -280 1270 -260
rect 1290 -280 1310 -260
rect 1330 -280 1350 -260
rect 1370 -280 1390 -260
rect 1410 -280 1430 -260
rect 1450 -280 1470 -260
rect 1490 -280 1510 -260
rect 1530 -280 1550 -260
rect 1570 -280 1590 -260
rect 1640 -280 1660 -260
rect 1680 -280 1700 -260
rect 1720 -280 1740 -260
rect 1760 -280 1780 -260
rect 1800 -280 1820 -260
rect 1840 -280 1860 -260
rect 1880 -280 1900 -260
rect 1920 -280 1940 -260
rect 1960 -280 1980 -260
rect 2000 -280 2020 -260
rect 2040 -280 2060 -260
rect 2080 -280 2100 -260
rect 2120 -280 2140 -260
rect 2160 -280 2180 -260
rect 2200 -280 2220 -260
rect 2240 -280 2260 -260
rect 2280 -280 2300 -260
rect 2320 -280 2340 -260
rect 2360 -280 2380 -260
rect 2400 -280 2420 -260
rect 2440 -280 2460 -260
rect 2480 -280 2500 -260
rect 2520 -280 2540 -260
rect 2560 -280 2580 -260
rect 2600 -280 2620 -260
rect 2640 -280 2660 -260
rect 2680 -280 2700 -260
rect 2720 -280 2740 -260
rect 2760 -280 2780 -260
rect 2800 -280 2820 -260
rect 2840 -280 2860 -260
rect 2880 -280 2900 -260
rect 2920 -280 2940 -260
rect 2960 -280 2980 -260
rect 3000 -280 3020 -260
rect 3040 -280 3060 -260
rect 3080 -280 3100 -260
rect 3120 -280 3140 -260
rect 3160 -280 3180 -260
rect 3200 -280 3220 -260
rect 3240 -280 3260 -260
rect 3280 -280 3300 -260
rect 3320 -280 3340 -260
rect 3360 -280 3380 -260
rect 3400 -280 3420 -260
rect 3440 -280 3460 -260
rect 3480 -280 3500 -260
rect 3520 -280 3540 -260
rect 3560 -280 3580 -260
rect 3600 -280 3615 -260
rect -3485 -295 3615 -280
rect -3485 -360 3615 -345
rect -3485 -380 -3470 -360
rect -3450 -380 -3430 -360
rect -3410 -380 -3390 -360
rect -3370 -380 -3350 -360
rect -3330 -380 -3310 -360
rect -3290 -380 -3270 -360
rect -3250 -380 -3230 -360
rect -3210 -380 -3190 -360
rect -3170 -380 -3150 -360
rect -3130 -380 -3110 -360
rect -3090 -380 -3070 -360
rect -3050 -380 -3030 -360
rect -3010 -380 -2990 -360
rect -2970 -380 -2950 -360
rect -2930 -380 -2910 -360
rect -2890 -380 -2870 -360
rect -2850 -380 -2830 -360
rect -2810 -380 -2790 -360
rect -2770 -380 -2750 -360
rect -2730 -380 -2710 -360
rect -2690 -380 -2670 -360
rect -2650 -380 -2630 -360
rect -2610 -380 -2590 -360
rect -2570 -380 -2550 -360
rect -2530 -380 -2510 -360
rect -2490 -380 -2470 -360
rect -2450 -380 -2430 -360
rect -2410 -380 -2390 -360
rect -2370 -380 -2350 -360
rect -2330 -380 -2310 -360
rect -2290 -380 -2270 -360
rect -2250 -380 -2230 -360
rect -2210 -380 -2190 -360
rect -2170 -380 -2150 -360
rect -2130 -380 -2110 -360
rect -2090 -380 -2070 -360
rect -2050 -380 -2030 -360
rect -2010 -380 -1990 -360
rect -1970 -380 -1950 -360
rect -1930 -380 -1910 -360
rect -1890 -380 -1870 -360
rect -1850 -380 -1830 -360
rect -1810 -380 -1790 -360
rect -1770 -380 -1750 -360
rect -1730 -380 -1710 -360
rect -1690 -380 -1670 -360
rect -1650 -380 -1630 -360
rect -1610 -380 -1590 -360
rect -1570 -380 -1550 -360
rect -1530 -380 -1510 -360
rect -1460 -380 -1440 -360
rect -1420 -380 -1400 -360
rect -1380 -380 -1360 -360
rect -1340 -380 -1320 -360
rect -1300 -380 -1280 -360
rect -1260 -380 -1240 -360
rect -1220 -380 -1200 -360
rect -1180 -380 -1160 -360
rect -1140 -380 -1120 -360
rect -1100 -380 -1080 -360
rect -1060 -380 -1040 -360
rect -1020 -380 -1000 -360
rect -980 -380 -960 -360
rect -940 -380 -920 -360
rect -900 -380 -880 -360
rect -860 -380 -840 -360
rect -820 -380 -800 -360
rect -780 -380 -760 -360
rect -740 -380 -720 -360
rect -700 -380 -680 -360
rect -660 -380 -640 -360
rect -620 -380 -600 -360
rect -580 -380 -560 -360
rect -540 -380 -520 -360
rect -500 -380 -480 -360
rect -460 -380 -440 -360
rect -420 -380 -400 -360
rect -380 -380 -360 -360
rect -340 -380 -320 -360
rect -300 -380 -280 -360
rect -260 -380 -230 -360
rect -210 -380 -190 -360
rect -170 -380 -150 -360
rect -130 -380 -110 -360
rect -90 -380 -70 -360
rect -50 -380 -30 -360
rect -10 -380 10 -360
rect 30 -380 50 -360
rect 80 -380 100 -360
rect 120 -380 140 -360
rect 160 -380 180 -360
rect 200 -380 220 -360
rect 240 -380 260 -360
rect 280 -380 300 -360
rect 320 -380 340 -360
rect 360 -380 390 -360
rect 410 -380 430 -360
rect 450 -380 470 -360
rect 490 -380 510 -360
rect 530 -380 550 -360
rect 570 -380 590 -360
rect 610 -380 630 -360
rect 650 -380 670 -360
rect 690 -380 710 -360
rect 730 -380 750 -360
rect 770 -380 790 -360
rect 810 -380 830 -360
rect 850 -380 870 -360
rect 890 -380 910 -360
rect 930 -380 950 -360
rect 970 -380 990 -360
rect 1010 -380 1030 -360
rect 1050 -380 1070 -360
rect 1090 -380 1110 -360
rect 1130 -380 1150 -360
rect 1170 -380 1190 -360
rect 1210 -380 1230 -360
rect 1250 -380 1270 -360
rect 1290 -380 1310 -360
rect 1330 -380 1350 -360
rect 1370 -380 1390 -360
rect 1410 -380 1430 -360
rect 1450 -380 1470 -360
rect 1490 -380 1510 -360
rect 1530 -380 1550 -360
rect 1570 -380 1590 -360
rect 1640 -380 1660 -360
rect 1680 -380 1700 -360
rect 1720 -380 1740 -360
rect 1760 -380 1780 -360
rect 1800 -380 1820 -360
rect 1840 -380 1860 -360
rect 1880 -380 1900 -360
rect 1920 -380 1940 -360
rect 1960 -380 1980 -360
rect 2000 -380 2020 -360
rect 2040 -380 2060 -360
rect 2080 -380 2100 -360
rect 2120 -380 2140 -360
rect 2160 -380 2180 -360
rect 2200 -380 2220 -360
rect 2240 -380 2260 -360
rect 2280 -380 2300 -360
rect 2320 -380 2340 -360
rect 2360 -380 2380 -360
rect 2400 -380 2420 -360
rect 2440 -380 2460 -360
rect 2480 -380 2500 -360
rect 2520 -380 2540 -360
rect 2560 -380 2580 -360
rect 2600 -380 2620 -360
rect 2640 -380 2660 -360
rect 2680 -380 2700 -360
rect 2720 -380 2740 -360
rect 2760 -380 2780 -360
rect 2800 -380 2820 -360
rect 2840 -380 2860 -360
rect 2880 -380 2900 -360
rect 2920 -380 2940 -360
rect 2960 -380 2980 -360
rect 3000 -380 3020 -360
rect 3040 -380 3060 -360
rect 3080 -380 3100 -360
rect 3120 -380 3140 -360
rect 3160 -380 3180 -360
rect 3200 -380 3220 -360
rect 3240 -380 3260 -360
rect 3280 -380 3300 -360
rect 3320 -380 3340 -360
rect 3360 -380 3380 -360
rect 3400 -380 3420 -360
rect 3440 -380 3460 -360
rect 3480 -380 3500 -360
rect 3520 -380 3540 -360
rect 3560 -380 3580 -360
rect 3600 -380 3615 -360
rect -3485 -395 3615 -380
rect -3485 -460 3615 -445
rect -3485 -480 -3470 -460
rect -3450 -480 -3430 -460
rect -3410 -480 -3390 -460
rect -3370 -480 -3350 -460
rect -3330 -480 -3310 -460
rect -3290 -480 -3270 -460
rect -3250 -480 -3230 -460
rect -3210 -480 -3190 -460
rect -3170 -480 -3150 -460
rect -3130 -480 -3110 -460
rect -3090 -480 -3070 -460
rect -3050 -480 -3030 -460
rect -3010 -480 -2990 -460
rect -2970 -480 -2950 -460
rect -2930 -480 -2910 -460
rect -2890 -480 -2870 -460
rect -2850 -480 -2830 -460
rect -2810 -480 -2790 -460
rect -2770 -480 -2750 -460
rect -2730 -480 -2710 -460
rect -2690 -480 -2670 -460
rect -2650 -480 -2630 -460
rect -2610 -480 -2590 -460
rect -2570 -480 -2550 -460
rect -2530 -480 -2510 -460
rect -2490 -480 -2470 -460
rect -2450 -480 -2430 -460
rect -2410 -480 -2390 -460
rect -2370 -480 -2350 -460
rect -2330 -480 -2310 -460
rect -2290 -480 -2270 -460
rect -2250 -480 -2230 -460
rect -2210 -480 -2190 -460
rect -2170 -480 -2150 -460
rect -2130 -480 -2110 -460
rect -2090 -480 -2070 -460
rect -2050 -480 -2030 -460
rect -2010 -480 -1990 -460
rect -1970 -480 -1950 -460
rect -1930 -480 -1910 -460
rect -1890 -480 -1870 -460
rect -1850 -480 -1830 -460
rect -1810 -480 -1790 -460
rect -1770 -480 -1750 -460
rect -1730 -480 -1710 -460
rect -1690 -480 -1670 -460
rect -1650 -480 -1630 -460
rect -1610 -480 -1590 -460
rect -1570 -480 -1550 -460
rect -1530 -480 -1510 -460
rect -1460 -480 -1440 -460
rect -1420 -480 -1400 -460
rect -1380 -480 -1360 -460
rect -1340 -480 -1320 -460
rect -1300 -480 -1280 -460
rect -1260 -480 -1240 -460
rect -1220 -480 -1200 -460
rect -1180 -480 -1160 -460
rect -1140 -480 -1120 -460
rect -1100 -480 -1080 -460
rect -1060 -480 -1040 -460
rect -1020 -480 -1000 -460
rect -980 -480 -960 -460
rect -940 -480 -920 -460
rect -900 -480 -880 -460
rect -860 -480 -840 -460
rect -820 -480 -800 -460
rect -780 -480 -760 -460
rect -740 -480 -720 -460
rect -700 -480 -680 -460
rect -660 -480 -640 -460
rect -620 -480 -600 -460
rect -580 -480 -560 -460
rect -540 -480 -520 -460
rect -500 -480 -480 -460
rect -460 -480 -440 -460
rect -420 -480 -400 -460
rect -380 -480 -360 -460
rect -340 -480 -320 -460
rect -300 -480 -280 -460
rect -260 -480 -230 -460
rect -210 -480 -190 -460
rect -170 -480 -150 -460
rect -130 -480 -110 -460
rect -90 -480 -70 -460
rect -50 -480 -30 -460
rect -10 -480 10 -460
rect 30 -480 50 -460
rect 80 -480 100 -460
rect 120 -480 140 -460
rect 160 -480 180 -460
rect 200 -480 220 -460
rect 240 -480 260 -460
rect 280 -480 300 -460
rect 320 -480 340 -460
rect 360 -480 390 -460
rect 410 -480 430 -460
rect 450 -480 470 -460
rect 490 -480 510 -460
rect 530 -480 550 -460
rect 570 -480 590 -460
rect 610 -480 630 -460
rect 650 -480 670 -460
rect 690 -480 710 -460
rect 730 -480 750 -460
rect 770 -480 790 -460
rect 810 -480 830 -460
rect 850 -480 870 -460
rect 890 -480 910 -460
rect 930 -480 950 -460
rect 970 -480 990 -460
rect 1010 -480 1030 -460
rect 1050 -480 1070 -460
rect 1090 -480 1110 -460
rect 1130 -480 1150 -460
rect 1170 -480 1190 -460
rect 1210 -480 1230 -460
rect 1250 -480 1270 -460
rect 1290 -480 1310 -460
rect 1330 -480 1350 -460
rect 1370 -480 1390 -460
rect 1410 -480 1430 -460
rect 1450 -480 1470 -460
rect 1490 -480 1510 -460
rect 1530 -480 1550 -460
rect 1570 -480 1590 -460
rect 1640 -480 1660 -460
rect 1680 -480 1700 -460
rect 1720 -480 1740 -460
rect 1760 -480 1780 -460
rect 1800 -480 1820 -460
rect 1840 -480 1860 -460
rect 1880 -480 1900 -460
rect 1920 -480 1940 -460
rect 1960 -480 1980 -460
rect 2000 -480 2020 -460
rect 2040 -480 2060 -460
rect 2080 -480 2100 -460
rect 2120 -480 2140 -460
rect 2160 -480 2180 -460
rect 2200 -480 2220 -460
rect 2240 -480 2260 -460
rect 2280 -480 2300 -460
rect 2320 -480 2340 -460
rect 2360 -480 2380 -460
rect 2400 -480 2420 -460
rect 2440 -480 2460 -460
rect 2480 -480 2500 -460
rect 2520 -480 2540 -460
rect 2560 -480 2580 -460
rect 2600 -480 2620 -460
rect 2640 -480 2660 -460
rect 2680 -480 2700 -460
rect 2720 -480 2740 -460
rect 2760 -480 2780 -460
rect 2800 -480 2820 -460
rect 2840 -480 2860 -460
rect 2880 -480 2900 -460
rect 2920 -480 2940 -460
rect 2960 -480 2980 -460
rect 3000 -480 3020 -460
rect 3040 -480 3060 -460
rect 3080 -480 3100 -460
rect 3120 -480 3140 -460
rect 3160 -480 3180 -460
rect 3200 -480 3220 -460
rect 3240 -480 3260 -460
rect 3280 -480 3300 -460
rect 3320 -480 3340 -460
rect 3360 -480 3380 -460
rect 3400 -480 3420 -460
rect 3440 -480 3460 -460
rect 3480 -480 3500 -460
rect 3520 -480 3540 -460
rect 3560 -480 3580 -460
rect 3600 -480 3615 -460
rect -3485 -495 3615 -480
rect -3485 -560 3615 -545
rect -3485 -580 -3470 -560
rect -3450 -580 -3430 -560
rect -3410 -580 -3390 -560
rect -3370 -580 -3350 -560
rect -3330 -580 -3310 -560
rect -3290 -580 -3270 -560
rect -3250 -580 -3230 -560
rect -3210 -580 -3190 -560
rect -3170 -580 -3150 -560
rect -3130 -580 -3110 -560
rect -3090 -580 -3070 -560
rect -3050 -580 -3030 -560
rect -3010 -580 -2990 -560
rect -2970 -580 -2950 -560
rect -2930 -580 -2910 -560
rect -2890 -580 -2870 -560
rect -2850 -580 -2830 -560
rect -2810 -580 -2790 -560
rect -2770 -580 -2750 -560
rect -2730 -580 -2710 -560
rect -2690 -580 -2670 -560
rect -2650 -580 -2630 -560
rect -2610 -580 -2590 -560
rect -2570 -580 -2550 -560
rect -2530 -580 -2510 -560
rect -2490 -580 -2470 -560
rect -2450 -580 -2430 -560
rect -2410 -580 -2390 -560
rect -2370 -580 -2350 -560
rect -2330 -580 -2310 -560
rect -2290 -580 -2270 -560
rect -2250 -580 -2230 -560
rect -2210 -580 -2190 -560
rect -2170 -580 -2150 -560
rect -2130 -580 -2110 -560
rect -2090 -580 -2070 -560
rect -2050 -580 -2030 -560
rect -2010 -580 -1990 -560
rect -1970 -580 -1950 -560
rect -1930 -580 -1910 -560
rect -1890 -580 -1870 -560
rect -1850 -580 -1830 -560
rect -1810 -580 -1790 -560
rect -1770 -580 -1750 -560
rect -1730 -580 -1710 -560
rect -1690 -580 -1670 -560
rect -1650 -580 -1630 -560
rect -1610 -580 -1590 -560
rect -1570 -580 -1550 -560
rect -1530 -580 -1510 -560
rect -1460 -580 -1440 -560
rect -1420 -580 -1400 -560
rect -1380 -580 -1360 -560
rect -1340 -580 -1320 -560
rect -1300 -580 -1280 -560
rect -1260 -580 -1240 -560
rect -1220 -580 -1200 -560
rect -1180 -580 -1160 -560
rect -1140 -580 -1120 -560
rect -1100 -580 -1080 -560
rect -1060 -580 -1040 -560
rect -1020 -580 -1000 -560
rect -980 -580 -960 -560
rect -940 -580 -920 -560
rect -900 -580 -880 -560
rect -860 -580 -840 -560
rect -820 -580 -800 -560
rect -780 -580 -760 -560
rect -740 -580 -720 -560
rect -700 -580 -680 -560
rect -660 -580 -640 -560
rect -620 -580 -600 -560
rect -580 -580 -560 -560
rect -540 -580 -520 -560
rect -500 -580 -480 -560
rect -460 -580 -440 -560
rect -420 -580 -400 -560
rect -380 -580 -360 -560
rect -340 -580 -320 -560
rect -300 -580 -280 -560
rect -260 -580 -230 -560
rect -210 -580 -190 -560
rect -170 -580 -150 -560
rect -130 -580 -110 -560
rect -90 -580 -70 -560
rect -50 -580 -30 -560
rect -10 -580 10 -560
rect 30 -580 50 -560
rect 80 -580 100 -560
rect 120 -580 140 -560
rect 160 -580 180 -560
rect 200 -580 220 -560
rect 240 -580 260 -560
rect 280 -580 300 -560
rect 320 -580 340 -560
rect 360 -580 390 -560
rect 410 -580 430 -560
rect 450 -580 470 -560
rect 490 -580 510 -560
rect 530 -580 550 -560
rect 570 -580 590 -560
rect 610 -580 630 -560
rect 650 -580 670 -560
rect 690 -580 710 -560
rect 730 -580 750 -560
rect 770 -580 790 -560
rect 810 -580 830 -560
rect 850 -580 870 -560
rect 890 -580 910 -560
rect 930 -580 950 -560
rect 970 -580 990 -560
rect 1010 -580 1030 -560
rect 1050 -580 1070 -560
rect 1090 -580 1110 -560
rect 1130 -580 1150 -560
rect 1170 -580 1190 -560
rect 1210 -580 1230 -560
rect 1250 -580 1270 -560
rect 1290 -580 1310 -560
rect 1330 -580 1350 -560
rect 1370 -580 1390 -560
rect 1410 -580 1430 -560
rect 1450 -580 1470 -560
rect 1490 -580 1510 -560
rect 1530 -580 1550 -560
rect 1570 -580 1590 -560
rect 1640 -580 1660 -560
rect 1680 -580 1700 -560
rect 1720 -580 1740 -560
rect 1760 -580 1780 -560
rect 1800 -580 1820 -560
rect 1840 -580 1860 -560
rect 1880 -580 1900 -560
rect 1920 -580 1940 -560
rect 1960 -580 1980 -560
rect 2000 -580 2020 -560
rect 2040 -580 2060 -560
rect 2080 -580 2100 -560
rect 2120 -580 2140 -560
rect 2160 -580 2180 -560
rect 2200 -580 2220 -560
rect 2240 -580 2260 -560
rect 2280 -580 2300 -560
rect 2320 -580 2340 -560
rect 2360 -580 2380 -560
rect 2400 -580 2420 -560
rect 2440 -580 2460 -560
rect 2480 -580 2500 -560
rect 2520 -580 2540 -560
rect 2560 -580 2580 -560
rect 2600 -580 2620 -560
rect 2640 -580 2660 -560
rect 2680 -580 2700 -560
rect 2720 -580 2740 -560
rect 2760 -580 2780 -560
rect 2800 -580 2820 -560
rect 2840 -580 2860 -560
rect 2880 -580 2900 -560
rect 2920 -580 2940 -560
rect 2960 -580 2980 -560
rect 3000 -580 3020 -560
rect 3040 -580 3060 -560
rect 3080 -580 3100 -560
rect 3120 -580 3140 -560
rect 3160 -580 3180 -560
rect 3200 -580 3220 -560
rect 3240 -580 3260 -560
rect 3280 -580 3300 -560
rect 3320 -580 3340 -560
rect 3360 -580 3380 -560
rect 3400 -580 3420 -560
rect 3440 -580 3460 -560
rect 3480 -580 3500 -560
rect 3520 -580 3540 -560
rect 3560 -580 3580 -560
rect 3600 -580 3615 -560
rect -3485 -595 3615 -580
rect -3485 -660 3615 -645
rect -3485 -680 -3470 -660
rect -3450 -680 -3430 -660
rect -3410 -680 -3390 -660
rect -3370 -680 -3350 -660
rect -3330 -680 -3310 -660
rect -3290 -680 -3270 -660
rect -3250 -680 -3230 -660
rect -3210 -680 -3190 -660
rect -3170 -680 -3150 -660
rect -3130 -680 -3110 -660
rect -3090 -680 -3070 -660
rect -3050 -680 -3030 -660
rect -3010 -680 -2990 -660
rect -2970 -680 -2950 -660
rect -2930 -680 -2910 -660
rect -2890 -680 -2870 -660
rect -2850 -680 -2830 -660
rect -2810 -680 -2790 -660
rect -2770 -680 -2750 -660
rect -2730 -680 -2710 -660
rect -2690 -680 -2670 -660
rect -2650 -680 -2630 -660
rect -2610 -680 -2590 -660
rect -2570 -680 -2550 -660
rect -2530 -680 -2510 -660
rect -2490 -680 -2470 -660
rect -2450 -680 -2430 -660
rect -2410 -680 -2390 -660
rect -2370 -680 -2350 -660
rect -2330 -680 -2310 -660
rect -2290 -680 -2270 -660
rect -2250 -680 -2230 -660
rect -2210 -680 -2190 -660
rect -2170 -680 -2150 -660
rect -2130 -680 -2110 -660
rect -2090 -680 -2070 -660
rect -2050 -680 -2030 -660
rect -2010 -680 -1990 -660
rect -1970 -680 -1950 -660
rect -1930 -680 -1910 -660
rect -1890 -680 -1870 -660
rect -1850 -680 -1830 -660
rect -1810 -680 -1790 -660
rect -1770 -680 -1750 -660
rect -1730 -680 -1710 -660
rect -1690 -680 -1670 -660
rect -1650 -680 -1630 -660
rect -1610 -680 -1590 -660
rect -1570 -680 -1550 -660
rect -1530 -680 -1510 -660
rect -1460 -680 -1440 -660
rect -1420 -680 -1400 -660
rect -1380 -680 -1360 -660
rect -1340 -680 -1320 -660
rect -1300 -680 -1280 -660
rect -1260 -680 -1240 -660
rect -1220 -680 -1200 -660
rect -1180 -680 -1160 -660
rect -1140 -680 -1120 -660
rect -1100 -680 -1080 -660
rect -1060 -680 -1040 -660
rect -1020 -680 -1000 -660
rect -980 -680 -960 -660
rect -940 -680 -920 -660
rect -900 -680 -880 -660
rect -860 -680 -840 -660
rect -820 -680 -800 -660
rect -780 -680 -760 -660
rect -740 -680 -720 -660
rect -700 -680 -680 -660
rect -660 -680 -640 -660
rect -620 -680 -600 -660
rect -580 -680 -560 -660
rect -540 -680 -520 -660
rect -500 -680 -480 -660
rect -460 -680 -440 -660
rect -420 -680 -400 -660
rect -380 -680 -360 -660
rect -340 -680 -320 -660
rect -300 -680 -280 -660
rect -260 -680 -230 -660
rect -210 -680 -190 -660
rect -170 -680 -150 -660
rect -130 -680 -110 -660
rect -90 -680 -70 -660
rect -50 -680 -30 -660
rect -10 -680 10 -660
rect 30 -680 50 -660
rect 80 -680 100 -660
rect 120 -680 140 -660
rect 160 -680 180 -660
rect 200 -680 220 -660
rect 240 -680 260 -660
rect 280 -680 300 -660
rect 320 -680 340 -660
rect 360 -680 390 -660
rect 410 -680 430 -660
rect 450 -680 470 -660
rect 490 -680 510 -660
rect 530 -680 550 -660
rect 570 -680 590 -660
rect 610 -680 630 -660
rect 650 -680 670 -660
rect 690 -680 710 -660
rect 730 -680 750 -660
rect 770 -680 790 -660
rect 810 -680 830 -660
rect 850 -680 870 -660
rect 890 -680 910 -660
rect 930 -680 950 -660
rect 970 -680 990 -660
rect 1010 -680 1030 -660
rect 1050 -680 1070 -660
rect 1090 -680 1110 -660
rect 1130 -680 1150 -660
rect 1170 -680 1190 -660
rect 1210 -680 1230 -660
rect 1250 -680 1270 -660
rect 1290 -680 1310 -660
rect 1330 -680 1350 -660
rect 1370 -680 1390 -660
rect 1410 -680 1430 -660
rect 1450 -680 1470 -660
rect 1490 -680 1510 -660
rect 1530 -680 1550 -660
rect 1570 -680 1590 -660
rect 1640 -680 1660 -660
rect 1680 -680 1700 -660
rect 1720 -680 1740 -660
rect 1760 -680 1780 -660
rect 1800 -680 1820 -660
rect 1840 -680 1860 -660
rect 1880 -680 1900 -660
rect 1920 -680 1940 -660
rect 1960 -680 1980 -660
rect 2000 -680 2020 -660
rect 2040 -680 2060 -660
rect 2080 -680 2100 -660
rect 2120 -680 2140 -660
rect 2160 -680 2180 -660
rect 2200 -680 2220 -660
rect 2240 -680 2260 -660
rect 2280 -680 2300 -660
rect 2320 -680 2340 -660
rect 2360 -680 2380 -660
rect 2400 -680 2420 -660
rect 2440 -680 2460 -660
rect 2480 -680 2500 -660
rect 2520 -680 2540 -660
rect 2560 -680 2580 -660
rect 2600 -680 2620 -660
rect 2640 -680 2660 -660
rect 2680 -680 2700 -660
rect 2720 -680 2740 -660
rect 2760 -680 2780 -660
rect 2800 -680 2820 -660
rect 2840 -680 2860 -660
rect 2880 -680 2900 -660
rect 2920 -680 2940 -660
rect 2960 -680 2980 -660
rect 3000 -680 3020 -660
rect 3040 -680 3060 -660
rect 3080 -680 3100 -660
rect 3120 -680 3140 -660
rect 3160 -680 3180 -660
rect 3200 -680 3220 -660
rect 3240 -680 3260 -660
rect 3280 -680 3300 -660
rect 3320 -680 3340 -660
rect 3360 -680 3380 -660
rect 3400 -680 3420 -660
rect 3440 -680 3460 -660
rect 3480 -680 3500 -660
rect 3520 -680 3540 -660
rect 3560 -680 3580 -660
rect 3600 -680 3615 -660
rect -3485 -695 3615 -680
rect -3485 -760 3615 -745
rect -3485 -780 -3470 -760
rect -3450 -780 -3430 -760
rect -3410 -780 -3390 -760
rect -3370 -780 -3350 -760
rect -3330 -780 -3310 -760
rect -3290 -780 -3270 -760
rect -3250 -780 -3230 -760
rect -3210 -780 -3190 -760
rect -3170 -780 -3150 -760
rect -3130 -780 -3110 -760
rect -3090 -780 -3070 -760
rect -3050 -780 -3030 -760
rect -3010 -780 -2990 -760
rect -2970 -780 -2950 -760
rect -2930 -780 -2910 -760
rect -2890 -780 -2870 -760
rect -2850 -780 -2830 -760
rect -2810 -780 -2790 -760
rect -2770 -780 -2750 -760
rect -2730 -780 -2710 -760
rect -2690 -780 -2670 -760
rect -2650 -780 -2630 -760
rect -2610 -780 -2590 -760
rect -2570 -780 -2550 -760
rect -2530 -780 -2510 -760
rect -2490 -780 -2470 -760
rect -2450 -780 -2430 -760
rect -2410 -780 -2390 -760
rect -2370 -780 -2350 -760
rect -2330 -780 -2310 -760
rect -2290 -780 -2270 -760
rect -2250 -780 -2230 -760
rect -2210 -780 -2190 -760
rect -2170 -780 -2150 -760
rect -2130 -780 -2110 -760
rect -2090 -780 -2070 -760
rect -2050 -780 -2030 -760
rect -2010 -780 -1990 -760
rect -1970 -780 -1950 -760
rect -1930 -780 -1910 -760
rect -1890 -780 -1870 -760
rect -1850 -780 -1830 -760
rect -1810 -780 -1790 -760
rect -1770 -780 -1750 -760
rect -1730 -780 -1710 -760
rect -1690 -780 -1670 -760
rect -1650 -780 -1630 -760
rect -1610 -780 -1590 -760
rect -1570 -780 -1550 -760
rect -1530 -780 -1510 -760
rect -1460 -780 -1440 -760
rect -1420 -780 -1400 -760
rect -1380 -780 -1360 -760
rect -1340 -780 -1320 -760
rect -1300 -780 -1280 -760
rect -1260 -780 -1240 -760
rect -1220 -780 -1200 -760
rect -1180 -780 -1160 -760
rect -1140 -780 -1120 -760
rect -1100 -780 -1080 -760
rect -1060 -780 -1040 -760
rect -1020 -780 -1000 -760
rect -980 -780 -960 -760
rect -940 -780 -920 -760
rect -900 -780 -880 -760
rect -860 -780 -840 -760
rect -820 -780 -800 -760
rect -780 -780 -760 -760
rect -740 -780 -720 -760
rect -700 -780 -680 -760
rect -660 -780 -640 -760
rect -620 -780 -600 -760
rect -580 -780 -560 -760
rect -540 -780 -520 -760
rect -500 -780 -480 -760
rect -460 -780 -440 -760
rect -420 -780 -400 -760
rect -380 -780 -360 -760
rect -340 -780 -320 -760
rect -300 -780 -280 -760
rect -260 -780 -230 -760
rect -210 -780 -190 -760
rect -170 -780 -150 -760
rect -130 -780 -110 -760
rect -90 -780 -70 -760
rect -50 -780 -30 -760
rect -10 -780 10 -760
rect 30 -780 50 -760
rect 80 -780 100 -760
rect 120 -780 140 -760
rect 160 -780 180 -760
rect 200 -780 220 -760
rect 240 -780 260 -760
rect 280 -780 300 -760
rect 320 -780 340 -760
rect 360 -780 390 -760
rect 410 -780 430 -760
rect 450 -780 470 -760
rect 490 -780 510 -760
rect 530 -780 550 -760
rect 570 -780 590 -760
rect 610 -780 630 -760
rect 650 -780 670 -760
rect 690 -780 710 -760
rect 730 -780 750 -760
rect 770 -780 790 -760
rect 810 -780 830 -760
rect 850 -780 870 -760
rect 890 -780 910 -760
rect 930 -780 950 -760
rect 970 -780 990 -760
rect 1010 -780 1030 -760
rect 1050 -780 1070 -760
rect 1090 -780 1110 -760
rect 1130 -780 1150 -760
rect 1170 -780 1190 -760
rect 1210 -780 1230 -760
rect 1250 -780 1270 -760
rect 1290 -780 1310 -760
rect 1330 -780 1350 -760
rect 1370 -780 1390 -760
rect 1410 -780 1430 -760
rect 1450 -780 1470 -760
rect 1490 -780 1510 -760
rect 1530 -780 1550 -760
rect 1570 -780 1590 -760
rect 1640 -780 1660 -760
rect 1680 -780 1700 -760
rect 1720 -780 1740 -760
rect 1760 -780 1780 -760
rect 1800 -780 1820 -760
rect 1840 -780 1860 -760
rect 1880 -780 1900 -760
rect 1920 -780 1940 -760
rect 1960 -780 1980 -760
rect 2000 -780 2020 -760
rect 2040 -780 2060 -760
rect 2080 -780 2100 -760
rect 2120 -780 2140 -760
rect 2160 -780 2180 -760
rect 2200 -780 2220 -760
rect 2240 -780 2260 -760
rect 2280 -780 2300 -760
rect 2320 -780 2340 -760
rect 2360 -780 2380 -760
rect 2400 -780 2420 -760
rect 2440 -780 2460 -760
rect 2480 -780 2500 -760
rect 2520 -780 2540 -760
rect 2560 -780 2580 -760
rect 2600 -780 2620 -760
rect 2640 -780 2660 -760
rect 2680 -780 2700 -760
rect 2720 -780 2740 -760
rect 2760 -780 2780 -760
rect 2800 -780 2820 -760
rect 2840 -780 2860 -760
rect 2880 -780 2900 -760
rect 2920 -780 2940 -760
rect 2960 -780 2980 -760
rect 3000 -780 3020 -760
rect 3040 -780 3060 -760
rect 3080 -780 3100 -760
rect 3120 -780 3140 -760
rect 3160 -780 3180 -760
rect 3200 -780 3220 -760
rect 3240 -780 3260 -760
rect 3280 -780 3300 -760
rect 3320 -780 3340 -760
rect 3360 -780 3380 -760
rect 3400 -780 3420 -760
rect 3440 -780 3460 -760
rect 3480 -780 3500 -760
rect 3520 -780 3540 -760
rect 3560 -780 3580 -760
rect 3600 -780 3615 -760
rect -3485 -795 3615 -780
rect -3485 -860 3615 -845
rect -3485 -880 -3470 -860
rect -3450 -880 -3430 -860
rect -3410 -880 -3390 -860
rect -3370 -880 -3350 -860
rect -3330 -880 -3310 -860
rect -3290 -880 -3270 -860
rect -3250 -880 -3230 -860
rect -3210 -880 -3190 -860
rect -3170 -880 -3150 -860
rect -3130 -880 -3110 -860
rect -3090 -880 -3070 -860
rect -3050 -880 -3030 -860
rect -3010 -880 -2990 -860
rect -2970 -880 -2950 -860
rect -2930 -880 -2910 -860
rect -2890 -880 -2870 -860
rect -2850 -880 -2830 -860
rect -2810 -880 -2790 -860
rect -2770 -880 -2750 -860
rect -2730 -880 -2710 -860
rect -2690 -880 -2670 -860
rect -2650 -880 -2630 -860
rect -2610 -880 -2590 -860
rect -2570 -880 -2550 -860
rect -2530 -880 -2510 -860
rect -2490 -880 -2470 -860
rect -2450 -880 -2430 -860
rect -2410 -880 -2390 -860
rect -2370 -880 -2350 -860
rect -2330 -880 -2310 -860
rect -2290 -880 -2270 -860
rect -2250 -880 -2230 -860
rect -2210 -880 -2190 -860
rect -2170 -880 -2150 -860
rect -2130 -880 -2110 -860
rect -2090 -880 -2070 -860
rect -2050 -880 -2030 -860
rect -2010 -880 -1990 -860
rect -1970 -880 -1950 -860
rect -1930 -880 -1910 -860
rect -1890 -880 -1870 -860
rect -1850 -880 -1830 -860
rect -1810 -880 -1790 -860
rect -1770 -880 -1750 -860
rect -1730 -880 -1710 -860
rect -1690 -880 -1670 -860
rect -1650 -880 -1630 -860
rect -1610 -880 -1590 -860
rect -1570 -880 -1550 -860
rect -1530 -880 -1510 -860
rect -1460 -880 -1440 -860
rect -1420 -880 -1400 -860
rect -1380 -880 -1360 -860
rect -1340 -880 -1320 -860
rect -1300 -880 -1280 -860
rect -1260 -880 -1240 -860
rect -1220 -880 -1200 -860
rect -1180 -880 -1160 -860
rect -1140 -880 -1120 -860
rect -1100 -880 -1080 -860
rect -1060 -880 -1040 -860
rect -1020 -880 -1000 -860
rect -980 -880 -960 -860
rect -940 -880 -920 -860
rect -900 -880 -880 -860
rect -860 -880 -840 -860
rect -820 -880 -800 -860
rect -780 -880 -760 -860
rect -740 -880 -720 -860
rect -700 -880 -680 -860
rect -660 -880 -640 -860
rect -620 -880 -600 -860
rect -580 -880 -560 -860
rect -540 -880 -520 -860
rect -500 -880 -480 -860
rect -460 -880 -440 -860
rect -420 -880 -400 -860
rect -380 -880 -360 -860
rect -340 -880 -320 -860
rect -300 -880 -280 -860
rect -260 -880 -230 -860
rect -210 -880 -190 -860
rect -170 -880 -150 -860
rect -130 -880 -110 -860
rect -90 -880 -70 -860
rect -50 -880 -30 -860
rect -10 -880 10 -860
rect 30 -880 50 -860
rect 80 -880 100 -860
rect 120 -880 140 -860
rect 160 -880 180 -860
rect 200 -880 220 -860
rect 240 -880 260 -860
rect 280 -880 300 -860
rect 320 -880 340 -860
rect 360 -880 390 -860
rect 410 -880 430 -860
rect 450 -880 470 -860
rect 490 -880 510 -860
rect 530 -880 550 -860
rect 570 -880 590 -860
rect 610 -880 630 -860
rect 650 -880 670 -860
rect 690 -880 710 -860
rect 730 -880 750 -860
rect 770 -880 790 -860
rect 810 -880 830 -860
rect 850 -880 870 -860
rect 890 -880 910 -860
rect 930 -880 950 -860
rect 970 -880 990 -860
rect 1010 -880 1030 -860
rect 1050 -880 1070 -860
rect 1090 -880 1110 -860
rect 1130 -880 1150 -860
rect 1170 -880 1190 -860
rect 1210 -880 1230 -860
rect 1250 -880 1270 -860
rect 1290 -880 1310 -860
rect 1330 -880 1350 -860
rect 1370 -880 1390 -860
rect 1410 -880 1430 -860
rect 1450 -880 1470 -860
rect 1490 -880 1510 -860
rect 1530 -880 1550 -860
rect 1570 -880 1590 -860
rect 1640 -880 1660 -860
rect 1680 -880 1700 -860
rect 1720 -880 1740 -860
rect 1760 -880 1780 -860
rect 1800 -880 1820 -860
rect 1840 -880 1860 -860
rect 1880 -880 1900 -860
rect 1920 -880 1940 -860
rect 1960 -880 1980 -860
rect 2000 -880 2020 -860
rect 2040 -880 2060 -860
rect 2080 -880 2100 -860
rect 2120 -880 2140 -860
rect 2160 -880 2180 -860
rect 2200 -880 2220 -860
rect 2240 -880 2260 -860
rect 2280 -880 2300 -860
rect 2320 -880 2340 -860
rect 2360 -880 2380 -860
rect 2400 -880 2420 -860
rect 2440 -880 2460 -860
rect 2480 -880 2500 -860
rect 2520 -880 2540 -860
rect 2560 -880 2580 -860
rect 2600 -880 2620 -860
rect 2640 -880 2660 -860
rect 2680 -880 2700 -860
rect 2720 -880 2740 -860
rect 2760 -880 2780 -860
rect 2800 -880 2820 -860
rect 2840 -880 2860 -860
rect 2880 -880 2900 -860
rect 2920 -880 2940 -860
rect 2960 -880 2980 -860
rect 3000 -880 3020 -860
rect 3040 -880 3060 -860
rect 3080 -880 3100 -860
rect 3120 -880 3140 -860
rect 3160 -880 3180 -860
rect 3200 -880 3220 -860
rect 3240 -880 3260 -860
rect 3280 -880 3300 -860
rect 3320 -880 3340 -860
rect 3360 -880 3380 -860
rect 3400 -880 3420 -860
rect 3440 -880 3460 -860
rect 3480 -880 3500 -860
rect 3520 -880 3540 -860
rect 3560 -880 3580 -860
rect 3600 -880 3615 -860
rect -3485 -895 3615 -880
rect -3485 -960 3615 -945
rect -3485 -980 -3470 -960
rect -3450 -980 -3430 -960
rect -3410 -980 -3390 -960
rect -3370 -980 -3350 -960
rect -3330 -980 -3310 -960
rect -3290 -980 -3270 -960
rect -3250 -980 -3230 -960
rect -3210 -980 -3190 -960
rect -3170 -980 -3150 -960
rect -3130 -980 -3110 -960
rect -3090 -980 -3070 -960
rect -3050 -980 -3030 -960
rect -3010 -980 -2990 -960
rect -2970 -980 -2950 -960
rect -2930 -980 -2910 -960
rect -2890 -980 -2870 -960
rect -2850 -980 -2830 -960
rect -2810 -980 -2790 -960
rect -2770 -980 -2750 -960
rect -2730 -980 -2710 -960
rect -2690 -980 -2670 -960
rect -2650 -980 -2630 -960
rect -2610 -980 -2590 -960
rect -2570 -980 -2550 -960
rect -2530 -980 -2510 -960
rect -2490 -980 -2470 -960
rect -2450 -980 -2430 -960
rect -2410 -980 -2390 -960
rect -2370 -980 -2350 -960
rect -2330 -980 -2310 -960
rect -2290 -980 -2270 -960
rect -2250 -980 -2230 -960
rect -2210 -980 -2190 -960
rect -2170 -980 -2150 -960
rect -2130 -980 -2110 -960
rect -2090 -980 -2070 -960
rect -2050 -980 -2030 -960
rect -2010 -980 -1990 -960
rect -1970 -980 -1950 -960
rect -1930 -980 -1910 -960
rect -1890 -980 -1870 -960
rect -1850 -980 -1830 -960
rect -1810 -980 -1790 -960
rect -1770 -980 -1750 -960
rect -1730 -980 -1710 -960
rect -1690 -980 -1670 -960
rect -1650 -980 -1630 -960
rect -1610 -980 -1590 -960
rect -1570 -980 -1550 -960
rect -1530 -980 -1510 -960
rect -1460 -980 -1440 -960
rect -1420 -980 -1400 -960
rect -1380 -980 -1360 -960
rect -1340 -980 -1320 -960
rect -1300 -980 -1280 -960
rect -1260 -980 -1240 -960
rect -1220 -980 -1200 -960
rect -1180 -980 -1160 -960
rect -1140 -980 -1120 -960
rect -1100 -980 -1080 -960
rect -1060 -980 -1040 -960
rect -1020 -980 -1000 -960
rect -980 -980 -960 -960
rect -940 -980 -920 -960
rect -900 -980 -880 -960
rect -860 -980 -840 -960
rect -820 -980 -800 -960
rect -780 -980 -760 -960
rect -740 -980 -720 -960
rect -700 -980 -680 -960
rect -660 -980 -640 -960
rect -620 -980 -600 -960
rect -580 -980 -560 -960
rect -540 -980 -520 -960
rect -500 -980 -480 -960
rect -460 -980 -440 -960
rect -420 -980 -400 -960
rect -380 -980 -360 -960
rect -340 -980 -320 -960
rect -300 -980 -280 -960
rect -260 -980 -230 -960
rect -210 -980 -190 -960
rect -170 -980 -150 -960
rect -130 -980 -110 -960
rect -90 -980 -70 -960
rect -50 -980 -30 -960
rect -10 -980 10 -960
rect 30 -980 50 -960
rect 80 -980 100 -960
rect 120 -980 140 -960
rect 160 -980 180 -960
rect 200 -980 220 -960
rect 240 -980 260 -960
rect 280 -980 300 -960
rect 320 -980 340 -960
rect 360 -980 390 -960
rect 410 -980 430 -960
rect 450 -980 470 -960
rect 490 -980 510 -960
rect 530 -980 550 -960
rect 570 -980 590 -960
rect 610 -980 630 -960
rect 650 -980 670 -960
rect 690 -980 710 -960
rect 730 -980 750 -960
rect 770 -980 790 -960
rect 810 -980 830 -960
rect 850 -980 870 -960
rect 890 -980 910 -960
rect 930 -980 950 -960
rect 970 -980 990 -960
rect 1010 -980 1030 -960
rect 1050 -980 1070 -960
rect 1090 -980 1110 -960
rect 1130 -980 1150 -960
rect 1170 -980 1190 -960
rect 1210 -980 1230 -960
rect 1250 -980 1270 -960
rect 1290 -980 1310 -960
rect 1330 -980 1350 -960
rect 1370 -980 1390 -960
rect 1410 -980 1430 -960
rect 1450 -980 1470 -960
rect 1490 -980 1510 -960
rect 1530 -980 1550 -960
rect 1570 -980 1590 -960
rect 1640 -980 1660 -960
rect 1680 -980 1700 -960
rect 1720 -980 1740 -960
rect 1760 -980 1780 -960
rect 1800 -980 1820 -960
rect 1840 -980 1860 -960
rect 1880 -980 1900 -960
rect 1920 -980 1940 -960
rect 1960 -980 1980 -960
rect 2000 -980 2020 -960
rect 2040 -980 2060 -960
rect 2080 -980 2100 -960
rect 2120 -980 2140 -960
rect 2160 -980 2180 -960
rect 2200 -980 2220 -960
rect 2240 -980 2260 -960
rect 2280 -980 2300 -960
rect 2320 -980 2340 -960
rect 2360 -980 2380 -960
rect 2400 -980 2420 -960
rect 2440 -980 2460 -960
rect 2480 -980 2500 -960
rect 2520 -980 2540 -960
rect 2560 -980 2580 -960
rect 2600 -980 2620 -960
rect 2640 -980 2660 -960
rect 2680 -980 2700 -960
rect 2720 -980 2740 -960
rect 2760 -980 2780 -960
rect 2800 -980 2820 -960
rect 2840 -980 2860 -960
rect 2880 -980 2900 -960
rect 2920 -980 2940 -960
rect 2960 -980 2980 -960
rect 3000 -980 3020 -960
rect 3040 -980 3060 -960
rect 3080 -980 3100 -960
rect 3120 -980 3140 -960
rect 3160 -980 3180 -960
rect 3200 -980 3220 -960
rect 3240 -980 3260 -960
rect 3280 -980 3300 -960
rect 3320 -980 3340 -960
rect 3360 -980 3380 -960
rect 3400 -980 3420 -960
rect 3440 -980 3460 -960
rect 3480 -980 3500 -960
rect 3520 -980 3540 -960
rect 3560 -980 3580 -960
rect 3600 -980 3615 -960
rect -3485 -995 3615 -980
rect -3485 -1060 3615 -1045
rect -3485 -1080 -3470 -1060
rect -3450 -1080 -3430 -1060
rect -3410 -1080 -3390 -1060
rect -3370 -1080 -3350 -1060
rect -3330 -1080 -3310 -1060
rect -3290 -1080 -3270 -1060
rect -3250 -1080 -3230 -1060
rect -3210 -1080 -3190 -1060
rect -3170 -1080 -3150 -1060
rect -3130 -1080 -3110 -1060
rect -3090 -1080 -3070 -1060
rect -3050 -1080 -3030 -1060
rect -3010 -1080 -2990 -1060
rect -2970 -1080 -2950 -1060
rect -2930 -1080 -2910 -1060
rect -2890 -1080 -2870 -1060
rect -2850 -1080 -2830 -1060
rect -2810 -1080 -2790 -1060
rect -2770 -1080 -2750 -1060
rect -2730 -1080 -2710 -1060
rect -2690 -1080 -2670 -1060
rect -2650 -1080 -2630 -1060
rect -2610 -1080 -2590 -1060
rect -2570 -1080 -2550 -1060
rect -2530 -1080 -2510 -1060
rect -2490 -1080 -2470 -1060
rect -2450 -1080 -2430 -1060
rect -2410 -1080 -2390 -1060
rect -2370 -1080 -2350 -1060
rect -2330 -1080 -2310 -1060
rect -2290 -1080 -2270 -1060
rect -2250 -1080 -2230 -1060
rect -2210 -1080 -2190 -1060
rect -2170 -1080 -2150 -1060
rect -2130 -1080 -2110 -1060
rect -2090 -1080 -2070 -1060
rect -2050 -1080 -2030 -1060
rect -2010 -1080 -1990 -1060
rect -1970 -1080 -1950 -1060
rect -1930 -1080 -1910 -1060
rect -1890 -1080 -1870 -1060
rect -1850 -1080 -1830 -1060
rect -1810 -1080 -1790 -1060
rect -1770 -1080 -1750 -1060
rect -1730 -1080 -1710 -1060
rect -1690 -1080 -1670 -1060
rect -1650 -1080 -1630 -1060
rect -1610 -1080 -1590 -1060
rect -1570 -1080 -1550 -1060
rect -1530 -1080 -1510 -1060
rect -1460 -1080 -1440 -1060
rect -1420 -1080 -1400 -1060
rect -1380 -1080 -1360 -1060
rect -1340 -1080 -1320 -1060
rect -1300 -1080 -1280 -1060
rect -1260 -1080 -1240 -1060
rect -1220 -1080 -1200 -1060
rect -1180 -1080 -1160 -1060
rect -1140 -1080 -1120 -1060
rect -1100 -1080 -1080 -1060
rect -1060 -1080 -1040 -1060
rect -1020 -1080 -1000 -1060
rect -980 -1080 -960 -1060
rect -940 -1080 -920 -1060
rect -900 -1080 -880 -1060
rect -860 -1080 -840 -1060
rect -820 -1080 -800 -1060
rect -780 -1080 -760 -1060
rect -740 -1080 -720 -1060
rect -700 -1080 -680 -1060
rect -660 -1080 -640 -1060
rect -620 -1080 -600 -1060
rect -580 -1080 -560 -1060
rect -540 -1080 -520 -1060
rect -500 -1080 -480 -1060
rect -460 -1080 -440 -1060
rect -420 -1080 -400 -1060
rect -380 -1080 -360 -1060
rect -340 -1080 -320 -1060
rect -300 -1080 -280 -1060
rect -260 -1080 -230 -1060
rect -210 -1080 -190 -1060
rect -170 -1080 -150 -1060
rect -130 -1080 -110 -1060
rect -90 -1080 -70 -1060
rect -50 -1080 -30 -1060
rect -10 -1080 10 -1060
rect 30 -1080 50 -1060
rect 80 -1080 100 -1060
rect 120 -1080 140 -1060
rect 160 -1080 180 -1060
rect 200 -1080 220 -1060
rect 240 -1080 260 -1060
rect 280 -1080 300 -1060
rect 320 -1080 340 -1060
rect 360 -1080 390 -1060
rect 410 -1080 430 -1060
rect 450 -1080 470 -1060
rect 490 -1080 510 -1060
rect 530 -1080 550 -1060
rect 570 -1080 590 -1060
rect 610 -1080 630 -1060
rect 650 -1080 670 -1060
rect 690 -1080 710 -1060
rect 730 -1080 750 -1060
rect 770 -1080 790 -1060
rect 810 -1080 830 -1060
rect 850 -1080 870 -1060
rect 890 -1080 910 -1060
rect 930 -1080 950 -1060
rect 970 -1080 990 -1060
rect 1010 -1080 1030 -1060
rect 1050 -1080 1070 -1060
rect 1090 -1080 1110 -1060
rect 1130 -1080 1150 -1060
rect 1170 -1080 1190 -1060
rect 1210 -1080 1230 -1060
rect 1250 -1080 1270 -1060
rect 1290 -1080 1310 -1060
rect 1330 -1080 1350 -1060
rect 1370 -1080 1390 -1060
rect 1410 -1080 1430 -1060
rect 1450 -1080 1470 -1060
rect 1490 -1080 1510 -1060
rect 1530 -1080 1550 -1060
rect 1570 -1080 1590 -1060
rect 1640 -1080 1660 -1060
rect 1680 -1080 1700 -1060
rect 1720 -1080 1740 -1060
rect 1760 -1080 1780 -1060
rect 1800 -1080 1820 -1060
rect 1840 -1080 1860 -1060
rect 1880 -1080 1900 -1060
rect 1920 -1080 1940 -1060
rect 1960 -1080 1980 -1060
rect 2000 -1080 2020 -1060
rect 2040 -1080 2060 -1060
rect 2080 -1080 2100 -1060
rect 2120 -1080 2140 -1060
rect 2160 -1080 2180 -1060
rect 2200 -1080 2220 -1060
rect 2240 -1080 2260 -1060
rect 2280 -1080 2300 -1060
rect 2320 -1080 2340 -1060
rect 2360 -1080 2380 -1060
rect 2400 -1080 2420 -1060
rect 2440 -1080 2460 -1060
rect 2480 -1080 2500 -1060
rect 2520 -1080 2540 -1060
rect 2560 -1080 2580 -1060
rect 2600 -1080 2620 -1060
rect 2640 -1080 2660 -1060
rect 2680 -1080 2700 -1060
rect 2720 -1080 2740 -1060
rect 2760 -1080 2780 -1060
rect 2800 -1080 2820 -1060
rect 2840 -1080 2860 -1060
rect 2880 -1080 2900 -1060
rect 2920 -1080 2940 -1060
rect 2960 -1080 2980 -1060
rect 3000 -1080 3020 -1060
rect 3040 -1080 3060 -1060
rect 3080 -1080 3100 -1060
rect 3120 -1080 3140 -1060
rect 3160 -1080 3180 -1060
rect 3200 -1080 3220 -1060
rect 3240 -1080 3260 -1060
rect 3280 -1080 3300 -1060
rect 3320 -1080 3340 -1060
rect 3360 -1080 3380 -1060
rect 3400 -1080 3420 -1060
rect 3440 -1080 3460 -1060
rect 3480 -1080 3500 -1060
rect 3520 -1080 3540 -1060
rect 3560 -1080 3580 -1060
rect 3600 -1080 3615 -1060
rect -3485 -1095 3615 -1080
rect -3485 -1160 3615 -1145
rect -3485 -1180 -3470 -1160
rect -3450 -1180 -3430 -1160
rect -3410 -1180 -3390 -1160
rect -3370 -1180 -3350 -1160
rect -3330 -1180 -3310 -1160
rect -3290 -1180 -3270 -1160
rect -3250 -1180 -3230 -1160
rect -3210 -1180 -3190 -1160
rect -3170 -1180 -3150 -1160
rect -3130 -1180 -3110 -1160
rect -3090 -1180 -3070 -1160
rect -3050 -1180 -3030 -1160
rect -3010 -1180 -2990 -1160
rect -2970 -1180 -2950 -1160
rect -2930 -1180 -2910 -1160
rect -2890 -1180 -2870 -1160
rect -2850 -1180 -2830 -1160
rect -2810 -1180 -2790 -1160
rect -2770 -1180 -2750 -1160
rect -2730 -1180 -2710 -1160
rect -2690 -1180 -2670 -1160
rect -2650 -1180 -2630 -1160
rect -2610 -1180 -2590 -1160
rect -2570 -1180 -2550 -1160
rect -2530 -1180 -2510 -1160
rect -2490 -1180 -2470 -1160
rect -2450 -1180 -2430 -1160
rect -2410 -1180 -2390 -1160
rect -2370 -1180 -2350 -1160
rect -2330 -1180 -2310 -1160
rect -2290 -1180 -2270 -1160
rect -2250 -1180 -2230 -1160
rect -2210 -1180 -2190 -1160
rect -2170 -1180 -2150 -1160
rect -2130 -1180 -2110 -1160
rect -2090 -1180 -2070 -1160
rect -2050 -1180 -2030 -1160
rect -2010 -1180 -1990 -1160
rect -1970 -1180 -1950 -1160
rect -1930 -1180 -1910 -1160
rect -1890 -1180 -1870 -1160
rect -1850 -1180 -1830 -1160
rect -1810 -1180 -1790 -1160
rect -1770 -1180 -1750 -1160
rect -1730 -1180 -1710 -1160
rect -1690 -1180 -1670 -1160
rect -1650 -1180 -1630 -1160
rect -1610 -1180 -1590 -1160
rect -1570 -1180 -1550 -1160
rect -1530 -1180 -1510 -1160
rect -1490 -1180 -1470 -1160
rect -1450 -1180 -1430 -1160
rect -1410 -1180 -1390 -1160
rect -1370 -1180 -1350 -1160
rect -1330 -1180 -1310 -1160
rect -1290 -1180 -1270 -1160
rect -1250 -1180 -1230 -1160
rect -1210 -1180 -1190 -1160
rect -1170 -1180 -1150 -1160
rect -1130 -1180 -1110 -1160
rect -1090 -1180 -1070 -1160
rect -1050 -1180 -1030 -1160
rect -1010 -1180 -990 -1160
rect -970 -1180 -950 -1160
rect -930 -1180 -910 -1160
rect -890 -1180 -870 -1160
rect -850 -1180 -830 -1160
rect -810 -1180 -790 -1160
rect -770 -1180 -750 -1160
rect -730 -1180 -710 -1160
rect -690 -1180 -670 -1160
rect -650 -1180 -630 -1160
rect -610 -1180 -590 -1160
rect -570 -1180 -550 -1160
rect -530 -1180 -510 -1160
rect -490 -1180 -470 -1160
rect -450 -1180 -430 -1160
rect -410 -1180 -390 -1160
rect -370 -1180 -350 -1160
rect -330 -1180 -310 -1160
rect -290 -1180 -270 -1160
rect -250 -1180 -230 -1160
rect -210 -1180 -190 -1160
rect -170 -1180 -150 -1160
rect -130 -1180 -110 -1160
rect -90 -1180 -70 -1160
rect -50 -1180 -30 -1160
rect -10 -1180 10 -1160
rect 30 -1180 50 -1160
rect 80 -1180 100 -1160
rect 120 -1180 140 -1160
rect 160 -1180 180 -1160
rect 200 -1180 220 -1160
rect 240 -1180 260 -1160
rect 280 -1180 300 -1160
rect 320 -1180 340 -1160
rect 360 -1180 380 -1160
rect 400 -1180 420 -1160
rect 440 -1180 460 -1160
rect 480 -1180 500 -1160
rect 520 -1180 540 -1160
rect 560 -1180 580 -1160
rect 600 -1180 620 -1160
rect 640 -1180 660 -1160
rect 680 -1180 700 -1160
rect 720 -1180 740 -1160
rect 760 -1180 780 -1160
rect 800 -1180 820 -1160
rect 840 -1180 860 -1160
rect 880 -1180 900 -1160
rect 920 -1180 940 -1160
rect 960 -1180 980 -1160
rect 1000 -1180 1020 -1160
rect 1040 -1180 1060 -1160
rect 1080 -1180 1100 -1160
rect 1120 -1180 1140 -1160
rect 1160 -1180 1180 -1160
rect 1200 -1180 1220 -1160
rect 1240 -1180 1260 -1160
rect 1280 -1180 1300 -1160
rect 1320 -1180 1340 -1160
rect 1360 -1180 1380 -1160
rect 1400 -1180 1420 -1160
rect 1440 -1180 1460 -1160
rect 1480 -1180 1500 -1160
rect 1520 -1180 1540 -1160
rect 1560 -1180 1580 -1160
rect 1600 -1180 1620 -1160
rect 1640 -1180 1660 -1160
rect 1680 -1180 1700 -1160
rect 1720 -1180 1740 -1160
rect 1760 -1180 1780 -1160
rect 1800 -1180 1820 -1160
rect 1840 -1180 1860 -1160
rect 1880 -1180 1900 -1160
rect 1920 -1180 1940 -1160
rect 1960 -1180 1980 -1160
rect 2000 -1180 2020 -1160
rect 2040 -1180 2060 -1160
rect 2080 -1180 2100 -1160
rect 2120 -1180 2140 -1160
rect 2160 -1180 2180 -1160
rect 2200 -1180 2220 -1160
rect 2240 -1180 2260 -1160
rect 2280 -1180 2300 -1160
rect 2320 -1180 2340 -1160
rect 2360 -1180 2380 -1160
rect 2400 -1180 2420 -1160
rect 2440 -1180 2460 -1160
rect 2480 -1180 2500 -1160
rect 2520 -1180 2540 -1160
rect 2560 -1180 2580 -1160
rect 2600 -1180 2620 -1160
rect 2640 -1180 2660 -1160
rect 2680 -1180 2700 -1160
rect 2720 -1180 2740 -1160
rect 2760 -1180 2780 -1160
rect 2800 -1180 2820 -1160
rect 2840 -1180 2860 -1160
rect 2880 -1180 2900 -1160
rect 2920 -1180 2940 -1160
rect 2960 -1180 2980 -1160
rect 3000 -1180 3020 -1160
rect 3040 -1180 3060 -1160
rect 3080 -1180 3100 -1160
rect 3120 -1180 3140 -1160
rect 3160 -1180 3180 -1160
rect 3200 -1180 3220 -1160
rect 3240 -1180 3260 -1160
rect 3280 -1180 3300 -1160
rect 3320 -1180 3340 -1160
rect 3360 -1180 3380 -1160
rect 3400 -1180 3420 -1160
rect 3440 -1180 3460 -1160
rect 3480 -1180 3500 -1160
rect 3520 -1180 3540 -1160
rect 3560 -1180 3580 -1160
rect 3600 -1180 3615 -1160
rect -3485 -1190 3615 -1180
<< ndiffc >>
rect -3470 -180 -3450 -160
rect -3430 -180 -3410 -160
rect -3390 -180 -3370 -160
rect -3350 -180 -3330 -160
rect -3310 -180 -3290 -160
rect -3270 -180 -3250 -160
rect -3230 -180 -3210 -160
rect -3190 -180 -3170 -160
rect -3150 -180 -3130 -160
rect -3110 -180 -3090 -160
rect -3070 -180 -3050 -160
rect -3030 -180 -3010 -160
rect -2990 -180 -2970 -160
rect -2950 -180 -2930 -160
rect -2910 -180 -2890 -160
rect -2870 -180 -2850 -160
rect -2830 -180 -2810 -160
rect -2790 -180 -2770 -160
rect -2750 -180 -2730 -160
rect -2710 -180 -2690 -160
rect -2670 -180 -2650 -160
rect -2630 -180 -2610 -160
rect -2590 -180 -2570 -160
rect -2550 -180 -2530 -160
rect -2510 -180 -2490 -160
rect -2470 -180 -2450 -160
rect -2430 -180 -2410 -160
rect -2390 -180 -2370 -160
rect -2350 -180 -2330 -160
rect -2310 -180 -2290 -160
rect -2270 -180 -2250 -160
rect -2230 -180 -2210 -160
rect -2190 -180 -2170 -160
rect -2150 -180 -2130 -160
rect -2110 -180 -2090 -160
rect -2070 -180 -2050 -160
rect -2030 -180 -2010 -160
rect -1990 -180 -1970 -160
rect -1950 -180 -1930 -160
rect -1910 -180 -1890 -160
rect -1870 -180 -1850 -160
rect -1830 -180 -1810 -160
rect -1790 -180 -1770 -160
rect -1750 -180 -1730 -160
rect -1710 -180 -1690 -160
rect -1670 -180 -1650 -160
rect -1630 -180 -1610 -160
rect -1590 -180 -1570 -160
rect -1550 -180 -1530 -160
rect -1510 -180 -1460 -160
rect -1440 -180 -1420 -160
rect -1400 -180 -1380 -160
rect -1360 -180 -1340 -160
rect -1320 -180 -1300 -160
rect -1280 -180 -1260 -160
rect -1240 -180 -1220 -160
rect -1200 -180 -1180 -160
rect -1160 -180 -1140 -160
rect -1120 -180 -1100 -160
rect -1080 -180 -1060 -160
rect -1040 -180 -1020 -160
rect -1000 -180 -980 -160
rect -960 -180 -940 -160
rect -920 -180 -900 -160
rect -880 -180 -860 -160
rect -840 -180 -820 -160
rect -800 -180 -780 -160
rect -760 -180 -740 -160
rect -720 -180 -700 -160
rect -680 -180 -660 -160
rect -640 -180 -620 -160
rect -600 -180 -580 -160
rect -560 -180 -540 -160
rect -520 -180 -500 -160
rect -480 -180 -460 -160
rect -440 -180 -420 -160
rect -400 -180 -380 -160
rect -360 -180 -340 -160
rect -320 -180 -300 -160
rect -280 -180 -260 -160
rect -230 -180 -210 -160
rect -190 -180 -170 -160
rect -150 -180 -130 -160
rect -110 -180 -90 -160
rect -70 -180 -50 -160
rect -30 -180 -10 -160
rect 10 -180 30 -160
rect 50 -180 80 -160
rect 100 -180 120 -160
rect 140 -180 160 -160
rect 180 -180 200 -160
rect 220 -180 240 -160
rect 260 -180 280 -160
rect 300 -180 320 -160
rect 340 -180 360 -160
rect 390 -180 410 -160
rect 430 -180 450 -160
rect 470 -180 490 -160
rect 510 -180 530 -160
rect 550 -180 570 -160
rect 590 -180 610 -160
rect 630 -180 650 -160
rect 670 -180 690 -160
rect 710 -180 730 -160
rect 750 -180 770 -160
rect 790 -180 810 -160
rect 830 -180 850 -160
rect 870 -180 890 -160
rect 910 -180 930 -160
rect 950 -180 970 -160
rect 990 -180 1010 -160
rect 1030 -180 1050 -160
rect 1070 -180 1090 -160
rect 1110 -180 1130 -160
rect 1150 -180 1170 -160
rect 1190 -180 1210 -160
rect 1230 -180 1250 -160
rect 1270 -180 1290 -160
rect 1310 -180 1330 -160
rect 1350 -180 1370 -160
rect 1390 -180 1410 -160
rect 1430 -180 1450 -160
rect 1470 -180 1490 -160
rect 1510 -180 1530 -160
rect 1550 -180 1570 -160
rect 1590 -180 1640 -160
rect 1660 -180 1680 -160
rect 1700 -180 1720 -160
rect 1740 -180 1760 -160
rect 1780 -180 1800 -160
rect 1820 -180 1840 -160
rect 1860 -180 1880 -160
rect 1900 -180 1920 -160
rect 1940 -180 1960 -160
rect 1980 -180 2000 -160
rect 2020 -180 2040 -160
rect 2060 -180 2080 -160
rect 2100 -180 2120 -160
rect 2140 -180 2160 -160
rect 2180 -180 2200 -160
rect 2220 -180 2240 -160
rect 2260 -180 2280 -160
rect 2300 -180 2320 -160
rect 2340 -180 2360 -160
rect 2380 -180 2400 -160
rect 2420 -180 2440 -160
rect 2460 -180 2480 -160
rect 2500 -180 2520 -160
rect 2540 -180 2560 -160
rect 2580 -180 2600 -160
rect 2620 -180 2640 -160
rect 2660 -180 2680 -160
rect 2700 -180 2720 -160
rect 2740 -180 2760 -160
rect 2780 -180 2800 -160
rect 2820 -180 2840 -160
rect 2860 -180 2880 -160
rect 2900 -180 2920 -160
rect 2940 -180 2960 -160
rect 2980 -180 3000 -160
rect 3020 -180 3040 -160
rect 3060 -180 3080 -160
rect 3100 -180 3120 -160
rect 3140 -180 3160 -160
rect 3180 -180 3200 -160
rect 3220 -180 3240 -160
rect 3260 -180 3280 -160
rect 3300 -180 3320 -160
rect 3340 -180 3360 -160
rect 3380 -180 3400 -160
rect 3420 -180 3440 -160
rect 3460 -180 3480 -160
rect 3500 -180 3520 -160
rect 3540 -180 3560 -160
rect 3580 -180 3600 -160
rect -3470 -280 -3450 -260
rect -3430 -280 -3410 -260
rect -3390 -280 -3370 -260
rect -3350 -280 -3330 -260
rect -3310 -280 -3290 -260
rect -3270 -280 -3250 -260
rect -3230 -280 -3210 -260
rect -3190 -280 -3170 -260
rect -3150 -280 -3130 -260
rect -3110 -280 -3090 -260
rect -3070 -280 -3050 -260
rect -3030 -280 -3010 -260
rect -2990 -280 -2970 -260
rect -2950 -280 -2930 -260
rect -2910 -280 -2890 -260
rect -2870 -280 -2850 -260
rect -2830 -280 -2810 -260
rect -2790 -280 -2770 -260
rect -2750 -280 -2730 -260
rect -2710 -280 -2690 -260
rect -2670 -280 -2650 -260
rect -2630 -280 -2610 -260
rect -2590 -280 -2570 -260
rect -2550 -280 -2530 -260
rect -2510 -280 -2490 -260
rect -2470 -280 -2450 -260
rect -2430 -280 -2410 -260
rect -2390 -280 -2370 -260
rect -2350 -280 -2330 -260
rect -2310 -280 -2290 -260
rect -2270 -280 -2250 -260
rect -2230 -280 -2210 -260
rect -2190 -280 -2170 -260
rect -2150 -280 -2130 -260
rect -2110 -280 -2090 -260
rect -2070 -280 -2050 -260
rect -2030 -280 -2010 -260
rect -1990 -280 -1970 -260
rect -1950 -280 -1930 -260
rect -1910 -280 -1890 -260
rect -1870 -280 -1850 -260
rect -1830 -280 -1810 -260
rect -1790 -280 -1770 -260
rect -1750 -280 -1730 -260
rect -1710 -280 -1690 -260
rect -1670 -280 -1650 -260
rect -1630 -280 -1610 -260
rect -1590 -280 -1570 -260
rect -1550 -280 -1530 -260
rect -1510 -280 -1460 -260
rect -1440 -280 -1420 -260
rect -1400 -280 -1380 -260
rect -1360 -280 -1340 -260
rect -1320 -280 -1300 -260
rect -1280 -280 -1260 -260
rect -1240 -280 -1220 -260
rect -1200 -280 -1180 -260
rect -1160 -280 -1140 -260
rect -1120 -280 -1100 -260
rect -1080 -280 -1060 -260
rect -1040 -280 -1020 -260
rect -1000 -280 -980 -260
rect -960 -280 -940 -260
rect -920 -280 -900 -260
rect -880 -280 -860 -260
rect -840 -280 -820 -260
rect -800 -280 -780 -260
rect -760 -280 -740 -260
rect -720 -280 -700 -260
rect -680 -280 -660 -260
rect -640 -280 -620 -260
rect -600 -280 -580 -260
rect -560 -280 -540 -260
rect -520 -280 -500 -260
rect -480 -280 -460 -260
rect -440 -280 -420 -260
rect -400 -280 -380 -260
rect -360 -280 -340 -260
rect -320 -280 -300 -260
rect -280 -280 -260 -260
rect -230 -280 -210 -260
rect -190 -280 -170 -260
rect -150 -280 -130 -260
rect -110 -280 -90 -260
rect -70 -280 -50 -260
rect -30 -280 -10 -260
rect 10 -280 30 -260
rect 50 -280 80 -260
rect 100 -280 120 -260
rect 140 -280 160 -260
rect 180 -280 200 -260
rect 220 -280 240 -260
rect 260 -280 280 -260
rect 300 -280 320 -260
rect 340 -280 360 -260
rect 390 -280 410 -260
rect 430 -280 450 -260
rect 470 -280 490 -260
rect 510 -280 530 -260
rect 550 -280 570 -260
rect 590 -280 610 -260
rect 630 -280 650 -260
rect 670 -280 690 -260
rect 710 -280 730 -260
rect 750 -280 770 -260
rect 790 -280 810 -260
rect 830 -280 850 -260
rect 870 -280 890 -260
rect 910 -280 930 -260
rect 950 -280 970 -260
rect 990 -280 1010 -260
rect 1030 -280 1050 -260
rect 1070 -280 1090 -260
rect 1110 -280 1130 -260
rect 1150 -280 1170 -260
rect 1190 -280 1210 -260
rect 1230 -280 1250 -260
rect 1270 -280 1290 -260
rect 1310 -280 1330 -260
rect 1350 -280 1370 -260
rect 1390 -280 1410 -260
rect 1430 -280 1450 -260
rect 1470 -280 1490 -260
rect 1510 -280 1530 -260
rect 1550 -280 1570 -260
rect 1590 -280 1640 -260
rect 1660 -280 1680 -260
rect 1700 -280 1720 -260
rect 1740 -280 1760 -260
rect 1780 -280 1800 -260
rect 1820 -280 1840 -260
rect 1860 -280 1880 -260
rect 1900 -280 1920 -260
rect 1940 -280 1960 -260
rect 1980 -280 2000 -260
rect 2020 -280 2040 -260
rect 2060 -280 2080 -260
rect 2100 -280 2120 -260
rect 2140 -280 2160 -260
rect 2180 -280 2200 -260
rect 2220 -280 2240 -260
rect 2260 -280 2280 -260
rect 2300 -280 2320 -260
rect 2340 -280 2360 -260
rect 2380 -280 2400 -260
rect 2420 -280 2440 -260
rect 2460 -280 2480 -260
rect 2500 -280 2520 -260
rect 2540 -280 2560 -260
rect 2580 -280 2600 -260
rect 2620 -280 2640 -260
rect 2660 -280 2680 -260
rect 2700 -280 2720 -260
rect 2740 -280 2760 -260
rect 2780 -280 2800 -260
rect 2820 -280 2840 -260
rect 2860 -280 2880 -260
rect 2900 -280 2920 -260
rect 2940 -280 2960 -260
rect 2980 -280 3000 -260
rect 3020 -280 3040 -260
rect 3060 -280 3080 -260
rect 3100 -280 3120 -260
rect 3140 -280 3160 -260
rect 3180 -280 3200 -260
rect 3220 -280 3240 -260
rect 3260 -280 3280 -260
rect 3300 -280 3320 -260
rect 3340 -280 3360 -260
rect 3380 -280 3400 -260
rect 3420 -280 3440 -260
rect 3460 -280 3480 -260
rect 3500 -280 3520 -260
rect 3540 -280 3560 -260
rect 3580 -280 3600 -260
rect -3470 -380 -3450 -360
rect -3430 -380 -3410 -360
rect -3390 -380 -3370 -360
rect -3350 -380 -3330 -360
rect -3310 -380 -3290 -360
rect -3270 -380 -3250 -360
rect -3230 -380 -3210 -360
rect -3190 -380 -3170 -360
rect -3150 -380 -3130 -360
rect -3110 -380 -3090 -360
rect -3070 -380 -3050 -360
rect -3030 -380 -3010 -360
rect -2990 -380 -2970 -360
rect -2950 -380 -2930 -360
rect -2910 -380 -2890 -360
rect -2870 -380 -2850 -360
rect -2830 -380 -2810 -360
rect -2790 -380 -2770 -360
rect -2750 -380 -2730 -360
rect -2710 -380 -2690 -360
rect -2670 -380 -2650 -360
rect -2630 -380 -2610 -360
rect -2590 -380 -2570 -360
rect -2550 -380 -2530 -360
rect -2510 -380 -2490 -360
rect -2470 -380 -2450 -360
rect -2430 -380 -2410 -360
rect -2390 -380 -2370 -360
rect -2350 -380 -2330 -360
rect -2310 -380 -2290 -360
rect -2270 -380 -2250 -360
rect -2230 -380 -2210 -360
rect -2190 -380 -2170 -360
rect -2150 -380 -2130 -360
rect -2110 -380 -2090 -360
rect -2070 -380 -2050 -360
rect -2030 -380 -2010 -360
rect -1990 -380 -1970 -360
rect -1950 -380 -1930 -360
rect -1910 -380 -1890 -360
rect -1870 -380 -1850 -360
rect -1830 -380 -1810 -360
rect -1790 -380 -1770 -360
rect -1750 -380 -1730 -360
rect -1710 -380 -1690 -360
rect -1670 -380 -1650 -360
rect -1630 -380 -1610 -360
rect -1590 -380 -1570 -360
rect -1550 -380 -1530 -360
rect -1510 -380 -1460 -360
rect -1440 -380 -1420 -360
rect -1400 -380 -1380 -360
rect -1360 -380 -1340 -360
rect -1320 -380 -1300 -360
rect -1280 -380 -1260 -360
rect -1240 -380 -1220 -360
rect -1200 -380 -1180 -360
rect -1160 -380 -1140 -360
rect -1120 -380 -1100 -360
rect -1080 -380 -1060 -360
rect -1040 -380 -1020 -360
rect -1000 -380 -980 -360
rect -960 -380 -940 -360
rect -920 -380 -900 -360
rect -880 -380 -860 -360
rect -840 -380 -820 -360
rect -800 -380 -780 -360
rect -760 -380 -740 -360
rect -720 -380 -700 -360
rect -680 -380 -660 -360
rect -640 -380 -620 -360
rect -600 -380 -580 -360
rect -560 -380 -540 -360
rect -520 -380 -500 -360
rect -480 -380 -460 -360
rect -440 -380 -420 -360
rect -400 -380 -380 -360
rect -360 -380 -340 -360
rect -320 -380 -300 -360
rect -280 -380 -260 -360
rect -230 -380 -210 -360
rect -190 -380 -170 -360
rect -150 -380 -130 -360
rect -110 -380 -90 -360
rect -70 -380 -50 -360
rect -30 -380 -10 -360
rect 10 -380 30 -360
rect 50 -380 80 -360
rect 100 -380 120 -360
rect 140 -380 160 -360
rect 180 -380 200 -360
rect 220 -380 240 -360
rect 260 -380 280 -360
rect 300 -380 320 -360
rect 340 -380 360 -360
rect 390 -380 410 -360
rect 430 -380 450 -360
rect 470 -380 490 -360
rect 510 -380 530 -360
rect 550 -380 570 -360
rect 590 -380 610 -360
rect 630 -380 650 -360
rect 670 -380 690 -360
rect 710 -380 730 -360
rect 750 -380 770 -360
rect 790 -380 810 -360
rect 830 -380 850 -360
rect 870 -380 890 -360
rect 910 -380 930 -360
rect 950 -380 970 -360
rect 990 -380 1010 -360
rect 1030 -380 1050 -360
rect 1070 -380 1090 -360
rect 1110 -380 1130 -360
rect 1150 -380 1170 -360
rect 1190 -380 1210 -360
rect 1230 -380 1250 -360
rect 1270 -380 1290 -360
rect 1310 -380 1330 -360
rect 1350 -380 1370 -360
rect 1390 -380 1410 -360
rect 1430 -380 1450 -360
rect 1470 -380 1490 -360
rect 1510 -380 1530 -360
rect 1550 -380 1570 -360
rect 1590 -380 1640 -360
rect 1660 -380 1680 -360
rect 1700 -380 1720 -360
rect 1740 -380 1760 -360
rect 1780 -380 1800 -360
rect 1820 -380 1840 -360
rect 1860 -380 1880 -360
rect 1900 -380 1920 -360
rect 1940 -380 1960 -360
rect 1980 -380 2000 -360
rect 2020 -380 2040 -360
rect 2060 -380 2080 -360
rect 2100 -380 2120 -360
rect 2140 -380 2160 -360
rect 2180 -380 2200 -360
rect 2220 -380 2240 -360
rect 2260 -380 2280 -360
rect 2300 -380 2320 -360
rect 2340 -380 2360 -360
rect 2380 -380 2400 -360
rect 2420 -380 2440 -360
rect 2460 -380 2480 -360
rect 2500 -380 2520 -360
rect 2540 -380 2560 -360
rect 2580 -380 2600 -360
rect 2620 -380 2640 -360
rect 2660 -380 2680 -360
rect 2700 -380 2720 -360
rect 2740 -380 2760 -360
rect 2780 -380 2800 -360
rect 2820 -380 2840 -360
rect 2860 -380 2880 -360
rect 2900 -380 2920 -360
rect 2940 -380 2960 -360
rect 2980 -380 3000 -360
rect 3020 -380 3040 -360
rect 3060 -380 3080 -360
rect 3100 -380 3120 -360
rect 3140 -380 3160 -360
rect 3180 -380 3200 -360
rect 3220 -380 3240 -360
rect 3260 -380 3280 -360
rect 3300 -380 3320 -360
rect 3340 -380 3360 -360
rect 3380 -380 3400 -360
rect 3420 -380 3440 -360
rect 3460 -380 3480 -360
rect 3500 -380 3520 -360
rect 3540 -380 3560 -360
rect 3580 -380 3600 -360
rect -3470 -480 -3450 -460
rect -3430 -480 -3410 -460
rect -3390 -480 -3370 -460
rect -3350 -480 -3330 -460
rect -3310 -480 -3290 -460
rect -3270 -480 -3250 -460
rect -3230 -480 -3210 -460
rect -3190 -480 -3170 -460
rect -3150 -480 -3130 -460
rect -3110 -480 -3090 -460
rect -3070 -480 -3050 -460
rect -3030 -480 -3010 -460
rect -2990 -480 -2970 -460
rect -2950 -480 -2930 -460
rect -2910 -480 -2890 -460
rect -2870 -480 -2850 -460
rect -2830 -480 -2810 -460
rect -2790 -480 -2770 -460
rect -2750 -480 -2730 -460
rect -2710 -480 -2690 -460
rect -2670 -480 -2650 -460
rect -2630 -480 -2610 -460
rect -2590 -480 -2570 -460
rect -2550 -480 -2530 -460
rect -2510 -480 -2490 -460
rect -2470 -480 -2450 -460
rect -2430 -480 -2410 -460
rect -2390 -480 -2370 -460
rect -2350 -480 -2330 -460
rect -2310 -480 -2290 -460
rect -2270 -480 -2250 -460
rect -2230 -480 -2210 -460
rect -2190 -480 -2170 -460
rect -2150 -480 -2130 -460
rect -2110 -480 -2090 -460
rect -2070 -480 -2050 -460
rect -2030 -480 -2010 -460
rect -1990 -480 -1970 -460
rect -1950 -480 -1930 -460
rect -1910 -480 -1890 -460
rect -1870 -480 -1850 -460
rect -1830 -480 -1810 -460
rect -1790 -480 -1770 -460
rect -1750 -480 -1730 -460
rect -1710 -480 -1690 -460
rect -1670 -480 -1650 -460
rect -1630 -480 -1610 -460
rect -1590 -480 -1570 -460
rect -1550 -480 -1530 -460
rect -1510 -480 -1460 -460
rect -1440 -480 -1420 -460
rect -1400 -480 -1380 -460
rect -1360 -480 -1340 -460
rect -1320 -480 -1300 -460
rect -1280 -480 -1260 -460
rect -1240 -480 -1220 -460
rect -1200 -480 -1180 -460
rect -1160 -480 -1140 -460
rect -1120 -480 -1100 -460
rect -1080 -480 -1060 -460
rect -1040 -480 -1020 -460
rect -1000 -480 -980 -460
rect -960 -480 -940 -460
rect -920 -480 -900 -460
rect -880 -480 -860 -460
rect -840 -480 -820 -460
rect -800 -480 -780 -460
rect -760 -480 -740 -460
rect -720 -480 -700 -460
rect -680 -480 -660 -460
rect -640 -480 -620 -460
rect -600 -480 -580 -460
rect -560 -480 -540 -460
rect -520 -480 -500 -460
rect -480 -480 -460 -460
rect -440 -480 -420 -460
rect -400 -480 -380 -460
rect -360 -480 -340 -460
rect -320 -480 -300 -460
rect -280 -480 -260 -460
rect -230 -480 -210 -460
rect -190 -480 -170 -460
rect -150 -480 -130 -460
rect -110 -480 -90 -460
rect -70 -480 -50 -460
rect -30 -480 -10 -460
rect 10 -480 30 -460
rect 50 -480 80 -460
rect 100 -480 120 -460
rect 140 -480 160 -460
rect 180 -480 200 -460
rect 220 -480 240 -460
rect 260 -480 280 -460
rect 300 -480 320 -460
rect 340 -480 360 -460
rect 390 -480 410 -460
rect 430 -480 450 -460
rect 470 -480 490 -460
rect 510 -480 530 -460
rect 550 -480 570 -460
rect 590 -480 610 -460
rect 630 -480 650 -460
rect 670 -480 690 -460
rect 710 -480 730 -460
rect 750 -480 770 -460
rect 790 -480 810 -460
rect 830 -480 850 -460
rect 870 -480 890 -460
rect 910 -480 930 -460
rect 950 -480 970 -460
rect 990 -480 1010 -460
rect 1030 -480 1050 -460
rect 1070 -480 1090 -460
rect 1110 -480 1130 -460
rect 1150 -480 1170 -460
rect 1190 -480 1210 -460
rect 1230 -480 1250 -460
rect 1270 -480 1290 -460
rect 1310 -480 1330 -460
rect 1350 -480 1370 -460
rect 1390 -480 1410 -460
rect 1430 -480 1450 -460
rect 1470 -480 1490 -460
rect 1510 -480 1530 -460
rect 1550 -480 1570 -460
rect 1590 -480 1640 -460
rect 1660 -480 1680 -460
rect 1700 -480 1720 -460
rect 1740 -480 1760 -460
rect 1780 -480 1800 -460
rect 1820 -480 1840 -460
rect 1860 -480 1880 -460
rect 1900 -480 1920 -460
rect 1940 -480 1960 -460
rect 1980 -480 2000 -460
rect 2020 -480 2040 -460
rect 2060 -480 2080 -460
rect 2100 -480 2120 -460
rect 2140 -480 2160 -460
rect 2180 -480 2200 -460
rect 2220 -480 2240 -460
rect 2260 -480 2280 -460
rect 2300 -480 2320 -460
rect 2340 -480 2360 -460
rect 2380 -480 2400 -460
rect 2420 -480 2440 -460
rect 2460 -480 2480 -460
rect 2500 -480 2520 -460
rect 2540 -480 2560 -460
rect 2580 -480 2600 -460
rect 2620 -480 2640 -460
rect 2660 -480 2680 -460
rect 2700 -480 2720 -460
rect 2740 -480 2760 -460
rect 2780 -480 2800 -460
rect 2820 -480 2840 -460
rect 2860 -480 2880 -460
rect 2900 -480 2920 -460
rect 2940 -480 2960 -460
rect 2980 -480 3000 -460
rect 3020 -480 3040 -460
rect 3060 -480 3080 -460
rect 3100 -480 3120 -460
rect 3140 -480 3160 -460
rect 3180 -480 3200 -460
rect 3220 -480 3240 -460
rect 3260 -480 3280 -460
rect 3300 -480 3320 -460
rect 3340 -480 3360 -460
rect 3380 -480 3400 -460
rect 3420 -480 3440 -460
rect 3460 -480 3480 -460
rect 3500 -480 3520 -460
rect 3540 -480 3560 -460
rect 3580 -480 3600 -460
rect -3470 -580 -3450 -560
rect -3430 -580 -3410 -560
rect -3390 -580 -3370 -560
rect -3350 -580 -3330 -560
rect -3310 -580 -3290 -560
rect -3270 -580 -3250 -560
rect -3230 -580 -3210 -560
rect -3190 -580 -3170 -560
rect -3150 -580 -3130 -560
rect -3110 -580 -3090 -560
rect -3070 -580 -3050 -560
rect -3030 -580 -3010 -560
rect -2990 -580 -2970 -560
rect -2950 -580 -2930 -560
rect -2910 -580 -2890 -560
rect -2870 -580 -2850 -560
rect -2830 -580 -2810 -560
rect -2790 -580 -2770 -560
rect -2750 -580 -2730 -560
rect -2710 -580 -2690 -560
rect -2670 -580 -2650 -560
rect -2630 -580 -2610 -560
rect -2590 -580 -2570 -560
rect -2550 -580 -2530 -560
rect -2510 -580 -2490 -560
rect -2470 -580 -2450 -560
rect -2430 -580 -2410 -560
rect -2390 -580 -2370 -560
rect -2350 -580 -2330 -560
rect -2310 -580 -2290 -560
rect -2270 -580 -2250 -560
rect -2230 -580 -2210 -560
rect -2190 -580 -2170 -560
rect -2150 -580 -2130 -560
rect -2110 -580 -2090 -560
rect -2070 -580 -2050 -560
rect -2030 -580 -2010 -560
rect -1990 -580 -1970 -560
rect -1950 -580 -1930 -560
rect -1910 -580 -1890 -560
rect -1870 -580 -1850 -560
rect -1830 -580 -1810 -560
rect -1790 -580 -1770 -560
rect -1750 -580 -1730 -560
rect -1710 -580 -1690 -560
rect -1670 -580 -1650 -560
rect -1630 -580 -1610 -560
rect -1590 -580 -1570 -560
rect -1550 -580 -1530 -560
rect -1510 -580 -1460 -560
rect -1440 -580 -1420 -560
rect -1400 -580 -1380 -560
rect -1360 -580 -1340 -560
rect -1320 -580 -1300 -560
rect -1280 -580 -1260 -560
rect -1240 -580 -1220 -560
rect -1200 -580 -1180 -560
rect -1160 -580 -1140 -560
rect -1120 -580 -1100 -560
rect -1080 -580 -1060 -560
rect -1040 -580 -1020 -560
rect -1000 -580 -980 -560
rect -960 -580 -940 -560
rect -920 -580 -900 -560
rect -880 -580 -860 -560
rect -840 -580 -820 -560
rect -800 -580 -780 -560
rect -760 -580 -740 -560
rect -720 -580 -700 -560
rect -680 -580 -660 -560
rect -640 -580 -620 -560
rect -600 -580 -580 -560
rect -560 -580 -540 -560
rect -520 -580 -500 -560
rect -480 -580 -460 -560
rect -440 -580 -420 -560
rect -400 -580 -380 -560
rect -360 -580 -340 -560
rect -320 -580 -300 -560
rect -280 -580 -260 -560
rect -230 -580 -210 -560
rect -190 -580 -170 -560
rect -150 -580 -130 -560
rect -110 -580 -90 -560
rect -70 -580 -50 -560
rect -30 -580 -10 -560
rect 10 -580 30 -560
rect 50 -580 80 -560
rect 100 -580 120 -560
rect 140 -580 160 -560
rect 180 -580 200 -560
rect 220 -580 240 -560
rect 260 -580 280 -560
rect 300 -580 320 -560
rect 340 -580 360 -560
rect 390 -580 410 -560
rect 430 -580 450 -560
rect 470 -580 490 -560
rect 510 -580 530 -560
rect 550 -580 570 -560
rect 590 -580 610 -560
rect 630 -580 650 -560
rect 670 -580 690 -560
rect 710 -580 730 -560
rect 750 -580 770 -560
rect 790 -580 810 -560
rect 830 -580 850 -560
rect 870 -580 890 -560
rect 910 -580 930 -560
rect 950 -580 970 -560
rect 990 -580 1010 -560
rect 1030 -580 1050 -560
rect 1070 -580 1090 -560
rect 1110 -580 1130 -560
rect 1150 -580 1170 -560
rect 1190 -580 1210 -560
rect 1230 -580 1250 -560
rect 1270 -580 1290 -560
rect 1310 -580 1330 -560
rect 1350 -580 1370 -560
rect 1390 -580 1410 -560
rect 1430 -580 1450 -560
rect 1470 -580 1490 -560
rect 1510 -580 1530 -560
rect 1550 -580 1570 -560
rect 1590 -580 1640 -560
rect 1660 -580 1680 -560
rect 1700 -580 1720 -560
rect 1740 -580 1760 -560
rect 1780 -580 1800 -560
rect 1820 -580 1840 -560
rect 1860 -580 1880 -560
rect 1900 -580 1920 -560
rect 1940 -580 1960 -560
rect 1980 -580 2000 -560
rect 2020 -580 2040 -560
rect 2060 -580 2080 -560
rect 2100 -580 2120 -560
rect 2140 -580 2160 -560
rect 2180 -580 2200 -560
rect 2220 -580 2240 -560
rect 2260 -580 2280 -560
rect 2300 -580 2320 -560
rect 2340 -580 2360 -560
rect 2380 -580 2400 -560
rect 2420 -580 2440 -560
rect 2460 -580 2480 -560
rect 2500 -580 2520 -560
rect 2540 -580 2560 -560
rect 2580 -580 2600 -560
rect 2620 -580 2640 -560
rect 2660 -580 2680 -560
rect 2700 -580 2720 -560
rect 2740 -580 2760 -560
rect 2780 -580 2800 -560
rect 2820 -580 2840 -560
rect 2860 -580 2880 -560
rect 2900 -580 2920 -560
rect 2940 -580 2960 -560
rect 2980 -580 3000 -560
rect 3020 -580 3040 -560
rect 3060 -580 3080 -560
rect 3100 -580 3120 -560
rect 3140 -580 3160 -560
rect 3180 -580 3200 -560
rect 3220 -580 3240 -560
rect 3260 -580 3280 -560
rect 3300 -580 3320 -560
rect 3340 -580 3360 -560
rect 3380 -580 3400 -560
rect 3420 -580 3440 -560
rect 3460 -580 3480 -560
rect 3500 -580 3520 -560
rect 3540 -580 3560 -560
rect 3580 -580 3600 -560
rect -3470 -680 -3450 -660
rect -3430 -680 -3410 -660
rect -3390 -680 -3370 -660
rect -3350 -680 -3330 -660
rect -3310 -680 -3290 -660
rect -3270 -680 -3250 -660
rect -3230 -680 -3210 -660
rect -3190 -680 -3170 -660
rect -3150 -680 -3130 -660
rect -3110 -680 -3090 -660
rect -3070 -680 -3050 -660
rect -3030 -680 -3010 -660
rect -2990 -680 -2970 -660
rect -2950 -680 -2930 -660
rect -2910 -680 -2890 -660
rect -2870 -680 -2850 -660
rect -2830 -680 -2810 -660
rect -2790 -680 -2770 -660
rect -2750 -680 -2730 -660
rect -2710 -680 -2690 -660
rect -2670 -680 -2650 -660
rect -2630 -680 -2610 -660
rect -2590 -680 -2570 -660
rect -2550 -680 -2530 -660
rect -2510 -680 -2490 -660
rect -2470 -680 -2450 -660
rect -2430 -680 -2410 -660
rect -2390 -680 -2370 -660
rect -2350 -680 -2330 -660
rect -2310 -680 -2290 -660
rect -2270 -680 -2250 -660
rect -2230 -680 -2210 -660
rect -2190 -680 -2170 -660
rect -2150 -680 -2130 -660
rect -2110 -680 -2090 -660
rect -2070 -680 -2050 -660
rect -2030 -680 -2010 -660
rect -1990 -680 -1970 -660
rect -1950 -680 -1930 -660
rect -1910 -680 -1890 -660
rect -1870 -680 -1850 -660
rect -1830 -680 -1810 -660
rect -1790 -680 -1770 -660
rect -1750 -680 -1730 -660
rect -1710 -680 -1690 -660
rect -1670 -680 -1650 -660
rect -1630 -680 -1610 -660
rect -1590 -680 -1570 -660
rect -1550 -680 -1530 -660
rect -1510 -680 -1460 -660
rect -1440 -680 -1420 -660
rect -1400 -680 -1380 -660
rect -1360 -680 -1340 -660
rect -1320 -680 -1300 -660
rect -1280 -680 -1260 -660
rect -1240 -680 -1220 -660
rect -1200 -680 -1180 -660
rect -1160 -680 -1140 -660
rect -1120 -680 -1100 -660
rect -1080 -680 -1060 -660
rect -1040 -680 -1020 -660
rect -1000 -680 -980 -660
rect -960 -680 -940 -660
rect -920 -680 -900 -660
rect -880 -680 -860 -660
rect -840 -680 -820 -660
rect -800 -680 -780 -660
rect -760 -680 -740 -660
rect -720 -680 -700 -660
rect -680 -680 -660 -660
rect -640 -680 -620 -660
rect -600 -680 -580 -660
rect -560 -680 -540 -660
rect -520 -680 -500 -660
rect -480 -680 -460 -660
rect -440 -680 -420 -660
rect -400 -680 -380 -660
rect -360 -680 -340 -660
rect -320 -680 -300 -660
rect -280 -680 -260 -660
rect -230 -680 -210 -660
rect -190 -680 -170 -660
rect -150 -680 -130 -660
rect -110 -680 -90 -660
rect -70 -680 -50 -660
rect -30 -680 -10 -660
rect 10 -680 30 -660
rect 50 -680 80 -660
rect 100 -680 120 -660
rect 140 -680 160 -660
rect 180 -680 200 -660
rect 220 -680 240 -660
rect 260 -680 280 -660
rect 300 -680 320 -660
rect 340 -680 360 -660
rect 390 -680 410 -660
rect 430 -680 450 -660
rect 470 -680 490 -660
rect 510 -680 530 -660
rect 550 -680 570 -660
rect 590 -680 610 -660
rect 630 -680 650 -660
rect 670 -680 690 -660
rect 710 -680 730 -660
rect 750 -680 770 -660
rect 790 -680 810 -660
rect 830 -680 850 -660
rect 870 -680 890 -660
rect 910 -680 930 -660
rect 950 -680 970 -660
rect 990 -680 1010 -660
rect 1030 -680 1050 -660
rect 1070 -680 1090 -660
rect 1110 -680 1130 -660
rect 1150 -680 1170 -660
rect 1190 -680 1210 -660
rect 1230 -680 1250 -660
rect 1270 -680 1290 -660
rect 1310 -680 1330 -660
rect 1350 -680 1370 -660
rect 1390 -680 1410 -660
rect 1430 -680 1450 -660
rect 1470 -680 1490 -660
rect 1510 -680 1530 -660
rect 1550 -680 1570 -660
rect 1590 -680 1640 -660
rect 1660 -680 1680 -660
rect 1700 -680 1720 -660
rect 1740 -680 1760 -660
rect 1780 -680 1800 -660
rect 1820 -680 1840 -660
rect 1860 -680 1880 -660
rect 1900 -680 1920 -660
rect 1940 -680 1960 -660
rect 1980 -680 2000 -660
rect 2020 -680 2040 -660
rect 2060 -680 2080 -660
rect 2100 -680 2120 -660
rect 2140 -680 2160 -660
rect 2180 -680 2200 -660
rect 2220 -680 2240 -660
rect 2260 -680 2280 -660
rect 2300 -680 2320 -660
rect 2340 -680 2360 -660
rect 2380 -680 2400 -660
rect 2420 -680 2440 -660
rect 2460 -680 2480 -660
rect 2500 -680 2520 -660
rect 2540 -680 2560 -660
rect 2580 -680 2600 -660
rect 2620 -680 2640 -660
rect 2660 -680 2680 -660
rect 2700 -680 2720 -660
rect 2740 -680 2760 -660
rect 2780 -680 2800 -660
rect 2820 -680 2840 -660
rect 2860 -680 2880 -660
rect 2900 -680 2920 -660
rect 2940 -680 2960 -660
rect 2980 -680 3000 -660
rect 3020 -680 3040 -660
rect 3060 -680 3080 -660
rect 3100 -680 3120 -660
rect 3140 -680 3160 -660
rect 3180 -680 3200 -660
rect 3220 -680 3240 -660
rect 3260 -680 3280 -660
rect 3300 -680 3320 -660
rect 3340 -680 3360 -660
rect 3380 -680 3400 -660
rect 3420 -680 3440 -660
rect 3460 -680 3480 -660
rect 3500 -680 3520 -660
rect 3540 -680 3560 -660
rect 3580 -680 3600 -660
rect -3470 -780 -3450 -760
rect -3430 -780 -3410 -760
rect -3390 -780 -3370 -760
rect -3350 -780 -3330 -760
rect -3310 -780 -3290 -760
rect -3270 -780 -3250 -760
rect -3230 -780 -3210 -760
rect -3190 -780 -3170 -760
rect -3150 -780 -3130 -760
rect -3110 -780 -3090 -760
rect -3070 -780 -3050 -760
rect -3030 -780 -3010 -760
rect -2990 -780 -2970 -760
rect -2950 -780 -2930 -760
rect -2910 -780 -2890 -760
rect -2870 -780 -2850 -760
rect -2830 -780 -2810 -760
rect -2790 -780 -2770 -760
rect -2750 -780 -2730 -760
rect -2710 -780 -2690 -760
rect -2670 -780 -2650 -760
rect -2630 -780 -2610 -760
rect -2590 -780 -2570 -760
rect -2550 -780 -2530 -760
rect -2510 -780 -2490 -760
rect -2470 -780 -2450 -760
rect -2430 -780 -2410 -760
rect -2390 -780 -2370 -760
rect -2350 -780 -2330 -760
rect -2310 -780 -2290 -760
rect -2270 -780 -2250 -760
rect -2230 -780 -2210 -760
rect -2190 -780 -2170 -760
rect -2150 -780 -2130 -760
rect -2110 -780 -2090 -760
rect -2070 -780 -2050 -760
rect -2030 -780 -2010 -760
rect -1990 -780 -1970 -760
rect -1950 -780 -1930 -760
rect -1910 -780 -1890 -760
rect -1870 -780 -1850 -760
rect -1830 -780 -1810 -760
rect -1790 -780 -1770 -760
rect -1750 -780 -1730 -760
rect -1710 -780 -1690 -760
rect -1670 -780 -1650 -760
rect -1630 -780 -1610 -760
rect -1590 -780 -1570 -760
rect -1550 -780 -1530 -760
rect -1510 -780 -1460 -760
rect -1440 -780 -1420 -760
rect -1400 -780 -1380 -760
rect -1360 -780 -1340 -760
rect -1320 -780 -1300 -760
rect -1280 -780 -1260 -760
rect -1240 -780 -1220 -760
rect -1200 -780 -1180 -760
rect -1160 -780 -1140 -760
rect -1120 -780 -1100 -760
rect -1080 -780 -1060 -760
rect -1040 -780 -1020 -760
rect -1000 -780 -980 -760
rect -960 -780 -940 -760
rect -920 -780 -900 -760
rect -880 -780 -860 -760
rect -840 -780 -820 -760
rect -800 -780 -780 -760
rect -760 -780 -740 -760
rect -720 -780 -700 -760
rect -680 -780 -660 -760
rect -640 -780 -620 -760
rect -600 -780 -580 -760
rect -560 -780 -540 -760
rect -520 -780 -500 -760
rect -480 -780 -460 -760
rect -440 -780 -420 -760
rect -400 -780 -380 -760
rect -360 -780 -340 -760
rect -320 -780 -300 -760
rect -280 -780 -260 -760
rect -230 -780 -210 -760
rect -190 -780 -170 -760
rect -150 -780 -130 -760
rect -110 -780 -90 -760
rect -70 -780 -50 -760
rect -30 -780 -10 -760
rect 10 -780 30 -760
rect 50 -780 80 -760
rect 100 -780 120 -760
rect 140 -780 160 -760
rect 180 -780 200 -760
rect 220 -780 240 -760
rect 260 -780 280 -760
rect 300 -780 320 -760
rect 340 -780 360 -760
rect 390 -780 410 -760
rect 430 -780 450 -760
rect 470 -780 490 -760
rect 510 -780 530 -760
rect 550 -780 570 -760
rect 590 -780 610 -760
rect 630 -780 650 -760
rect 670 -780 690 -760
rect 710 -780 730 -760
rect 750 -780 770 -760
rect 790 -780 810 -760
rect 830 -780 850 -760
rect 870 -780 890 -760
rect 910 -780 930 -760
rect 950 -780 970 -760
rect 990 -780 1010 -760
rect 1030 -780 1050 -760
rect 1070 -780 1090 -760
rect 1110 -780 1130 -760
rect 1150 -780 1170 -760
rect 1190 -780 1210 -760
rect 1230 -780 1250 -760
rect 1270 -780 1290 -760
rect 1310 -780 1330 -760
rect 1350 -780 1370 -760
rect 1390 -780 1410 -760
rect 1430 -780 1450 -760
rect 1470 -780 1490 -760
rect 1510 -780 1530 -760
rect 1550 -780 1570 -760
rect 1590 -780 1640 -760
rect 1660 -780 1680 -760
rect 1700 -780 1720 -760
rect 1740 -780 1760 -760
rect 1780 -780 1800 -760
rect 1820 -780 1840 -760
rect 1860 -780 1880 -760
rect 1900 -780 1920 -760
rect 1940 -780 1960 -760
rect 1980 -780 2000 -760
rect 2020 -780 2040 -760
rect 2060 -780 2080 -760
rect 2100 -780 2120 -760
rect 2140 -780 2160 -760
rect 2180 -780 2200 -760
rect 2220 -780 2240 -760
rect 2260 -780 2280 -760
rect 2300 -780 2320 -760
rect 2340 -780 2360 -760
rect 2380 -780 2400 -760
rect 2420 -780 2440 -760
rect 2460 -780 2480 -760
rect 2500 -780 2520 -760
rect 2540 -780 2560 -760
rect 2580 -780 2600 -760
rect 2620 -780 2640 -760
rect 2660 -780 2680 -760
rect 2700 -780 2720 -760
rect 2740 -780 2760 -760
rect 2780 -780 2800 -760
rect 2820 -780 2840 -760
rect 2860 -780 2880 -760
rect 2900 -780 2920 -760
rect 2940 -780 2960 -760
rect 2980 -780 3000 -760
rect 3020 -780 3040 -760
rect 3060 -780 3080 -760
rect 3100 -780 3120 -760
rect 3140 -780 3160 -760
rect 3180 -780 3200 -760
rect 3220 -780 3240 -760
rect 3260 -780 3280 -760
rect 3300 -780 3320 -760
rect 3340 -780 3360 -760
rect 3380 -780 3400 -760
rect 3420 -780 3440 -760
rect 3460 -780 3480 -760
rect 3500 -780 3520 -760
rect 3540 -780 3560 -760
rect 3580 -780 3600 -760
rect -3470 -880 -3450 -860
rect -3430 -880 -3410 -860
rect -3390 -880 -3370 -860
rect -3350 -880 -3330 -860
rect -3310 -880 -3290 -860
rect -3270 -880 -3250 -860
rect -3230 -880 -3210 -860
rect -3190 -880 -3170 -860
rect -3150 -880 -3130 -860
rect -3110 -880 -3090 -860
rect -3070 -880 -3050 -860
rect -3030 -880 -3010 -860
rect -2990 -880 -2970 -860
rect -2950 -880 -2930 -860
rect -2910 -880 -2890 -860
rect -2870 -880 -2850 -860
rect -2830 -880 -2810 -860
rect -2790 -880 -2770 -860
rect -2750 -880 -2730 -860
rect -2710 -880 -2690 -860
rect -2670 -880 -2650 -860
rect -2630 -880 -2610 -860
rect -2590 -880 -2570 -860
rect -2550 -880 -2530 -860
rect -2510 -880 -2490 -860
rect -2470 -880 -2450 -860
rect -2430 -880 -2410 -860
rect -2390 -880 -2370 -860
rect -2350 -880 -2330 -860
rect -2310 -880 -2290 -860
rect -2270 -880 -2250 -860
rect -2230 -880 -2210 -860
rect -2190 -880 -2170 -860
rect -2150 -880 -2130 -860
rect -2110 -880 -2090 -860
rect -2070 -880 -2050 -860
rect -2030 -880 -2010 -860
rect -1990 -880 -1970 -860
rect -1950 -880 -1930 -860
rect -1910 -880 -1890 -860
rect -1870 -880 -1850 -860
rect -1830 -880 -1810 -860
rect -1790 -880 -1770 -860
rect -1750 -880 -1730 -860
rect -1710 -880 -1690 -860
rect -1670 -880 -1650 -860
rect -1630 -880 -1610 -860
rect -1590 -880 -1570 -860
rect -1550 -880 -1530 -860
rect -1510 -880 -1460 -860
rect -1440 -880 -1420 -860
rect -1400 -880 -1380 -860
rect -1360 -880 -1340 -860
rect -1320 -880 -1300 -860
rect -1280 -880 -1260 -860
rect -1240 -880 -1220 -860
rect -1200 -880 -1180 -860
rect -1160 -880 -1140 -860
rect -1120 -880 -1100 -860
rect -1080 -880 -1060 -860
rect -1040 -880 -1020 -860
rect -1000 -880 -980 -860
rect -960 -880 -940 -860
rect -920 -880 -900 -860
rect -880 -880 -860 -860
rect -840 -880 -820 -860
rect -800 -880 -780 -860
rect -760 -880 -740 -860
rect -720 -880 -700 -860
rect -680 -880 -660 -860
rect -640 -880 -620 -860
rect -600 -880 -580 -860
rect -560 -880 -540 -860
rect -520 -880 -500 -860
rect -480 -880 -460 -860
rect -440 -880 -420 -860
rect -400 -880 -380 -860
rect -360 -880 -340 -860
rect -320 -880 -300 -860
rect -280 -880 -260 -860
rect -230 -880 -210 -860
rect -190 -880 -170 -860
rect -150 -880 -130 -860
rect -110 -880 -90 -860
rect -70 -880 -50 -860
rect -30 -880 -10 -860
rect 10 -880 30 -860
rect 50 -880 80 -860
rect 100 -880 120 -860
rect 140 -880 160 -860
rect 180 -880 200 -860
rect 220 -880 240 -860
rect 260 -880 280 -860
rect 300 -880 320 -860
rect 340 -880 360 -860
rect 390 -880 410 -860
rect 430 -880 450 -860
rect 470 -880 490 -860
rect 510 -880 530 -860
rect 550 -880 570 -860
rect 590 -880 610 -860
rect 630 -880 650 -860
rect 670 -880 690 -860
rect 710 -880 730 -860
rect 750 -880 770 -860
rect 790 -880 810 -860
rect 830 -880 850 -860
rect 870 -880 890 -860
rect 910 -880 930 -860
rect 950 -880 970 -860
rect 990 -880 1010 -860
rect 1030 -880 1050 -860
rect 1070 -880 1090 -860
rect 1110 -880 1130 -860
rect 1150 -880 1170 -860
rect 1190 -880 1210 -860
rect 1230 -880 1250 -860
rect 1270 -880 1290 -860
rect 1310 -880 1330 -860
rect 1350 -880 1370 -860
rect 1390 -880 1410 -860
rect 1430 -880 1450 -860
rect 1470 -880 1490 -860
rect 1510 -880 1530 -860
rect 1550 -880 1570 -860
rect 1590 -880 1640 -860
rect 1660 -880 1680 -860
rect 1700 -880 1720 -860
rect 1740 -880 1760 -860
rect 1780 -880 1800 -860
rect 1820 -880 1840 -860
rect 1860 -880 1880 -860
rect 1900 -880 1920 -860
rect 1940 -880 1960 -860
rect 1980 -880 2000 -860
rect 2020 -880 2040 -860
rect 2060 -880 2080 -860
rect 2100 -880 2120 -860
rect 2140 -880 2160 -860
rect 2180 -880 2200 -860
rect 2220 -880 2240 -860
rect 2260 -880 2280 -860
rect 2300 -880 2320 -860
rect 2340 -880 2360 -860
rect 2380 -880 2400 -860
rect 2420 -880 2440 -860
rect 2460 -880 2480 -860
rect 2500 -880 2520 -860
rect 2540 -880 2560 -860
rect 2580 -880 2600 -860
rect 2620 -880 2640 -860
rect 2660 -880 2680 -860
rect 2700 -880 2720 -860
rect 2740 -880 2760 -860
rect 2780 -880 2800 -860
rect 2820 -880 2840 -860
rect 2860 -880 2880 -860
rect 2900 -880 2920 -860
rect 2940 -880 2960 -860
rect 2980 -880 3000 -860
rect 3020 -880 3040 -860
rect 3060 -880 3080 -860
rect 3100 -880 3120 -860
rect 3140 -880 3160 -860
rect 3180 -880 3200 -860
rect 3220 -880 3240 -860
rect 3260 -880 3280 -860
rect 3300 -880 3320 -860
rect 3340 -880 3360 -860
rect 3380 -880 3400 -860
rect 3420 -880 3440 -860
rect 3460 -880 3480 -860
rect 3500 -880 3520 -860
rect 3540 -880 3560 -860
rect 3580 -880 3600 -860
rect -3470 -980 -3450 -960
rect -3430 -980 -3410 -960
rect -3390 -980 -3370 -960
rect -3350 -980 -3330 -960
rect -3310 -980 -3290 -960
rect -3270 -980 -3250 -960
rect -3230 -980 -3210 -960
rect -3190 -980 -3170 -960
rect -3150 -980 -3130 -960
rect -3110 -980 -3090 -960
rect -3070 -980 -3050 -960
rect -3030 -980 -3010 -960
rect -2990 -980 -2970 -960
rect -2950 -980 -2930 -960
rect -2910 -980 -2890 -960
rect -2870 -980 -2850 -960
rect -2830 -980 -2810 -960
rect -2790 -980 -2770 -960
rect -2750 -980 -2730 -960
rect -2710 -980 -2690 -960
rect -2670 -980 -2650 -960
rect -2630 -980 -2610 -960
rect -2590 -980 -2570 -960
rect -2550 -980 -2530 -960
rect -2510 -980 -2490 -960
rect -2470 -980 -2450 -960
rect -2430 -980 -2410 -960
rect -2390 -980 -2370 -960
rect -2350 -980 -2330 -960
rect -2310 -980 -2290 -960
rect -2270 -980 -2250 -960
rect -2230 -980 -2210 -960
rect -2190 -980 -2170 -960
rect -2150 -980 -2130 -960
rect -2110 -980 -2090 -960
rect -2070 -980 -2050 -960
rect -2030 -980 -2010 -960
rect -1990 -980 -1970 -960
rect -1950 -980 -1930 -960
rect -1910 -980 -1890 -960
rect -1870 -980 -1850 -960
rect -1830 -980 -1810 -960
rect -1790 -980 -1770 -960
rect -1750 -980 -1730 -960
rect -1710 -980 -1690 -960
rect -1670 -980 -1650 -960
rect -1630 -980 -1610 -960
rect -1590 -980 -1570 -960
rect -1550 -980 -1530 -960
rect -1510 -980 -1460 -960
rect -1440 -980 -1420 -960
rect -1400 -980 -1380 -960
rect -1360 -980 -1340 -960
rect -1320 -980 -1300 -960
rect -1280 -980 -1260 -960
rect -1240 -980 -1220 -960
rect -1200 -980 -1180 -960
rect -1160 -980 -1140 -960
rect -1120 -980 -1100 -960
rect -1080 -980 -1060 -960
rect -1040 -980 -1020 -960
rect -1000 -980 -980 -960
rect -960 -980 -940 -960
rect -920 -980 -900 -960
rect -880 -980 -860 -960
rect -840 -980 -820 -960
rect -800 -980 -780 -960
rect -760 -980 -740 -960
rect -720 -980 -700 -960
rect -680 -980 -660 -960
rect -640 -980 -620 -960
rect -600 -980 -580 -960
rect -560 -980 -540 -960
rect -520 -980 -500 -960
rect -480 -980 -460 -960
rect -440 -980 -420 -960
rect -400 -980 -380 -960
rect -360 -980 -340 -960
rect -320 -980 -300 -960
rect -280 -980 -260 -960
rect -230 -980 -210 -960
rect -190 -980 -170 -960
rect -150 -980 -130 -960
rect -110 -980 -90 -960
rect -70 -980 -50 -960
rect -30 -980 -10 -960
rect 10 -980 30 -960
rect 50 -980 80 -960
rect 100 -980 120 -960
rect 140 -980 160 -960
rect 180 -980 200 -960
rect 220 -980 240 -960
rect 260 -980 280 -960
rect 300 -980 320 -960
rect 340 -980 360 -960
rect 390 -980 410 -960
rect 430 -980 450 -960
rect 470 -980 490 -960
rect 510 -980 530 -960
rect 550 -980 570 -960
rect 590 -980 610 -960
rect 630 -980 650 -960
rect 670 -980 690 -960
rect 710 -980 730 -960
rect 750 -980 770 -960
rect 790 -980 810 -960
rect 830 -980 850 -960
rect 870 -980 890 -960
rect 910 -980 930 -960
rect 950 -980 970 -960
rect 990 -980 1010 -960
rect 1030 -980 1050 -960
rect 1070 -980 1090 -960
rect 1110 -980 1130 -960
rect 1150 -980 1170 -960
rect 1190 -980 1210 -960
rect 1230 -980 1250 -960
rect 1270 -980 1290 -960
rect 1310 -980 1330 -960
rect 1350 -980 1370 -960
rect 1390 -980 1410 -960
rect 1430 -980 1450 -960
rect 1470 -980 1490 -960
rect 1510 -980 1530 -960
rect 1550 -980 1570 -960
rect 1590 -980 1640 -960
rect 1660 -980 1680 -960
rect 1700 -980 1720 -960
rect 1740 -980 1760 -960
rect 1780 -980 1800 -960
rect 1820 -980 1840 -960
rect 1860 -980 1880 -960
rect 1900 -980 1920 -960
rect 1940 -980 1960 -960
rect 1980 -980 2000 -960
rect 2020 -980 2040 -960
rect 2060 -980 2080 -960
rect 2100 -980 2120 -960
rect 2140 -980 2160 -960
rect 2180 -980 2200 -960
rect 2220 -980 2240 -960
rect 2260 -980 2280 -960
rect 2300 -980 2320 -960
rect 2340 -980 2360 -960
rect 2380 -980 2400 -960
rect 2420 -980 2440 -960
rect 2460 -980 2480 -960
rect 2500 -980 2520 -960
rect 2540 -980 2560 -960
rect 2580 -980 2600 -960
rect 2620 -980 2640 -960
rect 2660 -980 2680 -960
rect 2700 -980 2720 -960
rect 2740 -980 2760 -960
rect 2780 -980 2800 -960
rect 2820 -980 2840 -960
rect 2860 -980 2880 -960
rect 2900 -980 2920 -960
rect 2940 -980 2960 -960
rect 2980 -980 3000 -960
rect 3020 -980 3040 -960
rect 3060 -980 3080 -960
rect 3100 -980 3120 -960
rect 3140 -980 3160 -960
rect 3180 -980 3200 -960
rect 3220 -980 3240 -960
rect 3260 -980 3280 -960
rect 3300 -980 3320 -960
rect 3340 -980 3360 -960
rect 3380 -980 3400 -960
rect 3420 -980 3440 -960
rect 3460 -980 3480 -960
rect 3500 -980 3520 -960
rect 3540 -980 3560 -960
rect 3580 -980 3600 -960
rect -3470 -1080 -3450 -1060
rect -3430 -1080 -3410 -1060
rect -3390 -1080 -3370 -1060
rect -3350 -1080 -3330 -1060
rect -3310 -1080 -3290 -1060
rect -3270 -1080 -3250 -1060
rect -3230 -1080 -3210 -1060
rect -3190 -1080 -3170 -1060
rect -3150 -1080 -3130 -1060
rect -3110 -1080 -3090 -1060
rect -3070 -1080 -3050 -1060
rect -3030 -1080 -3010 -1060
rect -2990 -1080 -2970 -1060
rect -2950 -1080 -2930 -1060
rect -2910 -1080 -2890 -1060
rect -2870 -1080 -2850 -1060
rect -2830 -1080 -2810 -1060
rect -2790 -1080 -2770 -1060
rect -2750 -1080 -2730 -1060
rect -2710 -1080 -2690 -1060
rect -2670 -1080 -2650 -1060
rect -2630 -1080 -2610 -1060
rect -2590 -1080 -2570 -1060
rect -2550 -1080 -2530 -1060
rect -2510 -1080 -2490 -1060
rect -2470 -1080 -2450 -1060
rect -2430 -1080 -2410 -1060
rect -2390 -1080 -2370 -1060
rect -2350 -1080 -2330 -1060
rect -2310 -1080 -2290 -1060
rect -2270 -1080 -2250 -1060
rect -2230 -1080 -2210 -1060
rect -2190 -1080 -2170 -1060
rect -2150 -1080 -2130 -1060
rect -2110 -1080 -2090 -1060
rect -2070 -1080 -2050 -1060
rect -2030 -1080 -2010 -1060
rect -1990 -1080 -1970 -1060
rect -1950 -1080 -1930 -1060
rect -1910 -1080 -1890 -1060
rect -1870 -1080 -1850 -1060
rect -1830 -1080 -1810 -1060
rect -1790 -1080 -1770 -1060
rect -1750 -1080 -1730 -1060
rect -1710 -1080 -1690 -1060
rect -1670 -1080 -1650 -1060
rect -1630 -1080 -1610 -1060
rect -1590 -1080 -1570 -1060
rect -1550 -1080 -1530 -1060
rect -1510 -1080 -1460 -1060
rect -1440 -1080 -1420 -1060
rect -1400 -1080 -1380 -1060
rect -1360 -1080 -1340 -1060
rect -1320 -1080 -1300 -1060
rect -1280 -1080 -1260 -1060
rect -1240 -1080 -1220 -1060
rect -1200 -1080 -1180 -1060
rect -1160 -1080 -1140 -1060
rect -1120 -1080 -1100 -1060
rect -1080 -1080 -1060 -1060
rect -1040 -1080 -1020 -1060
rect -1000 -1080 -980 -1060
rect -960 -1080 -940 -1060
rect -920 -1080 -900 -1060
rect -880 -1080 -860 -1060
rect -840 -1080 -820 -1060
rect -800 -1080 -780 -1060
rect -760 -1080 -740 -1060
rect -720 -1080 -700 -1060
rect -680 -1080 -660 -1060
rect -640 -1080 -620 -1060
rect -600 -1080 -580 -1060
rect -560 -1080 -540 -1060
rect -520 -1080 -500 -1060
rect -480 -1080 -460 -1060
rect -440 -1080 -420 -1060
rect -400 -1080 -380 -1060
rect -360 -1080 -340 -1060
rect -320 -1080 -300 -1060
rect -280 -1080 -260 -1060
rect -230 -1080 -210 -1060
rect -190 -1080 -170 -1060
rect -150 -1080 -130 -1060
rect -110 -1080 -90 -1060
rect -70 -1080 -50 -1060
rect -30 -1080 -10 -1060
rect 10 -1080 30 -1060
rect 50 -1080 80 -1060
rect 100 -1080 120 -1060
rect 140 -1080 160 -1060
rect 180 -1080 200 -1060
rect 220 -1080 240 -1060
rect 260 -1080 280 -1060
rect 300 -1080 320 -1060
rect 340 -1080 360 -1060
rect 390 -1080 410 -1060
rect 430 -1080 450 -1060
rect 470 -1080 490 -1060
rect 510 -1080 530 -1060
rect 550 -1080 570 -1060
rect 590 -1080 610 -1060
rect 630 -1080 650 -1060
rect 670 -1080 690 -1060
rect 710 -1080 730 -1060
rect 750 -1080 770 -1060
rect 790 -1080 810 -1060
rect 830 -1080 850 -1060
rect 870 -1080 890 -1060
rect 910 -1080 930 -1060
rect 950 -1080 970 -1060
rect 990 -1080 1010 -1060
rect 1030 -1080 1050 -1060
rect 1070 -1080 1090 -1060
rect 1110 -1080 1130 -1060
rect 1150 -1080 1170 -1060
rect 1190 -1080 1210 -1060
rect 1230 -1080 1250 -1060
rect 1270 -1080 1290 -1060
rect 1310 -1080 1330 -1060
rect 1350 -1080 1370 -1060
rect 1390 -1080 1410 -1060
rect 1430 -1080 1450 -1060
rect 1470 -1080 1490 -1060
rect 1510 -1080 1530 -1060
rect 1550 -1080 1570 -1060
rect 1590 -1080 1640 -1060
rect 1660 -1080 1680 -1060
rect 1700 -1080 1720 -1060
rect 1740 -1080 1760 -1060
rect 1780 -1080 1800 -1060
rect 1820 -1080 1840 -1060
rect 1860 -1080 1880 -1060
rect 1900 -1080 1920 -1060
rect 1940 -1080 1960 -1060
rect 1980 -1080 2000 -1060
rect 2020 -1080 2040 -1060
rect 2060 -1080 2080 -1060
rect 2100 -1080 2120 -1060
rect 2140 -1080 2160 -1060
rect 2180 -1080 2200 -1060
rect 2220 -1080 2240 -1060
rect 2260 -1080 2280 -1060
rect 2300 -1080 2320 -1060
rect 2340 -1080 2360 -1060
rect 2380 -1080 2400 -1060
rect 2420 -1080 2440 -1060
rect 2460 -1080 2480 -1060
rect 2500 -1080 2520 -1060
rect 2540 -1080 2560 -1060
rect 2580 -1080 2600 -1060
rect 2620 -1080 2640 -1060
rect 2660 -1080 2680 -1060
rect 2700 -1080 2720 -1060
rect 2740 -1080 2760 -1060
rect 2780 -1080 2800 -1060
rect 2820 -1080 2840 -1060
rect 2860 -1080 2880 -1060
rect 2900 -1080 2920 -1060
rect 2940 -1080 2960 -1060
rect 2980 -1080 3000 -1060
rect 3020 -1080 3040 -1060
rect 3060 -1080 3080 -1060
rect 3100 -1080 3120 -1060
rect 3140 -1080 3160 -1060
rect 3180 -1080 3200 -1060
rect 3220 -1080 3240 -1060
rect 3260 -1080 3280 -1060
rect 3300 -1080 3320 -1060
rect 3340 -1080 3360 -1060
rect 3380 -1080 3400 -1060
rect 3420 -1080 3440 -1060
rect 3460 -1080 3480 -1060
rect 3500 -1080 3520 -1060
rect 3540 -1080 3560 -1060
rect 3580 -1080 3600 -1060
rect -3470 -1180 -3450 -1160
rect -3430 -1180 -3410 -1160
rect -3390 -1180 -3370 -1160
rect -3350 -1180 -3330 -1160
rect -3310 -1180 -3290 -1160
rect -3270 -1180 -3250 -1160
rect -3230 -1180 -3210 -1160
rect -3190 -1180 -3170 -1160
rect -3150 -1180 -3130 -1160
rect -3110 -1180 -3090 -1160
rect -3070 -1180 -3050 -1160
rect -3030 -1180 -3010 -1160
rect -2990 -1180 -2970 -1160
rect -2950 -1180 -2930 -1160
rect -2910 -1180 -2890 -1160
rect -2870 -1180 -2850 -1160
rect -2830 -1180 -2810 -1160
rect -2790 -1180 -2770 -1160
rect -2750 -1180 -2730 -1160
rect -2710 -1180 -2690 -1160
rect -2670 -1180 -2650 -1160
rect -2630 -1180 -2610 -1160
rect -2590 -1180 -2570 -1160
rect -2550 -1180 -2530 -1160
rect -2510 -1180 -2490 -1160
rect -2470 -1180 -2450 -1160
rect -2430 -1180 -2410 -1160
rect -2390 -1180 -2370 -1160
rect -2350 -1180 -2330 -1160
rect -2310 -1180 -2290 -1160
rect -2270 -1180 -2250 -1160
rect -2230 -1180 -2210 -1160
rect -2190 -1180 -2170 -1160
rect -2150 -1180 -2130 -1160
rect -2110 -1180 -2090 -1160
rect -2070 -1180 -2050 -1160
rect -2030 -1180 -2010 -1160
rect -1990 -1180 -1970 -1160
rect -1950 -1180 -1930 -1160
rect -1910 -1180 -1890 -1160
rect -1870 -1180 -1850 -1160
rect -1830 -1180 -1810 -1160
rect -1790 -1180 -1770 -1160
rect -1750 -1180 -1730 -1160
rect -1710 -1180 -1690 -1160
rect -1670 -1180 -1650 -1160
rect -1630 -1180 -1610 -1160
rect -1590 -1180 -1570 -1160
rect -1550 -1180 -1530 -1160
rect -1510 -1180 -1490 -1160
rect -1470 -1180 -1450 -1160
rect -1430 -1180 -1410 -1160
rect -1390 -1180 -1370 -1160
rect -1350 -1180 -1330 -1160
rect -1310 -1180 -1290 -1160
rect -1270 -1180 -1250 -1160
rect -1230 -1180 -1210 -1160
rect -1190 -1180 -1170 -1160
rect -1150 -1180 -1130 -1160
rect -1110 -1180 -1090 -1160
rect -1070 -1180 -1050 -1160
rect -1030 -1180 -1010 -1160
rect -990 -1180 -970 -1160
rect -950 -1180 -930 -1160
rect -910 -1180 -890 -1160
rect -870 -1180 -850 -1160
rect -830 -1180 -810 -1160
rect -790 -1180 -770 -1160
rect -750 -1180 -730 -1160
rect -710 -1180 -690 -1160
rect -670 -1180 -650 -1160
rect -630 -1180 -610 -1160
rect -590 -1180 -570 -1160
rect -550 -1180 -530 -1160
rect -510 -1180 -490 -1160
rect -470 -1180 -450 -1160
rect -430 -1180 -410 -1160
rect -390 -1180 -370 -1160
rect -350 -1180 -330 -1160
rect -310 -1180 -290 -1160
rect -270 -1180 -250 -1160
rect -230 -1180 -210 -1160
rect -190 -1180 -170 -1160
rect -150 -1180 -130 -1160
rect -110 -1180 -90 -1160
rect -70 -1180 -50 -1160
rect -30 -1180 -10 -1160
rect 10 -1180 30 -1160
rect 50 -1180 80 -1160
rect 100 -1180 120 -1160
rect 140 -1180 160 -1160
rect 180 -1180 200 -1160
rect 220 -1180 240 -1160
rect 260 -1180 280 -1160
rect 300 -1180 320 -1160
rect 340 -1180 360 -1160
rect 380 -1180 400 -1160
rect 420 -1180 440 -1160
rect 460 -1180 480 -1160
rect 500 -1180 520 -1160
rect 540 -1180 560 -1160
rect 580 -1180 600 -1160
rect 620 -1180 640 -1160
rect 660 -1180 680 -1160
rect 700 -1180 720 -1160
rect 740 -1180 760 -1160
rect 780 -1180 800 -1160
rect 820 -1180 840 -1160
rect 860 -1180 880 -1160
rect 900 -1180 920 -1160
rect 940 -1180 960 -1160
rect 980 -1180 1000 -1160
rect 1020 -1180 1040 -1160
rect 1060 -1180 1080 -1160
rect 1100 -1180 1120 -1160
rect 1140 -1180 1160 -1160
rect 1180 -1180 1200 -1160
rect 1220 -1180 1240 -1160
rect 1260 -1180 1280 -1160
rect 1300 -1180 1320 -1160
rect 1340 -1180 1360 -1160
rect 1380 -1180 1400 -1160
rect 1420 -1180 1440 -1160
rect 1460 -1180 1480 -1160
rect 1500 -1180 1520 -1160
rect 1540 -1180 1560 -1160
rect 1580 -1180 1600 -1160
rect 1620 -1180 1640 -1160
rect 1660 -1180 1680 -1160
rect 1700 -1180 1720 -1160
rect 1740 -1180 1760 -1160
rect 1780 -1180 1800 -1160
rect 1820 -1180 1840 -1160
rect 1860 -1180 1880 -1160
rect 1900 -1180 1920 -1160
rect 1940 -1180 1960 -1160
rect 1980 -1180 2000 -1160
rect 2020 -1180 2040 -1160
rect 2060 -1180 2080 -1160
rect 2100 -1180 2120 -1160
rect 2140 -1180 2160 -1160
rect 2180 -1180 2200 -1160
rect 2220 -1180 2240 -1160
rect 2260 -1180 2280 -1160
rect 2300 -1180 2320 -1160
rect 2340 -1180 2360 -1160
rect 2380 -1180 2400 -1160
rect 2420 -1180 2440 -1160
rect 2460 -1180 2480 -1160
rect 2500 -1180 2520 -1160
rect 2540 -1180 2560 -1160
rect 2580 -1180 2600 -1160
rect 2620 -1180 2640 -1160
rect 2660 -1180 2680 -1160
rect 2700 -1180 2720 -1160
rect 2740 -1180 2760 -1160
rect 2780 -1180 2800 -1160
rect 2820 -1180 2840 -1160
rect 2860 -1180 2880 -1160
rect 2900 -1180 2920 -1160
rect 2940 -1180 2960 -1160
rect 2980 -1180 3000 -1160
rect 3020 -1180 3040 -1160
rect 3060 -1180 3080 -1160
rect 3100 -1180 3120 -1160
rect 3140 -1180 3160 -1160
rect 3180 -1180 3200 -1160
rect 3220 -1180 3240 -1160
rect 3260 -1180 3280 -1160
rect 3300 -1180 3320 -1160
rect 3340 -1180 3360 -1160
rect 3380 -1180 3400 -1160
rect 3420 -1180 3440 -1160
rect 3460 -1180 3480 -1160
rect 3500 -1180 3520 -1160
rect 3540 -1180 3560 -1160
rect 3580 -1180 3600 -1160
<< psubdiff >>
rect -3485 -120 3615 -110
rect -3485 -140 -3470 -120
rect -3450 -140 -3430 -120
rect -3410 -140 -3390 -120
rect -3370 -140 -3350 -120
rect -3330 -140 -3310 -120
rect -3290 -140 -3270 -120
rect -3250 -140 -3230 -120
rect -3210 -140 -3190 -120
rect -3170 -140 -3150 -120
rect -3130 -140 -3110 -120
rect -3090 -140 -3070 -120
rect -3050 -140 -3030 -120
rect -3010 -140 -2990 -120
rect -2970 -140 -2950 -120
rect -2930 -140 -2910 -120
rect -2890 -140 -2870 -120
rect -2850 -140 -2830 -120
rect -2810 -140 -2790 -120
rect -2770 -140 -2750 -120
rect -2730 -140 -2710 -120
rect -2690 -140 -2670 -120
rect -2650 -140 -2630 -120
rect -2610 -140 -2590 -120
rect -2570 -140 -2550 -120
rect -2530 -140 -2510 -120
rect -2490 -140 -2470 -120
rect -2450 -140 -2430 -120
rect -2410 -140 -2390 -120
rect -2370 -140 -2350 -120
rect -2330 -140 -2310 -120
rect -2290 -140 -2270 -120
rect -2250 -140 -2230 -120
rect -2210 -140 -2190 -120
rect -2170 -140 -2150 -120
rect -2130 -140 -2110 -120
rect -2090 -140 -2070 -120
rect -2050 -140 -2030 -120
rect -2010 -140 -1990 -120
rect -1970 -140 -1950 -120
rect -1930 -140 -1910 -120
rect -1890 -140 -1870 -120
rect -1850 -140 -1830 -120
rect -1810 -140 -1790 -120
rect -1770 -140 -1750 -120
rect -1730 -140 -1710 -120
rect -1690 -140 -1670 -120
rect -1650 -140 -1630 -120
rect -1610 -140 -1590 -120
rect -1570 -140 -1550 -120
rect -1530 -140 -1510 -120
rect -1460 -140 -1440 -120
rect -1420 -140 -1400 -120
rect -1380 -140 -1360 -120
rect -1340 -140 -1320 -120
rect -1300 -140 -1280 -120
rect -1260 -140 -1240 -120
rect -1220 -140 -1200 -120
rect -1180 -140 -1160 -120
rect -1140 -140 -1120 -120
rect -1100 -140 -1080 -120
rect -1060 -140 -1040 -120
rect -1020 -140 -1000 -120
rect -980 -140 -960 -120
rect -940 -140 -920 -120
rect -900 -140 -880 -120
rect -860 -140 -840 -120
rect -820 -140 -800 -120
rect -780 -140 -760 -120
rect -740 -140 -720 -120
rect -700 -140 -680 -120
rect -660 -140 -640 -120
rect -620 -140 -600 -120
rect -580 -140 -560 -120
rect -540 -140 -520 -120
rect -500 -140 -480 -120
rect -460 -140 -440 -120
rect -420 -140 -400 -120
rect -380 -140 -360 -120
rect -340 -140 -320 -120
rect -300 -140 -280 -120
rect -260 -140 -230 -120
rect -210 -140 -190 -120
rect -170 -140 -150 -120
rect -130 -140 -110 -120
rect -90 -140 -70 -120
rect -50 -140 -30 -120
rect -10 -140 10 -120
rect 30 -140 50 -120
rect 80 -140 100 -120
rect 120 -140 140 -120
rect 160 -140 180 -120
rect 200 -140 220 -120
rect 240 -140 260 -120
rect 280 -140 300 -120
rect 320 -140 340 -120
rect 360 -140 390 -120
rect 410 -140 430 -120
rect 450 -140 470 -120
rect 490 -140 510 -120
rect 530 -140 550 -120
rect 570 -140 590 -120
rect 610 -140 630 -120
rect 650 -140 670 -120
rect 690 -140 710 -120
rect 730 -140 750 -120
rect 770 -140 790 -120
rect 810 -140 830 -120
rect 850 -140 870 -120
rect 890 -140 910 -120
rect 930 -140 950 -120
rect 970 -140 990 -120
rect 1010 -140 1030 -120
rect 1050 -140 1070 -120
rect 1090 -140 1110 -120
rect 1130 -140 1150 -120
rect 1170 -140 1190 -120
rect 1210 -140 1230 -120
rect 1250 -140 1270 -120
rect 1290 -140 1310 -120
rect 1330 -140 1350 -120
rect 1370 -140 1390 -120
rect 1410 -140 1430 -120
rect 1450 -140 1470 -120
rect 1490 -140 1510 -120
rect 1530 -140 1550 -120
rect 1570 -140 1590 -120
rect 1640 -140 1660 -120
rect 1680 -140 1700 -120
rect 1720 -140 1740 -120
rect 1760 -140 1780 -120
rect 1800 -140 1820 -120
rect 1840 -140 1860 -120
rect 1880 -140 1900 -120
rect 1920 -140 1940 -120
rect 1960 -140 1980 -120
rect 2000 -140 2020 -120
rect 2040 -140 2060 -120
rect 2080 -140 2100 -120
rect 2120 -140 2140 -120
rect 2160 -140 2180 -120
rect 2200 -140 2220 -120
rect 2240 -140 2260 -120
rect 2280 -140 2300 -120
rect 2320 -140 2340 -120
rect 2360 -140 2380 -120
rect 2400 -140 2420 -120
rect 2440 -140 2460 -120
rect 2480 -140 2500 -120
rect 2520 -140 2540 -120
rect 2560 -140 2580 -120
rect 2600 -140 2620 -120
rect 2640 -140 2660 -120
rect 2680 -140 2700 -120
rect 2720 -140 2740 -120
rect 2760 -140 2780 -120
rect 2800 -140 2820 -120
rect 2840 -140 2860 -120
rect 2880 -140 2900 -120
rect 2920 -140 2940 -120
rect 2960 -140 2980 -120
rect 3000 -140 3020 -120
rect 3040 -140 3060 -120
rect 3080 -140 3100 -120
rect 3120 -140 3140 -120
rect 3160 -140 3180 -120
rect 3200 -140 3220 -120
rect 3240 -140 3260 -120
rect 3280 -140 3300 -120
rect 3320 -140 3340 -120
rect 3360 -140 3380 -120
rect 3400 -140 3420 -120
rect 3440 -140 3460 -120
rect 3480 -140 3500 -120
rect 3520 -140 3540 -120
rect 3560 -140 3580 -120
rect 3600 -140 3615 -120
rect -3485 -150 3615 -140
rect -3485 -1200 3615 -1190
rect -3485 -1220 -3470 -1200
rect -3450 -1220 -3430 -1200
rect -3410 -1220 -3390 -1200
rect -3370 -1220 -3350 -1200
rect -3330 -1220 -3310 -1200
rect -3290 -1220 -3270 -1200
rect -3250 -1220 -3230 -1200
rect -3210 -1220 -3190 -1200
rect -3170 -1220 -3150 -1200
rect -3130 -1220 -3110 -1200
rect -3090 -1220 -3070 -1200
rect -3050 -1220 -3030 -1200
rect -3010 -1220 -2990 -1200
rect -2970 -1220 -2950 -1200
rect -2930 -1220 -2910 -1200
rect -2890 -1220 -2870 -1200
rect -2850 -1220 -2830 -1200
rect -2810 -1220 -2790 -1200
rect -2770 -1220 -2750 -1200
rect -2730 -1220 -2710 -1200
rect -2690 -1220 -2670 -1200
rect -2650 -1220 -2630 -1200
rect -2610 -1220 -2590 -1200
rect -2570 -1220 -2550 -1200
rect -2530 -1220 -2510 -1200
rect -2490 -1220 -2470 -1200
rect -2450 -1220 -2430 -1200
rect -2410 -1220 -2390 -1200
rect -2370 -1220 -2350 -1200
rect -2330 -1220 -2310 -1200
rect -2290 -1220 -2270 -1200
rect -2250 -1220 -2230 -1200
rect -2210 -1220 -2190 -1200
rect -2170 -1220 -2150 -1200
rect -2130 -1220 -2110 -1200
rect -2090 -1220 -2070 -1200
rect -2050 -1220 -2030 -1200
rect -2010 -1220 -1990 -1200
rect -1970 -1220 -1950 -1200
rect -1930 -1220 -1910 -1200
rect -1890 -1220 -1870 -1200
rect -1850 -1220 -1830 -1200
rect -1810 -1220 -1790 -1200
rect -1770 -1220 -1750 -1200
rect -1730 -1220 -1710 -1200
rect -1690 -1220 -1670 -1200
rect -1650 -1220 -1630 -1200
rect -1610 -1220 -1590 -1200
rect -1570 -1220 -1550 -1200
rect -1530 -1220 -1510 -1200
rect -1490 -1220 -1470 -1200
rect -1450 -1220 -1430 -1200
rect -1410 -1220 -1390 -1200
rect -1370 -1220 -1350 -1200
rect -1330 -1220 -1310 -1200
rect -1290 -1220 -1270 -1200
rect -1250 -1220 -1230 -1200
rect -1210 -1220 -1190 -1200
rect -1170 -1220 -1150 -1200
rect -1130 -1220 -1110 -1200
rect -1090 -1220 -1070 -1200
rect -1050 -1220 -1030 -1200
rect -1010 -1220 -990 -1200
rect -970 -1220 -950 -1200
rect -930 -1220 -910 -1200
rect -890 -1220 -870 -1200
rect -850 -1220 -830 -1200
rect -810 -1220 -790 -1200
rect -770 -1220 -750 -1200
rect -730 -1220 -710 -1200
rect -690 -1220 -670 -1200
rect -650 -1220 -630 -1200
rect -610 -1220 -590 -1200
rect -570 -1220 -550 -1200
rect -530 -1220 -510 -1200
rect -490 -1220 -470 -1200
rect -450 -1220 -430 -1200
rect -410 -1220 -390 -1200
rect -370 -1220 -350 -1200
rect -330 -1220 -310 -1200
rect -290 -1220 -270 -1200
rect -250 -1220 -230 -1200
rect -210 -1220 -190 -1200
rect -170 -1220 -150 -1200
rect -130 -1220 -110 -1200
rect -90 -1220 -70 -1200
rect -50 -1220 -30 -1200
rect -10 -1220 10 -1200
rect 30 -1220 50 -1200
rect 80 -1220 100 -1200
rect 120 -1220 140 -1200
rect 160 -1220 180 -1200
rect 200 -1220 220 -1200
rect 240 -1220 260 -1200
rect 280 -1220 300 -1200
rect 320 -1220 340 -1200
rect 360 -1220 380 -1200
rect 400 -1220 420 -1200
rect 440 -1220 460 -1200
rect 480 -1220 500 -1200
rect 520 -1220 540 -1200
rect 560 -1220 580 -1200
rect 600 -1220 620 -1200
rect 640 -1220 660 -1200
rect 680 -1220 700 -1200
rect 720 -1220 740 -1200
rect 760 -1220 780 -1200
rect 800 -1220 820 -1200
rect 840 -1220 860 -1200
rect 880 -1220 900 -1200
rect 920 -1220 940 -1200
rect 960 -1220 980 -1200
rect 1000 -1220 1020 -1200
rect 1040 -1220 1060 -1200
rect 1080 -1220 1100 -1200
rect 1120 -1220 1140 -1200
rect 1160 -1220 1180 -1200
rect 1200 -1220 1220 -1200
rect 1240 -1220 1260 -1200
rect 1280 -1220 1300 -1200
rect 1320 -1220 1340 -1200
rect 1360 -1220 1380 -1200
rect 1400 -1220 1420 -1200
rect 1440 -1220 1460 -1200
rect 1480 -1220 1500 -1200
rect 1520 -1220 1540 -1200
rect 1560 -1220 1580 -1200
rect 1600 -1220 1620 -1200
rect 1640 -1220 1660 -1200
rect 1680 -1220 1700 -1200
rect 1720 -1220 1740 -1200
rect 1760 -1220 1780 -1200
rect 1800 -1220 1820 -1200
rect 1840 -1220 1860 -1200
rect 1880 -1220 1900 -1200
rect 1920 -1220 1940 -1200
rect 1960 -1220 1980 -1200
rect 2000 -1220 2020 -1200
rect 2040 -1220 2060 -1200
rect 2080 -1220 2100 -1200
rect 2120 -1220 2140 -1200
rect 2160 -1220 2180 -1200
rect 2200 -1220 2220 -1200
rect 2240 -1220 2260 -1200
rect 2280 -1220 2300 -1200
rect 2320 -1220 2340 -1200
rect 2360 -1220 2380 -1200
rect 2400 -1220 2420 -1200
rect 2440 -1220 2460 -1200
rect 2480 -1220 2500 -1200
rect 2520 -1220 2540 -1200
rect 2560 -1220 2580 -1200
rect 2600 -1220 2620 -1200
rect 2640 -1220 2660 -1200
rect 2680 -1220 2700 -1200
rect 2720 -1220 2740 -1200
rect 2760 -1220 2780 -1200
rect 2800 -1220 2820 -1200
rect 2840 -1220 2860 -1200
rect 2880 -1220 2900 -1200
rect 2920 -1220 2940 -1200
rect 2960 -1220 2980 -1200
rect 3000 -1220 3020 -1200
rect 3040 -1220 3060 -1200
rect 3080 -1220 3100 -1200
rect 3120 -1220 3140 -1200
rect 3160 -1220 3180 -1200
rect 3200 -1220 3220 -1200
rect 3240 -1220 3260 -1200
rect 3280 -1220 3300 -1200
rect 3320 -1220 3340 -1200
rect 3360 -1220 3380 -1200
rect 3400 -1220 3420 -1200
rect 3440 -1220 3460 -1200
rect 3480 -1220 3500 -1200
rect 3520 -1220 3540 -1200
rect 3560 -1220 3580 -1200
rect 3600 -1220 3615 -1200
rect -3485 -1230 3615 -1220
<< psubdiffcont >>
rect -3470 -140 -3450 -120
rect -3430 -140 -3410 -120
rect -3390 -140 -3370 -120
rect -3350 -140 -3330 -120
rect -3310 -140 -3290 -120
rect -3270 -140 -3250 -120
rect -3230 -140 -3210 -120
rect -3190 -140 -3170 -120
rect -3150 -140 -3130 -120
rect -3110 -140 -3090 -120
rect -3070 -140 -3050 -120
rect -3030 -140 -3010 -120
rect -2990 -140 -2970 -120
rect -2950 -140 -2930 -120
rect -2910 -140 -2890 -120
rect -2870 -140 -2850 -120
rect -2830 -140 -2810 -120
rect -2790 -140 -2770 -120
rect -2750 -140 -2730 -120
rect -2710 -140 -2690 -120
rect -2670 -140 -2650 -120
rect -2630 -140 -2610 -120
rect -2590 -140 -2570 -120
rect -2550 -140 -2530 -120
rect -2510 -140 -2490 -120
rect -2470 -140 -2450 -120
rect -2430 -140 -2410 -120
rect -2390 -140 -2370 -120
rect -2350 -140 -2330 -120
rect -2310 -140 -2290 -120
rect -2270 -140 -2250 -120
rect -2230 -140 -2210 -120
rect -2190 -140 -2170 -120
rect -2150 -140 -2130 -120
rect -2110 -140 -2090 -120
rect -2070 -140 -2050 -120
rect -2030 -140 -2010 -120
rect -1990 -140 -1970 -120
rect -1950 -140 -1930 -120
rect -1910 -140 -1890 -120
rect -1870 -140 -1850 -120
rect -1830 -140 -1810 -120
rect -1790 -140 -1770 -120
rect -1750 -140 -1730 -120
rect -1710 -140 -1690 -120
rect -1670 -140 -1650 -120
rect -1630 -140 -1610 -120
rect -1590 -140 -1570 -120
rect -1550 -140 -1530 -120
rect -1510 -140 -1460 -120
rect -1440 -140 -1420 -120
rect -1400 -140 -1380 -120
rect -1360 -140 -1340 -120
rect -1320 -140 -1300 -120
rect -1280 -140 -1260 -120
rect -1240 -140 -1220 -120
rect -1200 -140 -1180 -120
rect -1160 -140 -1140 -120
rect -1120 -140 -1100 -120
rect -1080 -140 -1060 -120
rect -1040 -140 -1020 -120
rect -1000 -140 -980 -120
rect -960 -140 -940 -120
rect -920 -140 -900 -120
rect -880 -140 -860 -120
rect -840 -140 -820 -120
rect -800 -140 -780 -120
rect -760 -140 -740 -120
rect -720 -140 -700 -120
rect -680 -140 -660 -120
rect -640 -140 -620 -120
rect -600 -140 -580 -120
rect -560 -140 -540 -120
rect -520 -140 -500 -120
rect -480 -140 -460 -120
rect -440 -140 -420 -120
rect -400 -140 -380 -120
rect -360 -140 -340 -120
rect -320 -140 -300 -120
rect -280 -140 -260 -120
rect -230 -140 -210 -120
rect -190 -140 -170 -120
rect -150 -140 -130 -120
rect -110 -140 -90 -120
rect -70 -140 -50 -120
rect -30 -140 -10 -120
rect 10 -140 30 -120
rect 50 -140 80 -120
rect 100 -140 120 -120
rect 140 -140 160 -120
rect 180 -140 200 -120
rect 220 -140 240 -120
rect 260 -140 280 -120
rect 300 -140 320 -120
rect 340 -140 360 -120
rect 390 -140 410 -120
rect 430 -140 450 -120
rect 470 -140 490 -120
rect 510 -140 530 -120
rect 550 -140 570 -120
rect 590 -140 610 -120
rect 630 -140 650 -120
rect 670 -140 690 -120
rect 710 -140 730 -120
rect 750 -140 770 -120
rect 790 -140 810 -120
rect 830 -140 850 -120
rect 870 -140 890 -120
rect 910 -140 930 -120
rect 950 -140 970 -120
rect 990 -140 1010 -120
rect 1030 -140 1050 -120
rect 1070 -140 1090 -120
rect 1110 -140 1130 -120
rect 1150 -140 1170 -120
rect 1190 -140 1210 -120
rect 1230 -140 1250 -120
rect 1270 -140 1290 -120
rect 1310 -140 1330 -120
rect 1350 -140 1370 -120
rect 1390 -140 1410 -120
rect 1430 -140 1450 -120
rect 1470 -140 1490 -120
rect 1510 -140 1530 -120
rect 1550 -140 1570 -120
rect 1590 -140 1640 -120
rect 1660 -140 1680 -120
rect 1700 -140 1720 -120
rect 1740 -140 1760 -120
rect 1780 -140 1800 -120
rect 1820 -140 1840 -120
rect 1860 -140 1880 -120
rect 1900 -140 1920 -120
rect 1940 -140 1960 -120
rect 1980 -140 2000 -120
rect 2020 -140 2040 -120
rect 2060 -140 2080 -120
rect 2100 -140 2120 -120
rect 2140 -140 2160 -120
rect 2180 -140 2200 -120
rect 2220 -140 2240 -120
rect 2260 -140 2280 -120
rect 2300 -140 2320 -120
rect 2340 -140 2360 -120
rect 2380 -140 2400 -120
rect 2420 -140 2440 -120
rect 2460 -140 2480 -120
rect 2500 -140 2520 -120
rect 2540 -140 2560 -120
rect 2580 -140 2600 -120
rect 2620 -140 2640 -120
rect 2660 -140 2680 -120
rect 2700 -140 2720 -120
rect 2740 -140 2760 -120
rect 2780 -140 2800 -120
rect 2820 -140 2840 -120
rect 2860 -140 2880 -120
rect 2900 -140 2920 -120
rect 2940 -140 2960 -120
rect 2980 -140 3000 -120
rect 3020 -140 3040 -120
rect 3060 -140 3080 -120
rect 3100 -140 3120 -120
rect 3140 -140 3160 -120
rect 3180 -140 3200 -120
rect 3220 -140 3240 -120
rect 3260 -140 3280 -120
rect 3300 -140 3320 -120
rect 3340 -140 3360 -120
rect 3380 -140 3400 -120
rect 3420 -140 3440 -120
rect 3460 -140 3480 -120
rect 3500 -140 3520 -120
rect 3540 -140 3560 -120
rect 3580 -140 3600 -120
rect -3470 -1220 -3450 -1200
rect -3430 -1220 -3410 -1200
rect -3390 -1220 -3370 -1200
rect -3350 -1220 -3330 -1200
rect -3310 -1220 -3290 -1200
rect -3270 -1220 -3250 -1200
rect -3230 -1220 -3210 -1200
rect -3190 -1220 -3170 -1200
rect -3150 -1220 -3130 -1200
rect -3110 -1220 -3090 -1200
rect -3070 -1220 -3050 -1200
rect -3030 -1220 -3010 -1200
rect -2990 -1220 -2970 -1200
rect -2950 -1220 -2930 -1200
rect -2910 -1220 -2890 -1200
rect -2870 -1220 -2850 -1200
rect -2830 -1220 -2810 -1200
rect -2790 -1220 -2770 -1200
rect -2750 -1220 -2730 -1200
rect -2710 -1220 -2690 -1200
rect -2670 -1220 -2650 -1200
rect -2630 -1220 -2610 -1200
rect -2590 -1220 -2570 -1200
rect -2550 -1220 -2530 -1200
rect -2510 -1220 -2490 -1200
rect -2470 -1220 -2450 -1200
rect -2430 -1220 -2410 -1200
rect -2390 -1220 -2370 -1200
rect -2350 -1220 -2330 -1200
rect -2310 -1220 -2290 -1200
rect -2270 -1220 -2250 -1200
rect -2230 -1220 -2210 -1200
rect -2190 -1220 -2170 -1200
rect -2150 -1220 -2130 -1200
rect -2110 -1220 -2090 -1200
rect -2070 -1220 -2050 -1200
rect -2030 -1220 -2010 -1200
rect -1990 -1220 -1970 -1200
rect -1950 -1220 -1930 -1200
rect -1910 -1220 -1890 -1200
rect -1870 -1220 -1850 -1200
rect -1830 -1220 -1810 -1200
rect -1790 -1220 -1770 -1200
rect -1750 -1220 -1730 -1200
rect -1710 -1220 -1690 -1200
rect -1670 -1220 -1650 -1200
rect -1630 -1220 -1610 -1200
rect -1590 -1220 -1570 -1200
rect -1550 -1220 -1530 -1200
rect -1510 -1220 -1490 -1200
rect -1470 -1220 -1450 -1200
rect -1430 -1220 -1410 -1200
rect -1390 -1220 -1370 -1200
rect -1350 -1220 -1330 -1200
rect -1310 -1220 -1290 -1200
rect -1270 -1220 -1250 -1200
rect -1230 -1220 -1210 -1200
rect -1190 -1220 -1170 -1200
rect -1150 -1220 -1130 -1200
rect -1110 -1220 -1090 -1200
rect -1070 -1220 -1050 -1200
rect -1030 -1220 -1010 -1200
rect -990 -1220 -970 -1200
rect -950 -1220 -930 -1200
rect -910 -1220 -890 -1200
rect -870 -1220 -850 -1200
rect -830 -1220 -810 -1200
rect -790 -1220 -770 -1200
rect -750 -1220 -730 -1200
rect -710 -1220 -690 -1200
rect -670 -1220 -650 -1200
rect -630 -1220 -610 -1200
rect -590 -1220 -570 -1200
rect -550 -1220 -530 -1200
rect -510 -1220 -490 -1200
rect -470 -1220 -450 -1200
rect -430 -1220 -410 -1200
rect -390 -1220 -370 -1200
rect -350 -1220 -330 -1200
rect -310 -1220 -290 -1200
rect -270 -1220 -250 -1200
rect -230 -1220 -210 -1200
rect -190 -1220 -170 -1200
rect -150 -1220 -130 -1200
rect -110 -1220 -90 -1200
rect -70 -1220 -50 -1200
rect -30 -1220 -10 -1200
rect 10 -1220 30 -1200
rect 50 -1220 80 -1200
rect 100 -1220 120 -1200
rect 140 -1220 160 -1200
rect 180 -1220 200 -1200
rect 220 -1220 240 -1200
rect 260 -1220 280 -1200
rect 300 -1220 320 -1200
rect 340 -1220 360 -1200
rect 380 -1220 400 -1200
rect 420 -1220 440 -1200
rect 460 -1220 480 -1200
rect 500 -1220 520 -1200
rect 540 -1220 560 -1200
rect 580 -1220 600 -1200
rect 620 -1220 640 -1200
rect 660 -1220 680 -1200
rect 700 -1220 720 -1200
rect 740 -1220 760 -1200
rect 780 -1220 800 -1200
rect 820 -1220 840 -1200
rect 860 -1220 880 -1200
rect 900 -1220 920 -1200
rect 940 -1220 960 -1200
rect 980 -1220 1000 -1200
rect 1020 -1220 1040 -1200
rect 1060 -1220 1080 -1200
rect 1100 -1220 1120 -1200
rect 1140 -1220 1160 -1200
rect 1180 -1220 1200 -1200
rect 1220 -1220 1240 -1200
rect 1260 -1220 1280 -1200
rect 1300 -1220 1320 -1200
rect 1340 -1220 1360 -1200
rect 1380 -1220 1400 -1200
rect 1420 -1220 1440 -1200
rect 1460 -1220 1480 -1200
rect 1500 -1220 1520 -1200
rect 1540 -1220 1560 -1200
rect 1580 -1220 1600 -1200
rect 1620 -1220 1640 -1200
rect 1660 -1220 1680 -1200
rect 1700 -1220 1720 -1200
rect 1740 -1220 1760 -1200
rect 1780 -1220 1800 -1200
rect 1820 -1220 1840 -1200
rect 1860 -1220 1880 -1200
rect 1900 -1220 1920 -1200
rect 1940 -1220 1960 -1200
rect 1980 -1220 2000 -1200
rect 2020 -1220 2040 -1200
rect 2060 -1220 2080 -1200
rect 2100 -1220 2120 -1200
rect 2140 -1220 2160 -1200
rect 2180 -1220 2200 -1200
rect 2220 -1220 2240 -1200
rect 2260 -1220 2280 -1200
rect 2300 -1220 2320 -1200
rect 2340 -1220 2360 -1200
rect 2380 -1220 2400 -1200
rect 2420 -1220 2440 -1200
rect 2460 -1220 2480 -1200
rect 2500 -1220 2520 -1200
rect 2540 -1220 2560 -1200
rect 2580 -1220 2600 -1200
rect 2620 -1220 2640 -1200
rect 2660 -1220 2680 -1200
rect 2700 -1220 2720 -1200
rect 2740 -1220 2760 -1200
rect 2780 -1220 2800 -1200
rect 2820 -1220 2840 -1200
rect 2860 -1220 2880 -1200
rect 2900 -1220 2920 -1200
rect 2940 -1220 2960 -1200
rect 2980 -1220 3000 -1200
rect 3020 -1220 3040 -1200
rect 3060 -1220 3080 -1200
rect 3100 -1220 3120 -1200
rect 3140 -1220 3160 -1200
rect 3180 -1220 3200 -1200
rect 3220 -1220 3240 -1200
rect 3260 -1220 3280 -1200
rect 3300 -1220 3320 -1200
rect 3340 -1220 3360 -1200
rect 3380 -1220 3400 -1200
rect 3420 -1220 3440 -1200
rect 3460 -1220 3480 -1200
rect 3500 -1220 3520 -1200
rect 3540 -1220 3560 -1200
rect 3580 -1220 3600 -1200
<< poly >>
rect -3500 -245 -3485 -195
rect 3615 -205 3790 -195
rect 3615 -235 3645 -205
rect 3665 -235 3685 -205
rect 3705 -235 3725 -205
rect 3745 -235 3765 -205
rect 3785 -235 3790 -205
rect 3615 -245 3790 -235
rect -3500 -345 -3485 -295
rect 3615 -305 3790 -295
rect 3615 -335 3645 -305
rect 3665 -335 3685 -305
rect 3705 -335 3725 -305
rect 3745 -335 3765 -305
rect 3785 -335 3790 -305
rect 3615 -345 3790 -335
rect -3500 -445 -3485 -395
rect 3615 -405 3790 -395
rect 3615 -435 3645 -405
rect 3665 -435 3685 -405
rect 3705 -435 3725 -405
rect 3745 -435 3765 -405
rect 3785 -435 3790 -405
rect 3615 -445 3790 -435
rect -3500 -545 -3485 -495
rect 3615 -505 3790 -495
rect 3615 -535 3645 -505
rect 3665 -535 3685 -505
rect 3705 -535 3725 -505
rect 3745 -535 3765 -505
rect 3785 -535 3790 -505
rect 3615 -545 3790 -535
rect -3500 -645 -3485 -595
rect 3615 -605 3790 -595
rect 3615 -635 3645 -605
rect 3665 -635 3685 -605
rect 3705 -635 3725 -605
rect 3745 -635 3765 -605
rect 3785 -635 3790 -605
rect 3615 -645 3790 -635
rect -3500 -745 -3485 -695
rect 3615 -705 3790 -695
rect 3615 -735 3645 -705
rect 3665 -735 3685 -705
rect 3705 -735 3725 -705
rect 3745 -735 3765 -705
rect 3785 -735 3790 -705
rect 3615 -745 3790 -735
rect -3500 -845 -3485 -795
rect 3615 -805 3790 -795
rect 3615 -835 3645 -805
rect 3665 -835 3685 -805
rect 3705 -835 3725 -805
rect 3745 -835 3765 -805
rect 3785 -835 3790 -805
rect 3615 -845 3790 -835
rect -3500 -945 -3485 -895
rect 3615 -905 3790 -895
rect 3615 -935 3645 -905
rect 3665 -935 3685 -905
rect 3705 -935 3725 -905
rect 3745 -935 3765 -905
rect 3785 -935 3790 -905
rect 3615 -945 3790 -935
rect -3500 -1045 -3485 -995
rect 3615 -1005 3790 -995
rect 3615 -1035 3645 -1005
rect 3665 -1035 3685 -1005
rect 3705 -1035 3725 -1005
rect 3745 -1035 3765 -1005
rect 3785 -1035 3790 -1005
rect 3615 -1045 3790 -1035
rect -3505 -1145 -3485 -1095
rect 3615 -1105 3790 -1095
rect 3615 -1135 3645 -1105
rect 3665 -1135 3685 -1105
rect 3705 -1135 3725 -1105
rect 3745 -1135 3765 -1105
rect 3785 -1135 3790 -1105
rect 3615 -1145 3790 -1135
<< polycont >>
rect 3645 -235 3665 -205
rect 3685 -235 3705 -205
rect 3725 -235 3745 -205
rect 3765 -235 3785 -205
rect 3645 -335 3665 -305
rect 3685 -335 3705 -305
rect 3725 -335 3745 -305
rect 3765 -335 3785 -305
rect 3645 -435 3665 -405
rect 3685 -435 3705 -405
rect 3725 -435 3745 -405
rect 3765 -435 3785 -405
rect 3645 -535 3665 -505
rect 3685 -535 3705 -505
rect 3725 -535 3745 -505
rect 3765 -535 3785 -505
rect 3645 -635 3665 -605
rect 3685 -635 3705 -605
rect 3725 -635 3745 -605
rect 3765 -635 3785 -605
rect 3645 -735 3665 -705
rect 3685 -735 3705 -705
rect 3725 -735 3745 -705
rect 3765 -735 3785 -705
rect 3645 -835 3665 -805
rect 3685 -835 3705 -805
rect 3725 -835 3745 -805
rect 3765 -835 3785 -805
rect 3645 -935 3665 -905
rect 3685 -935 3705 -905
rect 3725 -935 3745 -905
rect 3765 -935 3785 -905
rect 3645 -1035 3665 -1005
rect 3685 -1035 3705 -1005
rect 3725 -1035 3745 -1005
rect 3765 -1035 3785 -1005
rect 3645 -1135 3665 -1105
rect 3685 -1135 3705 -1105
rect 3725 -1135 3745 -1105
rect 3765 -1135 3785 -1105
<< locali >>
rect -3485 -120 3615 -110
rect -3485 -140 -3470 -120
rect -3450 -140 -3430 -120
rect -3410 -140 -3390 -120
rect -3370 -140 -3350 -120
rect -3330 -140 -3310 -120
rect -3290 -140 -3270 -120
rect -3250 -140 -3230 -120
rect -3210 -140 -3190 -120
rect -3170 -140 -3150 -120
rect -3130 -140 -3110 -120
rect -3090 -140 -3070 -120
rect -3050 -140 -3030 -120
rect -3010 -140 -2990 -120
rect -2970 -140 -2950 -120
rect -2930 -140 -2910 -120
rect -2890 -140 -2870 -120
rect -2850 -140 -2830 -120
rect -2810 -140 -2790 -120
rect -2770 -140 -2750 -120
rect -2730 -140 -2710 -120
rect -2690 -140 -2670 -120
rect -2650 -140 -2630 -120
rect -2610 -140 -2590 -120
rect -2570 -140 -2550 -120
rect -2530 -140 -2510 -120
rect -2490 -140 -2470 -120
rect -2450 -140 -2430 -120
rect -2410 -140 -2390 -120
rect -2370 -140 -2350 -120
rect -2330 -140 -2310 -120
rect -2290 -140 -2270 -120
rect -2250 -140 -2230 -120
rect -2210 -140 -2190 -120
rect -2170 -140 -2150 -120
rect -2130 -140 -2110 -120
rect -2090 -140 -2070 -120
rect -2050 -140 -2030 -120
rect -2010 -140 -1990 -120
rect -1970 -140 -1950 -120
rect -1930 -140 -1910 -120
rect -1890 -140 -1870 -120
rect -1850 -140 -1830 -120
rect -1810 -140 -1790 -120
rect -1770 -140 -1750 -120
rect -1730 -140 -1710 -120
rect -1690 -140 -1670 -120
rect -1650 -140 -1630 -120
rect -1610 -140 -1590 -120
rect -1570 -140 -1550 -120
rect -1530 -140 -1510 -120
rect -1460 -140 -1440 -120
rect -1420 -140 -1400 -120
rect -1380 -140 -1360 -120
rect -1340 -140 -1320 -120
rect -1300 -140 -1280 -120
rect -1260 -140 -1240 -120
rect -1220 -140 -1200 -120
rect -1180 -140 -1160 -120
rect -1140 -140 -1120 -120
rect -1100 -140 -1080 -120
rect -1060 -140 -1040 -120
rect -1020 -140 -1000 -120
rect -980 -140 -960 -120
rect -940 -140 -920 -120
rect -900 -140 -880 -120
rect -860 -140 -840 -120
rect -820 -140 -800 -120
rect -780 -140 -760 -120
rect -740 -140 -720 -120
rect -700 -140 -680 -120
rect -660 -140 -640 -120
rect -620 -140 -600 -120
rect -580 -140 -560 -120
rect -540 -140 -520 -120
rect -500 -140 -480 -120
rect -460 -140 -440 -120
rect -420 -140 -400 -120
rect -380 -140 -360 -120
rect -340 -140 -320 -120
rect -300 -140 -280 -120
rect -260 -140 -230 -120
rect -210 -140 -190 -120
rect -170 -140 -150 -120
rect -130 -140 -110 -120
rect -90 -140 -70 -120
rect -50 -140 -30 -120
rect -10 -140 10 -120
rect 30 -140 50 -120
rect 80 -140 100 -120
rect 120 -140 140 -120
rect 160 -140 180 -120
rect 200 -140 220 -120
rect 240 -140 260 -120
rect 280 -140 300 -120
rect 320 -140 340 -120
rect 360 -140 390 -120
rect 410 -140 430 -120
rect 450 -140 470 -120
rect 490 -140 510 -120
rect 530 -140 550 -120
rect 570 -140 590 -120
rect 610 -140 630 -120
rect 650 -140 670 -120
rect 690 -140 710 -120
rect 730 -140 750 -120
rect 770 -140 790 -120
rect 810 -140 830 -120
rect 850 -140 870 -120
rect 890 -140 910 -120
rect 930 -140 950 -120
rect 970 -140 990 -120
rect 1010 -140 1030 -120
rect 1050 -140 1070 -120
rect 1090 -140 1110 -120
rect 1130 -140 1150 -120
rect 1170 -140 1190 -120
rect 1210 -140 1230 -120
rect 1250 -140 1270 -120
rect 1290 -140 1310 -120
rect 1330 -140 1350 -120
rect 1370 -140 1390 -120
rect 1410 -140 1430 -120
rect 1450 -140 1470 -120
rect 1490 -140 1510 -120
rect 1530 -140 1550 -120
rect 1570 -140 1590 -120
rect 1640 -140 1660 -120
rect 1680 -140 1700 -120
rect 1720 -140 1740 -120
rect 1760 -140 1780 -120
rect 1800 -140 1820 -120
rect 1840 -140 1860 -120
rect 1880 -140 1900 -120
rect 1920 -140 1940 -120
rect 1960 -140 1980 -120
rect 2000 -140 2020 -120
rect 2040 -140 2060 -120
rect 2080 -140 2100 -120
rect 2120 -140 2140 -120
rect 2160 -140 2180 -120
rect 2200 -140 2220 -120
rect 2240 -140 2260 -120
rect 2280 -140 2300 -120
rect 2320 -140 2340 -120
rect 2360 -140 2380 -120
rect 2400 -140 2420 -120
rect 2440 -140 2460 -120
rect 2480 -140 2500 -120
rect 2520 -140 2540 -120
rect 2560 -140 2580 -120
rect 2600 -140 2620 -120
rect 2640 -140 2660 -120
rect 2680 -140 2700 -120
rect 2720 -140 2740 -120
rect 2760 -140 2780 -120
rect 2800 -140 2820 -120
rect 2840 -140 2860 -120
rect 2880 -140 2900 -120
rect 2920 -140 2940 -120
rect 2960 -140 2980 -120
rect 3000 -140 3020 -120
rect 3040 -140 3060 -120
rect 3080 -140 3100 -120
rect 3120 -140 3140 -120
rect 3160 -140 3180 -120
rect 3200 -140 3220 -120
rect 3240 -140 3260 -120
rect 3280 -140 3300 -120
rect 3320 -140 3340 -120
rect 3360 -140 3380 -120
rect 3400 -140 3420 -120
rect 3440 -140 3460 -120
rect 3480 -140 3500 -120
rect 3520 -140 3540 -120
rect 3560 -140 3580 -120
rect 3600 -140 3615 -120
rect -3485 -160 3615 -140
rect -3485 -180 -3470 -160
rect -3450 -180 -3430 -160
rect -3410 -180 -3390 -160
rect -3370 -180 -3350 -160
rect -3330 -180 -3310 -160
rect -3290 -180 -3270 -160
rect -3250 -180 -3230 -160
rect -3210 -180 -3190 -160
rect -3170 -180 -3150 -160
rect -3130 -180 -3110 -160
rect -3090 -180 -3070 -160
rect -3050 -180 -3030 -160
rect -3010 -180 -2990 -160
rect -2970 -180 -2950 -160
rect -2930 -180 -2910 -160
rect -2890 -180 -2870 -160
rect -2850 -180 -2830 -160
rect -2810 -180 -2790 -160
rect -2770 -180 -2750 -160
rect -2730 -180 -2710 -160
rect -2690 -180 -2670 -160
rect -2650 -180 -2630 -160
rect -2610 -180 -2590 -160
rect -2570 -180 -2550 -160
rect -2530 -180 -2510 -160
rect -2490 -180 -2470 -160
rect -2450 -180 -2430 -160
rect -2410 -180 -2390 -160
rect -2370 -180 -2350 -160
rect -2330 -180 -2310 -160
rect -2290 -180 -2270 -160
rect -2250 -180 -2230 -160
rect -2210 -180 -2190 -160
rect -2170 -180 -2150 -160
rect -2130 -180 -2110 -160
rect -2090 -180 -2070 -160
rect -2050 -180 -2030 -160
rect -2010 -180 -1990 -160
rect -1970 -180 -1950 -160
rect -1930 -180 -1910 -160
rect -1890 -180 -1870 -160
rect -1850 -180 -1830 -160
rect -1810 -180 -1790 -160
rect -1770 -180 -1750 -160
rect -1730 -180 -1710 -160
rect -1690 -180 -1670 -160
rect -1650 -180 -1630 -160
rect -1610 -180 -1590 -160
rect -1570 -180 -1550 -160
rect -1530 -180 -1510 -160
rect -1460 -180 -1440 -160
rect -1420 -180 -1400 -160
rect -1380 -180 -1360 -160
rect -1340 -180 -1320 -160
rect -1300 -180 -1280 -160
rect -1260 -180 -1240 -160
rect -1220 -180 -1200 -160
rect -1180 -180 -1160 -160
rect -1140 -180 -1120 -160
rect -1100 -180 -1080 -160
rect -1060 -180 -1040 -160
rect -1020 -180 -1000 -160
rect -980 -180 -960 -160
rect -940 -180 -920 -160
rect -900 -180 -880 -160
rect -860 -180 -840 -160
rect -820 -180 -800 -160
rect -780 -180 -760 -160
rect -740 -180 -720 -160
rect -700 -180 -680 -160
rect -660 -180 -640 -160
rect -620 -180 -600 -160
rect -580 -180 -560 -160
rect -540 -180 -520 -160
rect -500 -180 -480 -160
rect -460 -180 -440 -160
rect -420 -180 -400 -160
rect -380 -180 -360 -160
rect -340 -180 -320 -160
rect -300 -180 -280 -160
rect -260 -180 -230 -160
rect -210 -180 -190 -160
rect -170 -180 -150 -160
rect -130 -180 -110 -160
rect -90 -180 -70 -160
rect -50 -180 -30 -160
rect -10 -180 10 -160
rect 30 -180 50 -160
rect 80 -180 100 -160
rect 120 -180 140 -160
rect 160 -180 180 -160
rect 200 -180 220 -160
rect 240 -180 260 -160
rect 280 -180 300 -160
rect 320 -180 340 -160
rect 360 -180 390 -160
rect 410 -180 430 -160
rect 450 -180 470 -160
rect 490 -180 510 -160
rect 530 -180 550 -160
rect 570 -180 590 -160
rect 610 -180 630 -160
rect 650 -180 670 -160
rect 690 -180 710 -160
rect 730 -180 750 -160
rect 770 -180 790 -160
rect 810 -180 830 -160
rect 850 -180 870 -160
rect 890 -180 910 -160
rect 930 -180 950 -160
rect 970 -180 990 -160
rect 1010 -180 1030 -160
rect 1050 -180 1070 -160
rect 1090 -180 1110 -160
rect 1130 -180 1150 -160
rect 1170 -180 1190 -160
rect 1210 -180 1230 -160
rect 1250 -180 1270 -160
rect 1290 -180 1310 -160
rect 1330 -180 1350 -160
rect 1370 -180 1390 -160
rect 1410 -180 1430 -160
rect 1450 -180 1470 -160
rect 1490 -180 1510 -160
rect 1530 -180 1550 -160
rect 1570 -180 1590 -160
rect 1640 -180 1660 -160
rect 1680 -180 1700 -160
rect 1720 -180 1740 -160
rect 1760 -180 1780 -160
rect 1800 -180 1820 -160
rect 1840 -180 1860 -160
rect 1880 -180 1900 -160
rect 1920 -180 1940 -160
rect 1960 -180 1980 -160
rect 2000 -180 2020 -160
rect 2040 -180 2060 -160
rect 2080 -180 2100 -160
rect 2120 -180 2140 -160
rect 2160 -180 2180 -160
rect 2200 -180 2220 -160
rect 2240 -180 2260 -160
rect 2280 -180 2300 -160
rect 2320 -180 2340 -160
rect 2360 -180 2380 -160
rect 2400 -180 2420 -160
rect 2440 -180 2460 -160
rect 2480 -180 2500 -160
rect 2520 -180 2540 -160
rect 2560 -180 2580 -160
rect 2600 -180 2620 -160
rect 2640 -180 2660 -160
rect 2680 -180 2700 -160
rect 2720 -180 2740 -160
rect 2760 -180 2780 -160
rect 2800 -180 2820 -160
rect 2840 -180 2860 -160
rect 2880 -180 2900 -160
rect 2920 -180 2940 -160
rect 2960 -180 2980 -160
rect 3000 -180 3020 -160
rect 3040 -180 3060 -160
rect 3080 -180 3100 -160
rect 3120 -180 3140 -160
rect 3160 -180 3180 -160
rect 3200 -180 3220 -160
rect 3240 -180 3260 -160
rect 3280 -180 3300 -160
rect 3320 -180 3340 -160
rect 3360 -180 3380 -160
rect 3400 -180 3420 -160
rect 3440 -180 3460 -160
rect 3480 -180 3500 -160
rect 3520 -180 3540 -160
rect 3560 -180 3580 -160
rect 3600 -180 3615 -160
rect -3485 -190 3615 -180
rect 3635 -205 3790 -195
rect 3635 -235 3645 -205
rect 3665 -235 3685 -205
rect 3705 -235 3725 -205
rect 3745 -235 3765 -205
rect 3785 -235 3790 -205
rect 3635 -245 3790 -235
rect -3485 -260 3615 -250
rect -3485 -280 -3470 -260
rect -3450 -280 -3430 -260
rect -3410 -280 -3390 -260
rect -3370 -280 -3350 -260
rect -3330 -280 -3310 -260
rect -3290 -280 -3270 -260
rect -3250 -280 -3230 -260
rect -3210 -280 -3190 -260
rect -3170 -280 -3150 -260
rect -3130 -280 -3110 -260
rect -3090 -280 -3070 -260
rect -3050 -280 -3030 -260
rect -3010 -280 -2990 -260
rect -2970 -280 -2950 -260
rect -2930 -280 -2910 -260
rect -2890 -280 -2870 -260
rect -2850 -280 -2830 -260
rect -2810 -280 -2790 -260
rect -2770 -280 -2750 -260
rect -2730 -280 -2710 -260
rect -2690 -280 -2670 -260
rect -2650 -280 -2630 -260
rect -2610 -280 -2590 -260
rect -2570 -280 -2550 -260
rect -2530 -280 -2510 -260
rect -2490 -280 -2470 -260
rect -2450 -280 -2430 -260
rect -2410 -280 -2390 -260
rect -2370 -280 -2350 -260
rect -2330 -280 -2310 -260
rect -2290 -280 -2270 -260
rect -2250 -280 -2230 -260
rect -2210 -280 -2190 -260
rect -2170 -280 -2150 -260
rect -2130 -280 -2110 -260
rect -2090 -280 -2070 -260
rect -2050 -280 -2030 -260
rect -2010 -280 -1990 -260
rect -1970 -280 -1950 -260
rect -1930 -280 -1910 -260
rect -1890 -280 -1870 -260
rect -1850 -280 -1830 -260
rect -1810 -280 -1790 -260
rect -1770 -280 -1750 -260
rect -1730 -280 -1710 -260
rect -1690 -280 -1670 -260
rect -1650 -280 -1630 -260
rect -1610 -280 -1590 -260
rect -1570 -280 -1550 -260
rect -1530 -280 -1510 -260
rect -1460 -280 -1440 -260
rect -1420 -280 -1400 -260
rect -1380 -280 -1360 -260
rect -1340 -280 -1320 -260
rect -1300 -280 -1280 -260
rect -1260 -280 -1240 -260
rect -1220 -280 -1200 -260
rect -1180 -280 -1160 -260
rect -1140 -280 -1120 -260
rect -1100 -280 -1080 -260
rect -1060 -280 -1040 -260
rect -1020 -280 -1000 -260
rect -980 -280 -960 -260
rect -940 -280 -920 -260
rect -900 -280 -880 -260
rect -860 -280 -840 -260
rect -820 -280 -800 -260
rect -780 -280 -760 -260
rect -740 -280 -720 -260
rect -700 -280 -680 -260
rect -660 -280 -640 -260
rect -620 -280 -600 -260
rect -580 -280 -560 -260
rect -540 -280 -520 -260
rect -500 -280 -480 -260
rect -460 -280 -440 -260
rect -420 -280 -400 -260
rect -380 -280 -360 -260
rect -340 -280 -320 -260
rect -300 -280 -280 -260
rect -260 -280 -230 -260
rect -210 -280 -190 -260
rect -170 -280 -150 -260
rect -130 -280 -110 -260
rect -90 -280 -70 -260
rect -50 -280 -30 -260
rect -10 -280 10 -260
rect 30 -280 50 -260
rect 80 -280 100 -260
rect 120 -280 140 -260
rect 160 -280 180 -260
rect 200 -280 220 -260
rect 240 -280 260 -260
rect 280 -280 300 -260
rect 320 -280 340 -260
rect 360 -280 390 -260
rect 410 -280 430 -260
rect 450 -280 470 -260
rect 490 -280 510 -260
rect 530 -280 550 -260
rect 570 -280 590 -260
rect 610 -280 630 -260
rect 650 -280 670 -260
rect 690 -280 710 -260
rect 730 -280 750 -260
rect 770 -280 790 -260
rect 810 -280 830 -260
rect 850 -280 870 -260
rect 890 -280 910 -260
rect 930 -280 950 -260
rect 970 -280 990 -260
rect 1010 -280 1030 -260
rect 1050 -280 1070 -260
rect 1090 -280 1110 -260
rect 1130 -280 1150 -260
rect 1170 -280 1190 -260
rect 1210 -280 1230 -260
rect 1250 -280 1270 -260
rect 1290 -280 1310 -260
rect 1330 -280 1350 -260
rect 1370 -280 1390 -260
rect 1410 -280 1430 -260
rect 1450 -280 1470 -260
rect 1490 -280 1510 -260
rect 1530 -280 1550 -260
rect 1570 -280 1590 -260
rect 1640 -280 1660 -260
rect 1680 -280 1700 -260
rect 1720 -280 1740 -260
rect 1760 -280 1780 -260
rect 1800 -280 1820 -260
rect 1840 -280 1860 -260
rect 1880 -280 1900 -260
rect 1920 -280 1940 -260
rect 1960 -280 1980 -260
rect 2000 -280 2020 -260
rect 2040 -280 2060 -260
rect 2080 -280 2100 -260
rect 2120 -280 2140 -260
rect 2160 -280 2180 -260
rect 2200 -280 2220 -260
rect 2240 -280 2260 -260
rect 2280 -280 2300 -260
rect 2320 -280 2340 -260
rect 2360 -280 2380 -260
rect 2400 -280 2420 -260
rect 2440 -280 2460 -260
rect 2480 -280 2500 -260
rect 2520 -280 2540 -260
rect 2560 -280 2580 -260
rect 2600 -280 2620 -260
rect 2640 -280 2660 -260
rect 2680 -280 2700 -260
rect 2720 -280 2740 -260
rect 2760 -280 2780 -260
rect 2800 -280 2820 -260
rect 2840 -280 2860 -260
rect 2880 -280 2900 -260
rect 2920 -280 2940 -260
rect 2960 -280 2980 -260
rect 3000 -280 3020 -260
rect 3040 -280 3060 -260
rect 3080 -280 3100 -260
rect 3120 -280 3140 -260
rect 3160 -280 3180 -260
rect 3200 -280 3220 -260
rect 3240 -280 3260 -260
rect 3280 -280 3300 -260
rect 3320 -280 3340 -260
rect 3360 -280 3380 -260
rect 3400 -280 3420 -260
rect 3440 -280 3460 -260
rect 3480 -280 3500 -260
rect 3520 -280 3540 -260
rect 3560 -280 3580 -260
rect 3600 -280 3615 -260
rect -3485 -290 3615 -280
rect 3635 -305 3790 -295
rect 3635 -335 3645 -305
rect 3665 -335 3685 -305
rect 3705 -335 3725 -305
rect 3745 -335 3765 -305
rect 3785 -335 3790 -305
rect 3635 -345 3790 -335
rect -3485 -360 3615 -350
rect -3485 -380 -3470 -360
rect -3450 -380 -3430 -360
rect -3410 -380 -3390 -360
rect -3370 -380 -3350 -360
rect -3330 -380 -3310 -360
rect -3290 -380 -3270 -360
rect -3250 -380 -3230 -360
rect -3210 -380 -3190 -360
rect -3170 -380 -3150 -360
rect -3130 -380 -3110 -360
rect -3090 -380 -3070 -360
rect -3050 -380 -3030 -360
rect -3010 -380 -2990 -360
rect -2970 -380 -2950 -360
rect -2930 -380 -2910 -360
rect -2890 -380 -2870 -360
rect -2850 -380 -2830 -360
rect -2810 -380 -2790 -360
rect -2770 -380 -2750 -360
rect -2730 -380 -2710 -360
rect -2690 -380 -2670 -360
rect -2650 -380 -2630 -360
rect -2610 -380 -2590 -360
rect -2570 -380 -2550 -360
rect -2530 -380 -2510 -360
rect -2490 -380 -2470 -360
rect -2450 -380 -2430 -360
rect -2410 -380 -2390 -360
rect -2370 -380 -2350 -360
rect -2330 -380 -2310 -360
rect -2290 -380 -2270 -360
rect -2250 -380 -2230 -360
rect -2210 -380 -2190 -360
rect -2170 -380 -2150 -360
rect -2130 -380 -2110 -360
rect -2090 -380 -2070 -360
rect -2050 -380 -2030 -360
rect -2010 -380 -1990 -360
rect -1970 -380 -1950 -360
rect -1930 -380 -1910 -360
rect -1890 -380 -1870 -360
rect -1850 -380 -1830 -360
rect -1810 -380 -1790 -360
rect -1770 -380 -1750 -360
rect -1730 -380 -1710 -360
rect -1690 -380 -1670 -360
rect -1650 -380 -1630 -360
rect -1610 -380 -1590 -360
rect -1570 -380 -1550 -360
rect -1530 -380 -1510 -360
rect -1460 -380 -1440 -360
rect -1420 -380 -1400 -360
rect -1380 -380 -1360 -360
rect -1340 -380 -1320 -360
rect -1300 -380 -1280 -360
rect -1260 -380 -1240 -360
rect -1220 -380 -1200 -360
rect -1180 -380 -1160 -360
rect -1140 -380 -1120 -360
rect -1100 -380 -1080 -360
rect -1060 -380 -1040 -360
rect -1020 -380 -1000 -360
rect -980 -380 -960 -360
rect -940 -380 -920 -360
rect -900 -380 -880 -360
rect -860 -380 -840 -360
rect -820 -380 -800 -360
rect -780 -380 -760 -360
rect -740 -380 -720 -360
rect -700 -380 -680 -360
rect -660 -380 -640 -360
rect -620 -380 -600 -360
rect -580 -380 -560 -360
rect -540 -380 -520 -360
rect -500 -380 -480 -360
rect -460 -380 -440 -360
rect -420 -380 -400 -360
rect -380 -380 -360 -360
rect -340 -380 -320 -360
rect -300 -380 -280 -360
rect -260 -380 -230 -360
rect -210 -380 -190 -360
rect -170 -380 -150 -360
rect -130 -380 -110 -360
rect -90 -380 -70 -360
rect -50 -380 -30 -360
rect -10 -380 10 -360
rect 30 -380 50 -360
rect 80 -380 100 -360
rect 120 -380 140 -360
rect 160 -380 180 -360
rect 200 -380 220 -360
rect 240 -380 260 -360
rect 280 -380 300 -360
rect 320 -380 340 -360
rect 360 -380 390 -360
rect 410 -380 430 -360
rect 450 -380 470 -360
rect 490 -380 510 -360
rect 530 -380 550 -360
rect 570 -380 590 -360
rect 610 -380 630 -360
rect 650 -380 670 -360
rect 690 -380 710 -360
rect 730 -380 750 -360
rect 770 -380 790 -360
rect 810 -380 830 -360
rect 850 -380 870 -360
rect 890 -380 910 -360
rect 930 -380 950 -360
rect 970 -380 990 -360
rect 1010 -380 1030 -360
rect 1050 -380 1070 -360
rect 1090 -380 1110 -360
rect 1130 -380 1150 -360
rect 1170 -380 1190 -360
rect 1210 -380 1230 -360
rect 1250 -380 1270 -360
rect 1290 -380 1310 -360
rect 1330 -380 1350 -360
rect 1370 -380 1390 -360
rect 1410 -380 1430 -360
rect 1450 -380 1470 -360
rect 1490 -380 1510 -360
rect 1530 -380 1550 -360
rect 1570 -380 1590 -360
rect 1640 -380 1660 -360
rect 1680 -380 1700 -360
rect 1720 -380 1740 -360
rect 1760 -380 1780 -360
rect 1800 -380 1820 -360
rect 1840 -380 1860 -360
rect 1880 -380 1900 -360
rect 1920 -380 1940 -360
rect 1960 -380 1980 -360
rect 2000 -380 2020 -360
rect 2040 -380 2060 -360
rect 2080 -380 2100 -360
rect 2120 -380 2140 -360
rect 2160 -380 2180 -360
rect 2200 -380 2220 -360
rect 2240 -380 2260 -360
rect 2280 -380 2300 -360
rect 2320 -380 2340 -360
rect 2360 -380 2380 -360
rect 2400 -380 2420 -360
rect 2440 -380 2460 -360
rect 2480 -380 2500 -360
rect 2520 -380 2540 -360
rect 2560 -380 2580 -360
rect 2600 -380 2620 -360
rect 2640 -380 2660 -360
rect 2680 -380 2700 -360
rect 2720 -380 2740 -360
rect 2760 -380 2780 -360
rect 2800 -380 2820 -360
rect 2840 -380 2860 -360
rect 2880 -380 2900 -360
rect 2920 -380 2940 -360
rect 2960 -380 2980 -360
rect 3000 -380 3020 -360
rect 3040 -380 3060 -360
rect 3080 -380 3100 -360
rect 3120 -380 3140 -360
rect 3160 -380 3180 -360
rect 3200 -380 3220 -360
rect 3240 -380 3260 -360
rect 3280 -380 3300 -360
rect 3320 -380 3340 -360
rect 3360 -380 3380 -360
rect 3400 -380 3420 -360
rect 3440 -380 3460 -360
rect 3480 -380 3500 -360
rect 3520 -380 3540 -360
rect 3560 -380 3580 -360
rect 3600 -380 3615 -360
rect -3485 -390 3615 -380
rect 3635 -405 3790 -395
rect 3635 -435 3645 -405
rect 3665 -435 3685 -405
rect 3705 -435 3725 -405
rect 3745 -435 3765 -405
rect 3785 -435 3790 -405
rect 3635 -445 3790 -435
rect -3485 -460 3615 -450
rect -3485 -480 -3470 -460
rect -3450 -480 -3430 -460
rect -3410 -480 -3390 -460
rect -3370 -480 -3350 -460
rect -3330 -480 -3310 -460
rect -3290 -480 -3270 -460
rect -3250 -480 -3230 -460
rect -3210 -480 -3190 -460
rect -3170 -480 -3150 -460
rect -3130 -480 -3110 -460
rect -3090 -480 -3070 -460
rect -3050 -480 -3030 -460
rect -3010 -480 -2990 -460
rect -2970 -480 -2950 -460
rect -2930 -480 -2910 -460
rect -2890 -480 -2870 -460
rect -2850 -480 -2830 -460
rect -2810 -480 -2790 -460
rect -2770 -480 -2750 -460
rect -2730 -480 -2710 -460
rect -2690 -480 -2670 -460
rect -2650 -480 -2630 -460
rect -2610 -480 -2590 -460
rect -2570 -480 -2550 -460
rect -2530 -480 -2510 -460
rect -2490 -480 -2470 -460
rect -2450 -480 -2430 -460
rect -2410 -480 -2390 -460
rect -2370 -480 -2350 -460
rect -2330 -480 -2310 -460
rect -2290 -480 -2270 -460
rect -2250 -480 -2230 -460
rect -2210 -480 -2190 -460
rect -2170 -480 -2150 -460
rect -2130 -480 -2110 -460
rect -2090 -480 -2070 -460
rect -2050 -480 -2030 -460
rect -2010 -480 -1990 -460
rect -1970 -480 -1950 -460
rect -1930 -480 -1910 -460
rect -1890 -480 -1870 -460
rect -1850 -480 -1830 -460
rect -1810 -480 -1790 -460
rect -1770 -480 -1750 -460
rect -1730 -480 -1710 -460
rect -1690 -480 -1670 -460
rect -1650 -480 -1630 -460
rect -1610 -480 -1590 -460
rect -1570 -480 -1550 -460
rect -1530 -480 -1510 -460
rect -1460 -480 -1440 -460
rect -1420 -480 -1400 -460
rect -1380 -480 -1360 -460
rect -1340 -480 -1320 -460
rect -1300 -480 -1280 -460
rect -1260 -480 -1240 -460
rect -1220 -480 -1200 -460
rect -1180 -480 -1160 -460
rect -1140 -480 -1120 -460
rect -1100 -480 -1080 -460
rect -1060 -480 -1040 -460
rect -1020 -480 -1000 -460
rect -980 -480 -960 -460
rect -940 -480 -920 -460
rect -900 -480 -880 -460
rect -860 -480 -840 -460
rect -820 -480 -800 -460
rect -780 -480 -760 -460
rect -740 -480 -720 -460
rect -700 -480 -680 -460
rect -660 -480 -640 -460
rect -620 -480 -600 -460
rect -580 -480 -560 -460
rect -540 -480 -520 -460
rect -500 -480 -480 -460
rect -460 -480 -440 -460
rect -420 -480 -400 -460
rect -380 -480 -360 -460
rect -340 -480 -320 -460
rect -300 -480 -280 -460
rect -260 -480 -230 -460
rect -210 -480 -190 -460
rect -170 -480 -150 -460
rect -130 -480 -110 -460
rect -90 -480 -70 -460
rect -50 -480 -30 -460
rect -10 -480 10 -460
rect 30 -480 50 -460
rect 80 -480 100 -460
rect 120 -480 140 -460
rect 160 -480 180 -460
rect 200 -480 220 -460
rect 240 -480 260 -460
rect 280 -480 300 -460
rect 320 -480 340 -460
rect 360 -480 390 -460
rect 410 -480 430 -460
rect 450 -480 470 -460
rect 490 -480 510 -460
rect 530 -480 550 -460
rect 570 -480 590 -460
rect 610 -480 630 -460
rect 650 -480 670 -460
rect 690 -480 710 -460
rect 730 -480 750 -460
rect 770 -480 790 -460
rect 810 -480 830 -460
rect 850 -480 870 -460
rect 890 -480 910 -460
rect 930 -480 950 -460
rect 970 -480 990 -460
rect 1010 -480 1030 -460
rect 1050 -480 1070 -460
rect 1090 -480 1110 -460
rect 1130 -480 1150 -460
rect 1170 -480 1190 -460
rect 1210 -480 1230 -460
rect 1250 -480 1270 -460
rect 1290 -480 1310 -460
rect 1330 -480 1350 -460
rect 1370 -480 1390 -460
rect 1410 -480 1430 -460
rect 1450 -480 1470 -460
rect 1490 -480 1510 -460
rect 1530 -480 1550 -460
rect 1570 -480 1590 -460
rect 1640 -480 1660 -460
rect 1680 -480 1700 -460
rect 1720 -480 1740 -460
rect 1760 -480 1780 -460
rect 1800 -480 1820 -460
rect 1840 -480 1860 -460
rect 1880 -480 1900 -460
rect 1920 -480 1940 -460
rect 1960 -480 1980 -460
rect 2000 -480 2020 -460
rect 2040 -480 2060 -460
rect 2080 -480 2100 -460
rect 2120 -480 2140 -460
rect 2160 -480 2180 -460
rect 2200 -480 2220 -460
rect 2240 -480 2260 -460
rect 2280 -480 2300 -460
rect 2320 -480 2340 -460
rect 2360 -480 2380 -460
rect 2400 -480 2420 -460
rect 2440 -480 2460 -460
rect 2480 -480 2500 -460
rect 2520 -480 2540 -460
rect 2560 -480 2580 -460
rect 2600 -480 2620 -460
rect 2640 -480 2660 -460
rect 2680 -480 2700 -460
rect 2720 -480 2740 -460
rect 2760 -480 2780 -460
rect 2800 -480 2820 -460
rect 2840 -480 2860 -460
rect 2880 -480 2900 -460
rect 2920 -480 2940 -460
rect 2960 -480 2980 -460
rect 3000 -480 3020 -460
rect 3040 -480 3060 -460
rect 3080 -480 3100 -460
rect 3120 -480 3140 -460
rect 3160 -480 3180 -460
rect 3200 -480 3220 -460
rect 3240 -480 3260 -460
rect 3280 -480 3300 -460
rect 3320 -480 3340 -460
rect 3360 -480 3380 -460
rect 3400 -480 3420 -460
rect 3440 -480 3460 -460
rect 3480 -480 3500 -460
rect 3520 -480 3540 -460
rect 3560 -480 3580 -460
rect 3600 -480 3615 -460
rect -3485 -490 3615 -480
rect 3635 -505 3790 -495
rect 3635 -535 3645 -505
rect 3665 -535 3685 -505
rect 3705 -535 3725 -505
rect 3745 -535 3765 -505
rect 3785 -535 3790 -505
rect 3635 -545 3790 -535
rect -3485 -560 3615 -550
rect -3485 -580 -3470 -560
rect -3450 -580 -3430 -560
rect -3410 -580 -3390 -560
rect -3370 -580 -3350 -560
rect -3330 -580 -3310 -560
rect -3290 -580 -3270 -560
rect -3250 -580 -3230 -560
rect -3210 -580 -3190 -560
rect -3170 -580 -3150 -560
rect -3130 -580 -3110 -560
rect -3090 -580 -3070 -560
rect -3050 -580 -3030 -560
rect -3010 -580 -2990 -560
rect -2970 -580 -2950 -560
rect -2930 -580 -2910 -560
rect -2890 -580 -2870 -560
rect -2850 -580 -2830 -560
rect -2810 -580 -2790 -560
rect -2770 -580 -2750 -560
rect -2730 -580 -2710 -560
rect -2690 -580 -2670 -560
rect -2650 -580 -2630 -560
rect -2610 -580 -2590 -560
rect -2570 -580 -2550 -560
rect -2530 -580 -2510 -560
rect -2490 -580 -2470 -560
rect -2450 -580 -2430 -560
rect -2410 -580 -2390 -560
rect -2370 -580 -2350 -560
rect -2330 -580 -2310 -560
rect -2290 -580 -2270 -560
rect -2250 -580 -2230 -560
rect -2210 -580 -2190 -560
rect -2170 -580 -2150 -560
rect -2130 -580 -2110 -560
rect -2090 -580 -2070 -560
rect -2050 -580 -2030 -560
rect -2010 -580 -1990 -560
rect -1970 -580 -1950 -560
rect -1930 -580 -1910 -560
rect -1890 -580 -1870 -560
rect -1850 -580 -1830 -560
rect -1810 -580 -1790 -560
rect -1770 -580 -1750 -560
rect -1730 -580 -1710 -560
rect -1690 -580 -1670 -560
rect -1650 -580 -1630 -560
rect -1610 -580 -1590 -560
rect -1570 -580 -1550 -560
rect -1530 -580 -1510 -560
rect -1460 -580 -1440 -560
rect -1420 -580 -1400 -560
rect -1380 -580 -1360 -560
rect -1340 -580 -1320 -560
rect -1300 -580 -1280 -560
rect -1260 -580 -1240 -560
rect -1220 -580 -1200 -560
rect -1180 -580 -1160 -560
rect -1140 -580 -1120 -560
rect -1100 -580 -1080 -560
rect -1060 -580 -1040 -560
rect -1020 -580 -1000 -560
rect -980 -580 -960 -560
rect -940 -580 -920 -560
rect -900 -580 -880 -560
rect -860 -580 -840 -560
rect -820 -580 -800 -560
rect -780 -580 -760 -560
rect -740 -580 -720 -560
rect -700 -580 -680 -560
rect -660 -580 -640 -560
rect -620 -580 -600 -560
rect -580 -580 -560 -560
rect -540 -580 -520 -560
rect -500 -580 -480 -560
rect -460 -580 -440 -560
rect -420 -580 -400 -560
rect -380 -580 -360 -560
rect -340 -580 -320 -560
rect -300 -580 -280 -560
rect -260 -580 -230 -560
rect -210 -580 -190 -560
rect -170 -580 -150 -560
rect -130 -580 -110 -560
rect -90 -580 -70 -560
rect -50 -580 -30 -560
rect -10 -580 10 -560
rect 30 -580 50 -560
rect 80 -580 100 -560
rect 120 -580 140 -560
rect 160 -580 180 -560
rect 200 -580 220 -560
rect 240 -580 260 -560
rect 280 -580 300 -560
rect 320 -580 340 -560
rect 360 -580 390 -560
rect 410 -580 430 -560
rect 450 -580 470 -560
rect 490 -580 510 -560
rect 530 -580 550 -560
rect 570 -580 590 -560
rect 610 -580 630 -560
rect 650 -580 670 -560
rect 690 -580 710 -560
rect 730 -580 750 -560
rect 770 -580 790 -560
rect 810 -580 830 -560
rect 850 -580 870 -560
rect 890 -580 910 -560
rect 930 -580 950 -560
rect 970 -580 990 -560
rect 1010 -580 1030 -560
rect 1050 -580 1070 -560
rect 1090 -580 1110 -560
rect 1130 -580 1150 -560
rect 1170 -580 1190 -560
rect 1210 -580 1230 -560
rect 1250 -580 1270 -560
rect 1290 -580 1310 -560
rect 1330 -580 1350 -560
rect 1370 -580 1390 -560
rect 1410 -580 1430 -560
rect 1450 -580 1470 -560
rect 1490 -580 1510 -560
rect 1530 -580 1550 -560
rect 1570 -580 1590 -560
rect 1640 -580 1660 -560
rect 1680 -580 1700 -560
rect 1720 -580 1740 -560
rect 1760 -580 1780 -560
rect 1800 -580 1820 -560
rect 1840 -580 1860 -560
rect 1880 -580 1900 -560
rect 1920 -580 1940 -560
rect 1960 -580 1980 -560
rect 2000 -580 2020 -560
rect 2040 -580 2060 -560
rect 2080 -580 2100 -560
rect 2120 -580 2140 -560
rect 2160 -580 2180 -560
rect 2200 -580 2220 -560
rect 2240 -580 2260 -560
rect 2280 -580 2300 -560
rect 2320 -580 2340 -560
rect 2360 -580 2380 -560
rect 2400 -580 2420 -560
rect 2440 -580 2460 -560
rect 2480 -580 2500 -560
rect 2520 -580 2540 -560
rect 2560 -580 2580 -560
rect 2600 -580 2620 -560
rect 2640 -580 2660 -560
rect 2680 -580 2700 -560
rect 2720 -580 2740 -560
rect 2760 -580 2780 -560
rect 2800 -580 2820 -560
rect 2840 -580 2860 -560
rect 2880 -580 2900 -560
rect 2920 -580 2940 -560
rect 2960 -580 2980 -560
rect 3000 -580 3020 -560
rect 3040 -580 3060 -560
rect 3080 -580 3100 -560
rect 3120 -580 3140 -560
rect 3160 -580 3180 -560
rect 3200 -580 3220 -560
rect 3240 -580 3260 -560
rect 3280 -580 3300 -560
rect 3320 -580 3340 -560
rect 3360 -580 3380 -560
rect 3400 -580 3420 -560
rect 3440 -580 3460 -560
rect 3480 -580 3500 -560
rect 3520 -580 3540 -560
rect 3560 -580 3580 -560
rect 3600 -580 3615 -560
rect -3485 -590 3615 -580
rect 3635 -605 3790 -595
rect 3635 -635 3645 -605
rect 3665 -635 3685 -605
rect 3705 -635 3725 -605
rect 3745 -635 3765 -605
rect 3785 -635 3790 -605
rect 3635 -645 3790 -635
rect -3485 -660 3615 -650
rect -3485 -680 -3470 -660
rect -3450 -680 -3430 -660
rect -3410 -680 -3390 -660
rect -3370 -680 -3350 -660
rect -3330 -680 -3310 -660
rect -3290 -680 -3270 -660
rect -3250 -680 -3230 -660
rect -3210 -680 -3190 -660
rect -3170 -680 -3150 -660
rect -3130 -680 -3110 -660
rect -3090 -680 -3070 -660
rect -3050 -680 -3030 -660
rect -3010 -680 -2990 -660
rect -2970 -680 -2950 -660
rect -2930 -680 -2910 -660
rect -2890 -680 -2870 -660
rect -2850 -680 -2830 -660
rect -2810 -680 -2790 -660
rect -2770 -680 -2750 -660
rect -2730 -680 -2710 -660
rect -2690 -680 -2670 -660
rect -2650 -680 -2630 -660
rect -2610 -680 -2590 -660
rect -2570 -680 -2550 -660
rect -2530 -680 -2510 -660
rect -2490 -680 -2470 -660
rect -2450 -680 -2430 -660
rect -2410 -680 -2390 -660
rect -2370 -680 -2350 -660
rect -2330 -680 -2310 -660
rect -2290 -680 -2270 -660
rect -2250 -680 -2230 -660
rect -2210 -680 -2190 -660
rect -2170 -680 -2150 -660
rect -2130 -680 -2110 -660
rect -2090 -680 -2070 -660
rect -2050 -680 -2030 -660
rect -2010 -680 -1990 -660
rect -1970 -680 -1950 -660
rect -1930 -680 -1910 -660
rect -1890 -680 -1870 -660
rect -1850 -680 -1830 -660
rect -1810 -680 -1790 -660
rect -1770 -680 -1750 -660
rect -1730 -680 -1710 -660
rect -1690 -680 -1670 -660
rect -1650 -680 -1630 -660
rect -1610 -680 -1590 -660
rect -1570 -680 -1550 -660
rect -1530 -680 -1510 -660
rect -1460 -680 -1440 -660
rect -1420 -680 -1400 -660
rect -1380 -680 -1360 -660
rect -1340 -680 -1320 -660
rect -1300 -680 -1280 -660
rect -1260 -680 -1240 -660
rect -1220 -680 -1200 -660
rect -1180 -680 -1160 -660
rect -1140 -680 -1120 -660
rect -1100 -680 -1080 -660
rect -1060 -680 -1040 -660
rect -1020 -680 -1000 -660
rect -980 -680 -960 -660
rect -940 -680 -920 -660
rect -900 -680 -880 -660
rect -860 -680 -840 -660
rect -820 -680 -800 -660
rect -780 -680 -760 -660
rect -740 -680 -720 -660
rect -700 -680 -680 -660
rect -660 -680 -640 -660
rect -620 -680 -600 -660
rect -580 -680 -560 -660
rect -540 -680 -520 -660
rect -500 -680 -480 -660
rect -460 -680 -440 -660
rect -420 -680 -400 -660
rect -380 -680 -360 -660
rect -340 -680 -320 -660
rect -300 -680 -280 -660
rect -260 -680 -230 -660
rect -210 -680 -190 -660
rect -170 -680 -150 -660
rect -130 -680 -110 -660
rect -90 -680 -70 -660
rect -50 -680 -30 -660
rect -10 -680 10 -660
rect 30 -680 50 -660
rect 80 -680 100 -660
rect 120 -680 140 -660
rect 160 -680 180 -660
rect 200 -680 220 -660
rect 240 -680 260 -660
rect 280 -680 300 -660
rect 320 -680 340 -660
rect 360 -680 390 -660
rect 410 -680 430 -660
rect 450 -680 470 -660
rect 490 -680 510 -660
rect 530 -680 550 -660
rect 570 -680 590 -660
rect 610 -680 630 -660
rect 650 -680 670 -660
rect 690 -680 710 -660
rect 730 -680 750 -660
rect 770 -680 790 -660
rect 810 -680 830 -660
rect 850 -680 870 -660
rect 890 -680 910 -660
rect 930 -680 950 -660
rect 970 -680 990 -660
rect 1010 -680 1030 -660
rect 1050 -680 1070 -660
rect 1090 -680 1110 -660
rect 1130 -680 1150 -660
rect 1170 -680 1190 -660
rect 1210 -680 1230 -660
rect 1250 -680 1270 -660
rect 1290 -680 1310 -660
rect 1330 -680 1350 -660
rect 1370 -680 1390 -660
rect 1410 -680 1430 -660
rect 1450 -680 1470 -660
rect 1490 -680 1510 -660
rect 1530 -680 1550 -660
rect 1570 -680 1590 -660
rect 1640 -680 1660 -660
rect 1680 -680 1700 -660
rect 1720 -680 1740 -660
rect 1760 -680 1780 -660
rect 1800 -680 1820 -660
rect 1840 -680 1860 -660
rect 1880 -680 1900 -660
rect 1920 -680 1940 -660
rect 1960 -680 1980 -660
rect 2000 -680 2020 -660
rect 2040 -680 2060 -660
rect 2080 -680 2100 -660
rect 2120 -680 2140 -660
rect 2160 -680 2180 -660
rect 2200 -680 2220 -660
rect 2240 -680 2260 -660
rect 2280 -680 2300 -660
rect 2320 -680 2340 -660
rect 2360 -680 2380 -660
rect 2400 -680 2420 -660
rect 2440 -680 2460 -660
rect 2480 -680 2500 -660
rect 2520 -680 2540 -660
rect 2560 -680 2580 -660
rect 2600 -680 2620 -660
rect 2640 -680 2660 -660
rect 2680 -680 2700 -660
rect 2720 -680 2740 -660
rect 2760 -680 2780 -660
rect 2800 -680 2820 -660
rect 2840 -680 2860 -660
rect 2880 -680 2900 -660
rect 2920 -680 2940 -660
rect 2960 -680 2980 -660
rect 3000 -680 3020 -660
rect 3040 -680 3060 -660
rect 3080 -680 3100 -660
rect 3120 -680 3140 -660
rect 3160 -680 3180 -660
rect 3200 -680 3220 -660
rect 3240 -680 3260 -660
rect 3280 -680 3300 -660
rect 3320 -680 3340 -660
rect 3360 -680 3380 -660
rect 3400 -680 3420 -660
rect 3440 -680 3460 -660
rect 3480 -680 3500 -660
rect 3520 -680 3540 -660
rect 3560 -680 3580 -660
rect 3600 -680 3615 -660
rect -3485 -690 3615 -680
rect 3635 -705 3790 -695
rect 3635 -735 3645 -705
rect 3665 -735 3685 -705
rect 3705 -735 3725 -705
rect 3745 -735 3765 -705
rect 3785 -735 3790 -705
rect 3635 -745 3790 -735
rect -3485 -760 3615 -750
rect -3485 -780 -3470 -760
rect -3450 -780 -3430 -760
rect -3410 -780 -3390 -760
rect -3370 -780 -3350 -760
rect -3330 -780 -3310 -760
rect -3290 -780 -3270 -760
rect -3250 -780 -3230 -760
rect -3210 -780 -3190 -760
rect -3170 -780 -3150 -760
rect -3130 -780 -3110 -760
rect -3090 -780 -3070 -760
rect -3050 -780 -3030 -760
rect -3010 -780 -2990 -760
rect -2970 -780 -2950 -760
rect -2930 -780 -2910 -760
rect -2890 -780 -2870 -760
rect -2850 -780 -2830 -760
rect -2810 -780 -2790 -760
rect -2770 -780 -2750 -760
rect -2730 -780 -2710 -760
rect -2690 -780 -2670 -760
rect -2650 -780 -2630 -760
rect -2610 -780 -2590 -760
rect -2570 -780 -2550 -760
rect -2530 -780 -2510 -760
rect -2490 -780 -2470 -760
rect -2450 -780 -2430 -760
rect -2410 -780 -2390 -760
rect -2370 -780 -2350 -760
rect -2330 -780 -2310 -760
rect -2290 -780 -2270 -760
rect -2250 -780 -2230 -760
rect -2210 -780 -2190 -760
rect -2170 -780 -2150 -760
rect -2130 -780 -2110 -760
rect -2090 -780 -2070 -760
rect -2050 -780 -2030 -760
rect -2010 -780 -1990 -760
rect -1970 -780 -1950 -760
rect -1930 -780 -1910 -760
rect -1890 -780 -1870 -760
rect -1850 -780 -1830 -760
rect -1810 -780 -1790 -760
rect -1770 -780 -1750 -760
rect -1730 -780 -1710 -760
rect -1690 -780 -1670 -760
rect -1650 -780 -1630 -760
rect -1610 -780 -1590 -760
rect -1570 -780 -1550 -760
rect -1530 -780 -1510 -760
rect -1460 -780 -1440 -760
rect -1420 -780 -1400 -760
rect -1380 -780 -1360 -760
rect -1340 -780 -1320 -760
rect -1300 -780 -1280 -760
rect -1260 -780 -1240 -760
rect -1220 -780 -1200 -760
rect -1180 -780 -1160 -760
rect -1140 -780 -1120 -760
rect -1100 -780 -1080 -760
rect -1060 -780 -1040 -760
rect -1020 -780 -1000 -760
rect -980 -780 -960 -760
rect -940 -780 -920 -760
rect -900 -780 -880 -760
rect -860 -780 -840 -760
rect -820 -780 -800 -760
rect -780 -780 -760 -760
rect -740 -780 -720 -760
rect -700 -780 -680 -760
rect -660 -780 -640 -760
rect -620 -780 -600 -760
rect -580 -780 -560 -760
rect -540 -780 -520 -760
rect -500 -780 -480 -760
rect -460 -780 -440 -760
rect -420 -780 -400 -760
rect -380 -780 -360 -760
rect -340 -780 -320 -760
rect -300 -780 -280 -760
rect -260 -780 -230 -760
rect -210 -780 -190 -760
rect -170 -780 -150 -760
rect -130 -780 -110 -760
rect -90 -780 -70 -760
rect -50 -780 -30 -760
rect -10 -780 10 -760
rect 30 -780 50 -760
rect 80 -780 100 -760
rect 120 -780 140 -760
rect 160 -780 180 -760
rect 200 -780 220 -760
rect 240 -780 260 -760
rect 280 -780 300 -760
rect 320 -780 340 -760
rect 360 -780 390 -760
rect 410 -780 430 -760
rect 450 -780 470 -760
rect 490 -780 510 -760
rect 530 -780 550 -760
rect 570 -780 590 -760
rect 610 -780 630 -760
rect 650 -780 670 -760
rect 690 -780 710 -760
rect 730 -780 750 -760
rect 770 -780 790 -760
rect 810 -780 830 -760
rect 850 -780 870 -760
rect 890 -780 910 -760
rect 930 -780 950 -760
rect 970 -780 990 -760
rect 1010 -780 1030 -760
rect 1050 -780 1070 -760
rect 1090 -780 1110 -760
rect 1130 -780 1150 -760
rect 1170 -780 1190 -760
rect 1210 -780 1230 -760
rect 1250 -780 1270 -760
rect 1290 -780 1310 -760
rect 1330 -780 1350 -760
rect 1370 -780 1390 -760
rect 1410 -780 1430 -760
rect 1450 -780 1470 -760
rect 1490 -780 1510 -760
rect 1530 -780 1550 -760
rect 1570 -780 1590 -760
rect 1640 -780 1660 -760
rect 1680 -780 1700 -760
rect 1720 -780 1740 -760
rect 1760 -780 1780 -760
rect 1800 -780 1820 -760
rect 1840 -780 1860 -760
rect 1880 -780 1900 -760
rect 1920 -780 1940 -760
rect 1960 -780 1980 -760
rect 2000 -780 2020 -760
rect 2040 -780 2060 -760
rect 2080 -780 2100 -760
rect 2120 -780 2140 -760
rect 2160 -780 2180 -760
rect 2200 -780 2220 -760
rect 2240 -780 2260 -760
rect 2280 -780 2300 -760
rect 2320 -780 2340 -760
rect 2360 -780 2380 -760
rect 2400 -780 2420 -760
rect 2440 -780 2460 -760
rect 2480 -780 2500 -760
rect 2520 -780 2540 -760
rect 2560 -780 2580 -760
rect 2600 -780 2620 -760
rect 2640 -780 2660 -760
rect 2680 -780 2700 -760
rect 2720 -780 2740 -760
rect 2760 -780 2780 -760
rect 2800 -780 2820 -760
rect 2840 -780 2860 -760
rect 2880 -780 2900 -760
rect 2920 -780 2940 -760
rect 2960 -780 2980 -760
rect 3000 -780 3020 -760
rect 3040 -780 3060 -760
rect 3080 -780 3100 -760
rect 3120 -780 3140 -760
rect 3160 -780 3180 -760
rect 3200 -780 3220 -760
rect 3240 -780 3260 -760
rect 3280 -780 3300 -760
rect 3320 -780 3340 -760
rect 3360 -780 3380 -760
rect 3400 -780 3420 -760
rect 3440 -780 3460 -760
rect 3480 -780 3500 -760
rect 3520 -780 3540 -760
rect 3560 -780 3580 -760
rect 3600 -780 3615 -760
rect -3485 -790 3615 -780
rect 3635 -805 3790 -795
rect 3635 -835 3645 -805
rect 3665 -835 3685 -805
rect 3705 -835 3725 -805
rect 3745 -835 3765 -805
rect 3785 -835 3790 -805
rect 3635 -845 3790 -835
rect -3485 -860 3615 -850
rect -3485 -880 -3470 -860
rect -3450 -880 -3430 -860
rect -3410 -880 -3390 -860
rect -3370 -880 -3350 -860
rect -3330 -880 -3310 -860
rect -3290 -880 -3270 -860
rect -3250 -880 -3230 -860
rect -3210 -880 -3190 -860
rect -3170 -880 -3150 -860
rect -3130 -880 -3110 -860
rect -3090 -880 -3070 -860
rect -3050 -880 -3030 -860
rect -3010 -880 -2990 -860
rect -2970 -880 -2950 -860
rect -2930 -880 -2910 -860
rect -2890 -880 -2870 -860
rect -2850 -880 -2830 -860
rect -2810 -880 -2790 -860
rect -2770 -880 -2750 -860
rect -2730 -880 -2710 -860
rect -2690 -880 -2670 -860
rect -2650 -880 -2630 -860
rect -2610 -880 -2590 -860
rect -2570 -880 -2550 -860
rect -2530 -880 -2510 -860
rect -2490 -880 -2470 -860
rect -2450 -880 -2430 -860
rect -2410 -880 -2390 -860
rect -2370 -880 -2350 -860
rect -2330 -880 -2310 -860
rect -2290 -880 -2270 -860
rect -2250 -880 -2230 -860
rect -2210 -880 -2190 -860
rect -2170 -880 -2150 -860
rect -2130 -880 -2110 -860
rect -2090 -880 -2070 -860
rect -2050 -880 -2030 -860
rect -2010 -880 -1990 -860
rect -1970 -880 -1950 -860
rect -1930 -880 -1910 -860
rect -1890 -880 -1870 -860
rect -1850 -880 -1830 -860
rect -1810 -880 -1790 -860
rect -1770 -880 -1750 -860
rect -1730 -880 -1710 -860
rect -1690 -880 -1670 -860
rect -1650 -880 -1630 -860
rect -1610 -880 -1590 -860
rect -1570 -880 -1550 -860
rect -1530 -880 -1510 -860
rect -1460 -880 -1440 -860
rect -1420 -880 -1400 -860
rect -1380 -880 -1360 -860
rect -1340 -880 -1320 -860
rect -1300 -880 -1280 -860
rect -1260 -880 -1240 -860
rect -1220 -880 -1200 -860
rect -1180 -880 -1160 -860
rect -1140 -880 -1120 -860
rect -1100 -880 -1080 -860
rect -1060 -880 -1040 -860
rect -1020 -880 -1000 -860
rect -980 -880 -960 -860
rect -940 -880 -920 -860
rect -900 -880 -880 -860
rect -860 -880 -840 -860
rect -820 -880 -800 -860
rect -780 -880 -760 -860
rect -740 -880 -720 -860
rect -700 -880 -680 -860
rect -660 -880 -640 -860
rect -620 -880 -600 -860
rect -580 -880 -560 -860
rect -540 -880 -520 -860
rect -500 -880 -480 -860
rect -460 -880 -440 -860
rect -420 -880 -400 -860
rect -380 -880 -360 -860
rect -340 -880 -320 -860
rect -300 -880 -280 -860
rect -260 -880 -230 -860
rect -210 -880 -190 -860
rect -170 -880 -150 -860
rect -130 -880 -110 -860
rect -90 -880 -70 -860
rect -50 -880 -30 -860
rect -10 -880 10 -860
rect 30 -880 50 -860
rect 80 -880 100 -860
rect 120 -880 140 -860
rect 160 -880 180 -860
rect 200 -880 220 -860
rect 240 -880 260 -860
rect 280 -880 300 -860
rect 320 -880 340 -860
rect 360 -880 390 -860
rect 410 -880 430 -860
rect 450 -880 470 -860
rect 490 -880 510 -860
rect 530 -880 550 -860
rect 570 -880 590 -860
rect 610 -880 630 -860
rect 650 -880 670 -860
rect 690 -880 710 -860
rect 730 -880 750 -860
rect 770 -880 790 -860
rect 810 -880 830 -860
rect 850 -880 870 -860
rect 890 -880 910 -860
rect 930 -880 950 -860
rect 970 -880 990 -860
rect 1010 -880 1030 -860
rect 1050 -880 1070 -860
rect 1090 -880 1110 -860
rect 1130 -880 1150 -860
rect 1170 -880 1190 -860
rect 1210 -880 1230 -860
rect 1250 -880 1270 -860
rect 1290 -880 1310 -860
rect 1330 -880 1350 -860
rect 1370 -880 1390 -860
rect 1410 -880 1430 -860
rect 1450 -880 1470 -860
rect 1490 -880 1510 -860
rect 1530 -880 1550 -860
rect 1570 -880 1590 -860
rect 1640 -880 1660 -860
rect 1680 -880 1700 -860
rect 1720 -880 1740 -860
rect 1760 -880 1780 -860
rect 1800 -880 1820 -860
rect 1840 -880 1860 -860
rect 1880 -880 1900 -860
rect 1920 -880 1940 -860
rect 1960 -880 1980 -860
rect 2000 -880 2020 -860
rect 2040 -880 2060 -860
rect 2080 -880 2100 -860
rect 2120 -880 2140 -860
rect 2160 -880 2180 -860
rect 2200 -880 2220 -860
rect 2240 -880 2260 -860
rect 2280 -880 2300 -860
rect 2320 -880 2340 -860
rect 2360 -880 2380 -860
rect 2400 -880 2420 -860
rect 2440 -880 2460 -860
rect 2480 -880 2500 -860
rect 2520 -880 2540 -860
rect 2560 -880 2580 -860
rect 2600 -880 2620 -860
rect 2640 -880 2660 -860
rect 2680 -880 2700 -860
rect 2720 -880 2740 -860
rect 2760 -880 2780 -860
rect 2800 -880 2820 -860
rect 2840 -880 2860 -860
rect 2880 -880 2900 -860
rect 2920 -880 2940 -860
rect 2960 -880 2980 -860
rect 3000 -880 3020 -860
rect 3040 -880 3060 -860
rect 3080 -880 3100 -860
rect 3120 -880 3140 -860
rect 3160 -880 3180 -860
rect 3200 -880 3220 -860
rect 3240 -880 3260 -860
rect 3280 -880 3300 -860
rect 3320 -880 3340 -860
rect 3360 -880 3380 -860
rect 3400 -880 3420 -860
rect 3440 -880 3460 -860
rect 3480 -880 3500 -860
rect 3520 -880 3540 -860
rect 3560 -880 3580 -860
rect 3600 -880 3615 -860
rect -3485 -890 3615 -880
rect 3635 -905 3790 -895
rect 3635 -935 3645 -905
rect 3665 -935 3685 -905
rect 3705 -935 3725 -905
rect 3745 -935 3765 -905
rect 3785 -935 3790 -905
rect 3635 -945 3790 -935
rect -3485 -960 3615 -950
rect -3485 -980 -3470 -960
rect -3450 -980 -3430 -960
rect -3410 -980 -3390 -960
rect -3370 -980 -3350 -960
rect -3330 -980 -3310 -960
rect -3290 -980 -3270 -960
rect -3250 -980 -3230 -960
rect -3210 -980 -3190 -960
rect -3170 -980 -3150 -960
rect -3130 -980 -3110 -960
rect -3090 -980 -3070 -960
rect -3050 -980 -3030 -960
rect -3010 -980 -2990 -960
rect -2970 -980 -2950 -960
rect -2930 -980 -2910 -960
rect -2890 -980 -2870 -960
rect -2850 -980 -2830 -960
rect -2810 -980 -2790 -960
rect -2770 -980 -2750 -960
rect -2730 -980 -2710 -960
rect -2690 -980 -2670 -960
rect -2650 -980 -2630 -960
rect -2610 -980 -2590 -960
rect -2570 -980 -2550 -960
rect -2530 -980 -2510 -960
rect -2490 -980 -2470 -960
rect -2450 -980 -2430 -960
rect -2410 -980 -2390 -960
rect -2370 -980 -2350 -960
rect -2330 -980 -2310 -960
rect -2290 -980 -2270 -960
rect -2250 -980 -2230 -960
rect -2210 -980 -2190 -960
rect -2170 -980 -2150 -960
rect -2130 -980 -2110 -960
rect -2090 -980 -2070 -960
rect -2050 -980 -2030 -960
rect -2010 -980 -1990 -960
rect -1970 -980 -1950 -960
rect -1930 -980 -1910 -960
rect -1890 -980 -1870 -960
rect -1850 -980 -1830 -960
rect -1810 -980 -1790 -960
rect -1770 -980 -1750 -960
rect -1730 -980 -1710 -960
rect -1690 -980 -1670 -960
rect -1650 -980 -1630 -960
rect -1610 -980 -1590 -960
rect -1570 -980 -1550 -960
rect -1530 -980 -1510 -960
rect -1460 -980 -1440 -960
rect -1420 -980 -1400 -960
rect -1380 -980 -1360 -960
rect -1340 -980 -1320 -960
rect -1300 -980 -1280 -960
rect -1260 -980 -1240 -960
rect -1220 -980 -1200 -960
rect -1180 -980 -1160 -960
rect -1140 -980 -1120 -960
rect -1100 -980 -1080 -960
rect -1060 -980 -1040 -960
rect -1020 -980 -1000 -960
rect -980 -980 -960 -960
rect -940 -980 -920 -960
rect -900 -980 -880 -960
rect -860 -980 -840 -960
rect -820 -980 -800 -960
rect -780 -980 -760 -960
rect -740 -980 -720 -960
rect -700 -980 -680 -960
rect -660 -980 -640 -960
rect -620 -980 -600 -960
rect -580 -980 -560 -960
rect -540 -980 -520 -960
rect -500 -980 -480 -960
rect -460 -980 -440 -960
rect -420 -980 -400 -960
rect -380 -980 -360 -960
rect -340 -980 -320 -960
rect -300 -980 -280 -960
rect -260 -980 -230 -960
rect -210 -980 -190 -960
rect -170 -980 -150 -960
rect -130 -980 -110 -960
rect -90 -980 -70 -960
rect -50 -980 -30 -960
rect -10 -980 10 -960
rect 30 -980 50 -960
rect 80 -980 100 -960
rect 120 -980 140 -960
rect 160 -980 180 -960
rect 200 -980 220 -960
rect 240 -980 260 -960
rect 280 -980 300 -960
rect 320 -980 340 -960
rect 360 -980 390 -960
rect 410 -980 430 -960
rect 450 -980 470 -960
rect 490 -980 510 -960
rect 530 -980 550 -960
rect 570 -980 590 -960
rect 610 -980 630 -960
rect 650 -980 670 -960
rect 690 -980 710 -960
rect 730 -980 750 -960
rect 770 -980 790 -960
rect 810 -980 830 -960
rect 850 -980 870 -960
rect 890 -980 910 -960
rect 930 -980 950 -960
rect 970 -980 990 -960
rect 1010 -980 1030 -960
rect 1050 -980 1070 -960
rect 1090 -980 1110 -960
rect 1130 -980 1150 -960
rect 1170 -980 1190 -960
rect 1210 -980 1230 -960
rect 1250 -980 1270 -960
rect 1290 -980 1310 -960
rect 1330 -980 1350 -960
rect 1370 -980 1390 -960
rect 1410 -980 1430 -960
rect 1450 -980 1470 -960
rect 1490 -980 1510 -960
rect 1530 -980 1550 -960
rect 1570 -980 1590 -960
rect 1640 -980 1660 -960
rect 1680 -980 1700 -960
rect 1720 -980 1740 -960
rect 1760 -980 1780 -960
rect 1800 -980 1820 -960
rect 1840 -980 1860 -960
rect 1880 -980 1900 -960
rect 1920 -980 1940 -960
rect 1960 -980 1980 -960
rect 2000 -980 2020 -960
rect 2040 -980 2060 -960
rect 2080 -980 2100 -960
rect 2120 -980 2140 -960
rect 2160 -980 2180 -960
rect 2200 -980 2220 -960
rect 2240 -980 2260 -960
rect 2280 -980 2300 -960
rect 2320 -980 2340 -960
rect 2360 -980 2380 -960
rect 2400 -980 2420 -960
rect 2440 -980 2460 -960
rect 2480 -980 2500 -960
rect 2520 -980 2540 -960
rect 2560 -980 2580 -960
rect 2600 -980 2620 -960
rect 2640 -980 2660 -960
rect 2680 -980 2700 -960
rect 2720 -980 2740 -960
rect 2760 -980 2780 -960
rect 2800 -980 2820 -960
rect 2840 -980 2860 -960
rect 2880 -980 2900 -960
rect 2920 -980 2940 -960
rect 2960 -980 2980 -960
rect 3000 -980 3020 -960
rect 3040 -980 3060 -960
rect 3080 -980 3100 -960
rect 3120 -980 3140 -960
rect 3160 -980 3180 -960
rect 3200 -980 3220 -960
rect 3240 -980 3260 -960
rect 3280 -980 3300 -960
rect 3320 -980 3340 -960
rect 3360 -980 3380 -960
rect 3400 -980 3420 -960
rect 3440 -980 3460 -960
rect 3480 -980 3500 -960
rect 3520 -980 3540 -960
rect 3560 -980 3580 -960
rect 3600 -980 3615 -960
rect -3485 -990 3615 -980
rect 3635 -1005 3790 -995
rect 3635 -1035 3645 -1005
rect 3665 -1035 3685 -1005
rect 3705 -1035 3725 -1005
rect 3745 -1035 3765 -1005
rect 3785 -1035 3790 -1005
rect 3635 -1045 3790 -1035
rect -3485 -1060 3615 -1050
rect -3485 -1080 -3470 -1060
rect -3450 -1080 -3430 -1060
rect -3410 -1080 -3390 -1060
rect -3370 -1080 -3350 -1060
rect -3330 -1080 -3310 -1060
rect -3290 -1080 -3270 -1060
rect -3250 -1080 -3230 -1060
rect -3210 -1080 -3190 -1060
rect -3170 -1080 -3150 -1060
rect -3130 -1080 -3110 -1060
rect -3090 -1080 -3070 -1060
rect -3050 -1080 -3030 -1060
rect -3010 -1080 -2990 -1060
rect -2970 -1080 -2950 -1060
rect -2930 -1080 -2910 -1060
rect -2890 -1080 -2870 -1060
rect -2850 -1080 -2830 -1060
rect -2810 -1080 -2790 -1060
rect -2770 -1080 -2750 -1060
rect -2730 -1080 -2710 -1060
rect -2690 -1080 -2670 -1060
rect -2650 -1080 -2630 -1060
rect -2610 -1080 -2590 -1060
rect -2570 -1080 -2550 -1060
rect -2530 -1080 -2510 -1060
rect -2490 -1080 -2470 -1060
rect -2450 -1080 -2430 -1060
rect -2410 -1080 -2390 -1060
rect -2370 -1080 -2350 -1060
rect -2330 -1080 -2310 -1060
rect -2290 -1080 -2270 -1060
rect -2250 -1080 -2230 -1060
rect -2210 -1080 -2190 -1060
rect -2170 -1080 -2150 -1060
rect -2130 -1080 -2110 -1060
rect -2090 -1080 -2070 -1060
rect -2050 -1080 -2030 -1060
rect -2010 -1080 -1990 -1060
rect -1970 -1080 -1950 -1060
rect -1930 -1080 -1910 -1060
rect -1890 -1080 -1870 -1060
rect -1850 -1080 -1830 -1060
rect -1810 -1080 -1790 -1060
rect -1770 -1080 -1750 -1060
rect -1730 -1080 -1710 -1060
rect -1690 -1080 -1670 -1060
rect -1650 -1080 -1630 -1060
rect -1610 -1080 -1590 -1060
rect -1570 -1080 -1550 -1060
rect -1530 -1080 -1510 -1060
rect -1460 -1080 -1440 -1060
rect -1420 -1080 -1400 -1060
rect -1380 -1080 -1360 -1060
rect -1340 -1080 -1320 -1060
rect -1300 -1080 -1280 -1060
rect -1260 -1080 -1240 -1060
rect -1220 -1080 -1200 -1060
rect -1180 -1080 -1160 -1060
rect -1140 -1080 -1120 -1060
rect -1100 -1080 -1080 -1060
rect -1060 -1080 -1040 -1060
rect -1020 -1080 -1000 -1060
rect -980 -1080 -960 -1060
rect -940 -1080 -920 -1060
rect -900 -1080 -880 -1060
rect -860 -1080 -840 -1060
rect -820 -1080 -800 -1060
rect -780 -1080 -760 -1060
rect -740 -1080 -720 -1060
rect -700 -1080 -680 -1060
rect -660 -1080 -640 -1060
rect -620 -1080 -600 -1060
rect -580 -1080 -560 -1060
rect -540 -1080 -520 -1060
rect -500 -1080 -480 -1060
rect -460 -1080 -440 -1060
rect -420 -1080 -400 -1060
rect -380 -1080 -360 -1060
rect -340 -1080 -320 -1060
rect -300 -1080 -280 -1060
rect -260 -1080 -230 -1060
rect -210 -1080 -190 -1060
rect -170 -1080 -150 -1060
rect -130 -1080 -110 -1060
rect -90 -1080 -70 -1060
rect -50 -1080 -30 -1060
rect -10 -1080 10 -1060
rect 30 -1080 50 -1060
rect 80 -1080 100 -1060
rect 120 -1080 140 -1060
rect 160 -1080 180 -1060
rect 200 -1080 220 -1060
rect 240 -1080 260 -1060
rect 280 -1080 300 -1060
rect 320 -1080 340 -1060
rect 360 -1080 390 -1060
rect 410 -1080 430 -1060
rect 450 -1080 470 -1060
rect 490 -1080 510 -1060
rect 530 -1080 550 -1060
rect 570 -1080 590 -1060
rect 610 -1080 630 -1060
rect 650 -1080 670 -1060
rect 690 -1080 710 -1060
rect 730 -1080 750 -1060
rect 770 -1080 790 -1060
rect 810 -1080 830 -1060
rect 850 -1080 870 -1060
rect 890 -1080 910 -1060
rect 930 -1080 950 -1060
rect 970 -1080 990 -1060
rect 1010 -1080 1030 -1060
rect 1050 -1080 1070 -1060
rect 1090 -1080 1110 -1060
rect 1130 -1080 1150 -1060
rect 1170 -1080 1190 -1060
rect 1210 -1080 1230 -1060
rect 1250 -1080 1270 -1060
rect 1290 -1080 1310 -1060
rect 1330 -1080 1350 -1060
rect 1370 -1080 1390 -1060
rect 1410 -1080 1430 -1060
rect 1450 -1080 1470 -1060
rect 1490 -1080 1510 -1060
rect 1530 -1080 1550 -1060
rect 1570 -1080 1590 -1060
rect 1640 -1080 1660 -1060
rect 1680 -1080 1700 -1060
rect 1720 -1080 1740 -1060
rect 1760 -1080 1780 -1060
rect 1800 -1080 1820 -1060
rect 1840 -1080 1860 -1060
rect 1880 -1080 1900 -1060
rect 1920 -1080 1940 -1060
rect 1960 -1080 1980 -1060
rect 2000 -1080 2020 -1060
rect 2040 -1080 2060 -1060
rect 2080 -1080 2100 -1060
rect 2120 -1080 2140 -1060
rect 2160 -1080 2180 -1060
rect 2200 -1080 2220 -1060
rect 2240 -1080 2260 -1060
rect 2280 -1080 2300 -1060
rect 2320 -1080 2340 -1060
rect 2360 -1080 2380 -1060
rect 2400 -1080 2420 -1060
rect 2440 -1080 2460 -1060
rect 2480 -1080 2500 -1060
rect 2520 -1080 2540 -1060
rect 2560 -1080 2580 -1060
rect 2600 -1080 2620 -1060
rect 2640 -1080 2660 -1060
rect 2680 -1080 2700 -1060
rect 2720 -1080 2740 -1060
rect 2760 -1080 2780 -1060
rect 2800 -1080 2820 -1060
rect 2840 -1080 2860 -1060
rect 2880 -1080 2900 -1060
rect 2920 -1080 2940 -1060
rect 2960 -1080 2980 -1060
rect 3000 -1080 3020 -1060
rect 3040 -1080 3060 -1060
rect 3080 -1080 3100 -1060
rect 3120 -1080 3140 -1060
rect 3160 -1080 3180 -1060
rect 3200 -1080 3220 -1060
rect 3240 -1080 3260 -1060
rect 3280 -1080 3300 -1060
rect 3320 -1080 3340 -1060
rect 3360 -1080 3380 -1060
rect 3400 -1080 3420 -1060
rect 3440 -1080 3460 -1060
rect 3480 -1080 3500 -1060
rect 3520 -1080 3540 -1060
rect 3560 -1080 3580 -1060
rect 3600 -1080 3615 -1060
rect -3485 -1090 3615 -1080
rect 3635 -1105 3790 -1095
rect 3635 -1135 3645 -1105
rect 3665 -1135 3685 -1105
rect 3705 -1135 3725 -1105
rect 3745 -1135 3765 -1105
rect 3785 -1135 3790 -1105
rect 3635 -1145 3790 -1135
rect -3485 -1160 3615 -1150
rect -3485 -1180 -3470 -1160
rect -3450 -1180 -3430 -1160
rect -3410 -1180 -3390 -1160
rect -3370 -1180 -3350 -1160
rect -3330 -1180 -3310 -1160
rect -3290 -1180 -3270 -1160
rect -3250 -1180 -3230 -1160
rect -3210 -1180 -3190 -1160
rect -3170 -1180 -3150 -1160
rect -3130 -1180 -3110 -1160
rect -3090 -1180 -3070 -1160
rect -3050 -1180 -3030 -1160
rect -3010 -1180 -2990 -1160
rect -2970 -1180 -2950 -1160
rect -2930 -1180 -2910 -1160
rect -2890 -1180 -2870 -1160
rect -2850 -1180 -2830 -1160
rect -2810 -1180 -2790 -1160
rect -2770 -1180 -2750 -1160
rect -2730 -1180 -2710 -1160
rect -2690 -1180 -2670 -1160
rect -2650 -1180 -2630 -1160
rect -2610 -1180 -2590 -1160
rect -2570 -1180 -2550 -1160
rect -2530 -1180 -2510 -1160
rect -2490 -1180 -2470 -1160
rect -2450 -1180 -2430 -1160
rect -2410 -1180 -2390 -1160
rect -2370 -1180 -2350 -1160
rect -2330 -1180 -2310 -1160
rect -2290 -1180 -2270 -1160
rect -2250 -1180 -2230 -1160
rect -2210 -1180 -2190 -1160
rect -2170 -1180 -2150 -1160
rect -2130 -1180 -2110 -1160
rect -2090 -1180 -2070 -1160
rect -2050 -1180 -2030 -1160
rect -2010 -1180 -1990 -1160
rect -1970 -1180 -1950 -1160
rect -1930 -1180 -1910 -1160
rect -1890 -1180 -1870 -1160
rect -1850 -1180 -1830 -1160
rect -1810 -1180 -1790 -1160
rect -1770 -1180 -1750 -1160
rect -1730 -1180 -1710 -1160
rect -1690 -1180 -1670 -1160
rect -1650 -1180 -1630 -1160
rect -1610 -1180 -1590 -1160
rect -1570 -1180 -1550 -1160
rect -1530 -1180 -1510 -1160
rect -1490 -1180 -1470 -1160
rect -1450 -1180 -1430 -1160
rect -1410 -1180 -1390 -1160
rect -1370 -1180 -1350 -1160
rect -1330 -1180 -1310 -1160
rect -1290 -1180 -1270 -1160
rect -1250 -1180 -1230 -1160
rect -1210 -1180 -1190 -1160
rect -1170 -1180 -1150 -1160
rect -1130 -1180 -1110 -1160
rect -1090 -1180 -1070 -1160
rect -1050 -1180 -1030 -1160
rect -1010 -1180 -990 -1160
rect -970 -1180 -950 -1160
rect -930 -1180 -910 -1160
rect -890 -1180 -870 -1160
rect -850 -1180 -830 -1160
rect -810 -1180 -790 -1160
rect -770 -1180 -750 -1160
rect -730 -1180 -710 -1160
rect -690 -1180 -670 -1160
rect -650 -1180 -630 -1160
rect -610 -1180 -590 -1160
rect -570 -1180 -550 -1160
rect -530 -1180 -510 -1160
rect -490 -1180 -470 -1160
rect -450 -1180 -430 -1160
rect -410 -1180 -390 -1160
rect -370 -1180 -350 -1160
rect -330 -1180 -310 -1160
rect -290 -1180 -270 -1160
rect -250 -1180 -230 -1160
rect -210 -1180 -190 -1160
rect -170 -1180 -150 -1160
rect -130 -1180 -110 -1160
rect -90 -1180 -70 -1160
rect -50 -1180 -30 -1160
rect -10 -1180 10 -1160
rect 30 -1180 50 -1160
rect 80 -1180 100 -1160
rect 120 -1180 140 -1160
rect 160 -1180 180 -1160
rect 200 -1180 220 -1160
rect 240 -1180 260 -1160
rect 280 -1180 300 -1160
rect 320 -1180 340 -1160
rect 360 -1180 380 -1160
rect 400 -1180 420 -1160
rect 440 -1180 460 -1160
rect 480 -1180 500 -1160
rect 520 -1180 540 -1160
rect 560 -1180 580 -1160
rect 600 -1180 620 -1160
rect 640 -1180 660 -1160
rect 680 -1180 700 -1160
rect 720 -1180 740 -1160
rect 760 -1180 780 -1160
rect 800 -1180 820 -1160
rect 840 -1180 860 -1160
rect 880 -1180 900 -1160
rect 920 -1180 940 -1160
rect 960 -1180 980 -1160
rect 1000 -1180 1020 -1160
rect 1040 -1180 1060 -1160
rect 1080 -1180 1100 -1160
rect 1120 -1180 1140 -1160
rect 1160 -1180 1180 -1160
rect 1200 -1180 1220 -1160
rect 1240 -1180 1260 -1160
rect 1280 -1180 1300 -1160
rect 1320 -1180 1340 -1160
rect 1360 -1180 1380 -1160
rect 1400 -1180 1420 -1160
rect 1440 -1180 1460 -1160
rect 1480 -1180 1500 -1160
rect 1520 -1180 1540 -1160
rect 1560 -1180 1580 -1160
rect 1600 -1180 1620 -1160
rect 1640 -1180 1660 -1160
rect 1680 -1180 1700 -1160
rect 1720 -1180 1740 -1160
rect 1760 -1180 1780 -1160
rect 1800 -1180 1820 -1160
rect 1840 -1180 1860 -1160
rect 1880 -1180 1900 -1160
rect 1920 -1180 1940 -1160
rect 1960 -1180 1980 -1160
rect 2000 -1180 2020 -1160
rect 2040 -1180 2060 -1160
rect 2080 -1180 2100 -1160
rect 2120 -1180 2140 -1160
rect 2160 -1180 2180 -1160
rect 2200 -1180 2220 -1160
rect 2240 -1180 2260 -1160
rect 2280 -1180 2300 -1160
rect 2320 -1180 2340 -1160
rect 2360 -1180 2380 -1160
rect 2400 -1180 2420 -1160
rect 2440 -1180 2460 -1160
rect 2480 -1180 2500 -1160
rect 2520 -1180 2540 -1160
rect 2560 -1180 2580 -1160
rect 2600 -1180 2620 -1160
rect 2640 -1180 2660 -1160
rect 2680 -1180 2700 -1160
rect 2720 -1180 2740 -1160
rect 2760 -1180 2780 -1160
rect 2800 -1180 2820 -1160
rect 2840 -1180 2860 -1160
rect 2880 -1180 2900 -1160
rect 2920 -1180 2940 -1160
rect 2960 -1180 2980 -1160
rect 3000 -1180 3020 -1160
rect 3040 -1180 3060 -1160
rect 3080 -1180 3100 -1160
rect 3120 -1180 3140 -1160
rect 3160 -1180 3180 -1160
rect 3200 -1180 3220 -1160
rect 3240 -1180 3260 -1160
rect 3280 -1180 3300 -1160
rect 3320 -1180 3340 -1160
rect 3360 -1180 3380 -1160
rect 3400 -1180 3420 -1160
rect 3440 -1180 3460 -1160
rect 3480 -1180 3500 -1160
rect 3520 -1180 3540 -1160
rect 3560 -1180 3580 -1160
rect 3600 -1180 3615 -1160
rect -3485 -1200 3615 -1180
rect -3485 -1220 -3470 -1200
rect -3450 -1220 -3430 -1200
rect -3410 -1220 -3390 -1200
rect -3370 -1220 -3350 -1200
rect -3330 -1220 -3310 -1200
rect -3290 -1220 -3270 -1200
rect -3250 -1220 -3230 -1200
rect -3210 -1220 -3190 -1200
rect -3170 -1220 -3150 -1200
rect -3130 -1220 -3110 -1200
rect -3090 -1220 -3070 -1200
rect -3050 -1220 -3030 -1200
rect -3010 -1220 -2990 -1200
rect -2970 -1220 -2950 -1200
rect -2930 -1220 -2910 -1200
rect -2890 -1220 -2870 -1200
rect -2850 -1220 -2830 -1200
rect -2810 -1220 -2790 -1200
rect -2770 -1220 -2750 -1200
rect -2730 -1220 -2710 -1200
rect -2690 -1220 -2670 -1200
rect -2650 -1220 -2630 -1200
rect -2610 -1220 -2590 -1200
rect -2570 -1220 -2550 -1200
rect -2530 -1220 -2510 -1200
rect -2490 -1220 -2470 -1200
rect -2450 -1220 -2430 -1200
rect -2410 -1220 -2390 -1200
rect -2370 -1220 -2350 -1200
rect -2330 -1220 -2310 -1200
rect -2290 -1220 -2270 -1200
rect -2250 -1220 -2230 -1200
rect -2210 -1220 -2190 -1200
rect -2170 -1220 -2150 -1200
rect -2130 -1220 -2110 -1200
rect -2090 -1220 -2070 -1200
rect -2050 -1220 -2030 -1200
rect -2010 -1220 -1990 -1200
rect -1970 -1220 -1950 -1200
rect -1930 -1220 -1910 -1200
rect -1890 -1220 -1870 -1200
rect -1850 -1220 -1830 -1200
rect -1810 -1220 -1790 -1200
rect -1770 -1220 -1750 -1200
rect -1730 -1220 -1710 -1200
rect -1690 -1220 -1670 -1200
rect -1650 -1220 -1630 -1200
rect -1610 -1220 -1590 -1200
rect -1570 -1220 -1550 -1200
rect -1530 -1220 -1510 -1200
rect -1490 -1220 -1470 -1200
rect -1450 -1220 -1430 -1200
rect -1410 -1220 -1390 -1200
rect -1370 -1220 -1350 -1200
rect -1330 -1220 -1310 -1200
rect -1290 -1220 -1270 -1200
rect -1250 -1220 -1230 -1200
rect -1210 -1220 -1190 -1200
rect -1170 -1220 -1150 -1200
rect -1130 -1220 -1110 -1200
rect -1090 -1220 -1070 -1200
rect -1050 -1220 -1030 -1200
rect -1010 -1220 -990 -1200
rect -970 -1220 -950 -1200
rect -930 -1220 -910 -1200
rect -890 -1220 -870 -1200
rect -850 -1220 -830 -1200
rect -810 -1220 -790 -1200
rect -770 -1220 -750 -1200
rect -730 -1220 -710 -1200
rect -690 -1220 -670 -1200
rect -650 -1220 -630 -1200
rect -610 -1220 -590 -1200
rect -570 -1220 -550 -1200
rect -530 -1220 -510 -1200
rect -490 -1220 -470 -1200
rect -450 -1220 -430 -1200
rect -410 -1220 -390 -1200
rect -370 -1220 -350 -1200
rect -330 -1220 -310 -1200
rect -290 -1220 -270 -1200
rect -250 -1220 -230 -1200
rect -210 -1220 -190 -1200
rect -170 -1220 -150 -1200
rect -130 -1220 -110 -1200
rect -90 -1220 -70 -1200
rect -50 -1220 -30 -1200
rect -10 -1220 10 -1200
rect 30 -1220 50 -1200
rect 80 -1220 100 -1200
rect 120 -1220 140 -1200
rect 160 -1220 180 -1200
rect 200 -1220 220 -1200
rect 240 -1220 260 -1200
rect 280 -1220 300 -1200
rect 320 -1220 340 -1200
rect 360 -1220 380 -1200
rect 400 -1220 420 -1200
rect 440 -1220 460 -1200
rect 480 -1220 500 -1200
rect 520 -1220 540 -1200
rect 560 -1220 580 -1200
rect 600 -1220 620 -1200
rect 640 -1220 660 -1200
rect 680 -1220 700 -1200
rect 720 -1220 740 -1200
rect 760 -1220 780 -1200
rect 800 -1220 820 -1200
rect 840 -1220 860 -1200
rect 880 -1220 900 -1200
rect 920 -1220 940 -1200
rect 960 -1220 980 -1200
rect 1000 -1220 1020 -1200
rect 1040 -1220 1060 -1200
rect 1080 -1220 1100 -1200
rect 1120 -1220 1140 -1200
rect 1160 -1220 1180 -1200
rect 1200 -1220 1220 -1200
rect 1240 -1220 1260 -1200
rect 1280 -1220 1300 -1200
rect 1320 -1220 1340 -1200
rect 1360 -1220 1380 -1200
rect 1400 -1220 1420 -1200
rect 1440 -1220 1460 -1200
rect 1480 -1220 1500 -1200
rect 1520 -1220 1540 -1200
rect 1560 -1220 1580 -1200
rect 1600 -1220 1620 -1200
rect 1640 -1220 1660 -1200
rect 1680 -1220 1700 -1200
rect 1720 -1220 1740 -1200
rect 1760 -1220 1780 -1200
rect 1800 -1220 1820 -1200
rect 1840 -1220 1860 -1200
rect 1880 -1220 1900 -1200
rect 1920 -1220 1940 -1200
rect 1960 -1220 1980 -1200
rect 2000 -1220 2020 -1200
rect 2040 -1220 2060 -1200
rect 2080 -1220 2100 -1200
rect 2120 -1220 2140 -1200
rect 2160 -1220 2180 -1200
rect 2200 -1220 2220 -1200
rect 2240 -1220 2260 -1200
rect 2280 -1220 2300 -1200
rect 2320 -1220 2340 -1200
rect 2360 -1220 2380 -1200
rect 2400 -1220 2420 -1200
rect 2440 -1220 2460 -1200
rect 2480 -1220 2500 -1200
rect 2520 -1220 2540 -1200
rect 2560 -1220 2580 -1200
rect 2600 -1220 2620 -1200
rect 2640 -1220 2660 -1200
rect 2680 -1220 2700 -1200
rect 2720 -1220 2740 -1200
rect 2760 -1220 2780 -1200
rect 2800 -1220 2820 -1200
rect 2840 -1220 2860 -1200
rect 2880 -1220 2900 -1200
rect 2920 -1220 2940 -1200
rect 2960 -1220 2980 -1200
rect 3000 -1220 3020 -1200
rect 3040 -1220 3060 -1200
rect 3080 -1220 3100 -1200
rect 3120 -1220 3140 -1200
rect 3160 -1220 3180 -1200
rect 3200 -1220 3220 -1200
rect 3240 -1220 3260 -1200
rect 3280 -1220 3300 -1200
rect 3320 -1220 3340 -1200
rect 3360 -1220 3380 -1200
rect 3400 -1220 3420 -1200
rect 3440 -1220 3460 -1200
rect 3480 -1220 3500 -1200
rect 3520 -1220 3540 -1200
rect 3560 -1220 3580 -1200
rect 3600 -1220 3615 -1200
rect -3485 -1230 3615 -1220
<< viali >>
rect -3110 -140 -3090 -120
rect -3070 -140 -3050 -120
rect -3030 -140 -3010 -120
rect -2990 -140 -2970 -120
rect -2950 -140 -2930 -120
rect -2910 -140 -2890 -120
rect -2870 -140 -2850 -120
rect -2830 -140 -2810 -120
rect -2790 -140 -2770 -120
rect -2750 -140 -2730 -120
rect -2710 -140 -2690 -120
rect -2670 -140 -2650 -120
rect -2630 -140 -2610 -120
rect -2590 -140 -2570 -120
rect -2550 -140 -2530 -120
rect -2510 -140 -2490 -120
rect -2470 -140 -2450 -120
rect -2430 -140 -2410 -120
rect -2390 -140 -2370 -120
rect -2350 -140 -2330 -120
rect 2460 -140 2480 -120
rect 2500 -140 2520 -120
rect 2540 -140 2560 -120
rect 2580 -140 2600 -120
rect 2620 -140 2640 -120
rect 2660 -140 2680 -120
rect 2700 -140 2720 -120
rect 2740 -140 2760 -120
rect 2780 -140 2800 -120
rect 2820 -140 2840 -120
rect 2860 -140 2880 -120
rect 2900 -140 2920 -120
rect 2940 -140 2960 -120
rect 2980 -140 3000 -120
rect 3020 -140 3040 -120
rect 3060 -140 3080 -120
rect 3100 -140 3120 -120
rect 3140 -140 3160 -120
rect 3180 -140 3200 -120
rect 3220 -140 3240 -120
rect -3110 -180 -3090 -160
rect -3070 -180 -3050 -160
rect -3030 -180 -3010 -160
rect -2990 -180 -2970 -160
rect -2950 -180 -2930 -160
rect -2910 -180 -2890 -160
rect -2870 -180 -2850 -160
rect -2830 -180 -2810 -160
rect -2790 -180 -2770 -160
rect -2750 -180 -2730 -160
rect -2710 -180 -2690 -160
rect -2670 -180 -2650 -160
rect -2630 -180 -2610 -160
rect -2590 -180 -2570 -160
rect -2550 -180 -2530 -160
rect -2510 -180 -2490 -160
rect -2470 -180 -2450 -160
rect -2430 -180 -2410 -160
rect -2390 -180 -2370 -160
rect -2350 -180 -2330 -160
rect 2460 -180 2480 -160
rect 2500 -180 2520 -160
rect 2540 -180 2560 -160
rect 2580 -180 2600 -160
rect 2620 -180 2640 -160
rect 2660 -180 2680 -160
rect 2700 -180 2720 -160
rect 2740 -180 2760 -160
rect 2780 -180 2800 -160
rect 2820 -180 2840 -160
rect 2860 -180 2880 -160
rect 2900 -180 2920 -160
rect 2940 -180 2960 -160
rect 2980 -180 3000 -160
rect 3020 -180 3040 -160
rect 3060 -180 3080 -160
rect 3100 -180 3120 -160
rect 3140 -180 3160 -160
rect 3180 -180 3200 -160
rect 3220 -180 3240 -160
rect 3645 -235 3665 -205
rect 3685 -235 3705 -205
rect 3725 -235 3745 -205
rect 3765 -235 3785 -205
rect -1040 -280 -1020 -260
rect -1000 -280 -980 -260
rect -960 -280 -940 -260
rect -920 -280 -900 -260
rect -880 -280 -860 -260
rect -840 -280 -820 -260
rect -800 -280 -780 -260
rect -760 -280 -740 -260
rect -720 -280 -700 -260
rect -680 -280 -660 -260
rect -640 -280 -620 -260
rect -600 -280 -580 -260
rect -560 -280 -540 -260
rect -520 -280 -500 -260
rect -480 -280 -460 -260
rect -440 -280 -420 -260
rect -400 -280 -380 -260
rect -360 -280 -340 -260
rect -320 -280 -300 -260
rect -280 -280 -260 -260
rect 390 -280 410 -260
rect 430 -280 450 -260
rect 470 -280 490 -260
rect 510 -280 530 -260
rect 550 -280 570 -260
rect 590 -280 610 -260
rect 630 -280 650 -260
rect 670 -280 690 -260
rect 710 -280 730 -260
rect 750 -280 770 -260
rect 790 -280 810 -260
rect 830 -280 850 -260
rect 870 -280 890 -260
rect 910 -280 930 -260
rect 950 -280 970 -260
rect 990 -280 1010 -260
rect 1030 -280 1050 -260
rect 1070 -280 1090 -260
rect 1110 -280 1130 -260
rect 1150 -280 1170 -260
rect 3645 -335 3665 -305
rect 3685 -335 3705 -305
rect 3725 -335 3745 -305
rect 3765 -335 3785 -305
rect -3110 -380 -3090 -360
rect -3070 -380 -3050 -360
rect -3030 -380 -3010 -360
rect -2990 -380 -2970 -360
rect -2950 -380 -2930 -360
rect -2910 -380 -2890 -360
rect -2870 -380 -2850 -360
rect -2830 -380 -2810 -360
rect -2790 -380 -2770 -360
rect -2750 -380 -2730 -360
rect -2710 -380 -2690 -360
rect -2670 -380 -2650 -360
rect -2630 -380 -2610 -360
rect -2590 -380 -2570 -360
rect -2550 -380 -2530 -360
rect -2510 -380 -2490 -360
rect -2470 -380 -2450 -360
rect -2430 -380 -2410 -360
rect -2390 -380 -2370 -360
rect -2350 -380 -2330 -360
rect 2460 -380 2480 -360
rect 2500 -380 2520 -360
rect 2540 -380 2560 -360
rect 2580 -380 2600 -360
rect 2620 -380 2640 -360
rect 2660 -380 2680 -360
rect 2700 -380 2720 -360
rect 2740 -380 2760 -360
rect 2780 -380 2800 -360
rect 2820 -380 2840 -360
rect 2860 -380 2880 -360
rect 2900 -380 2920 -360
rect 2940 -380 2960 -360
rect 2980 -380 3000 -360
rect 3020 -380 3040 -360
rect 3060 -380 3080 -360
rect 3100 -380 3120 -360
rect 3140 -380 3160 -360
rect 3180 -380 3200 -360
rect 3220 -380 3240 -360
rect 3645 -435 3665 -405
rect 3685 -435 3705 -405
rect 3725 -435 3745 -405
rect 3765 -435 3785 -405
rect -1040 -480 -1020 -460
rect -1000 -480 -980 -460
rect -960 -480 -940 -460
rect -920 -480 -900 -460
rect -880 -480 -860 -460
rect -840 -480 -820 -460
rect -800 -480 -780 -460
rect -760 -480 -740 -460
rect -720 -480 -700 -460
rect -680 -480 -660 -460
rect -640 -480 -620 -460
rect -600 -480 -580 -460
rect -560 -480 -540 -460
rect -520 -480 -500 -460
rect -480 -480 -460 -460
rect -440 -480 -420 -460
rect -400 -480 -380 -460
rect -360 -480 -340 -460
rect -320 -480 -300 -460
rect -280 -480 -260 -460
rect 390 -480 410 -460
rect 430 -480 450 -460
rect 470 -480 490 -460
rect 510 -480 530 -460
rect 550 -480 570 -460
rect 590 -480 610 -460
rect 630 -480 650 -460
rect 670 -480 690 -460
rect 710 -480 730 -460
rect 750 -480 770 -460
rect 790 -480 810 -460
rect 830 -480 850 -460
rect 870 -480 890 -460
rect 910 -480 930 -460
rect 950 -480 970 -460
rect 990 -480 1010 -460
rect 1030 -480 1050 -460
rect 1070 -480 1090 -460
rect 1110 -480 1130 -460
rect 1150 -480 1170 -460
rect 3645 -535 3665 -505
rect 3685 -535 3705 -505
rect 3725 -535 3745 -505
rect 3765 -535 3785 -505
rect -3110 -580 -3090 -560
rect -3070 -580 -3050 -560
rect -3030 -580 -3010 -560
rect -2990 -580 -2970 -560
rect -2950 -580 -2930 -560
rect -2910 -580 -2890 -560
rect -2870 -580 -2850 -560
rect -2830 -580 -2810 -560
rect -2790 -580 -2770 -560
rect -2750 -580 -2730 -560
rect -2710 -580 -2690 -560
rect -2670 -580 -2650 -560
rect -2630 -580 -2610 -560
rect -2590 -580 -2570 -560
rect -2550 -580 -2530 -560
rect -2510 -580 -2490 -560
rect -2470 -580 -2450 -560
rect -2430 -580 -2410 -560
rect -2390 -580 -2370 -560
rect -2350 -580 -2330 -560
rect 2460 -580 2480 -560
rect 2500 -580 2520 -560
rect 2540 -580 2560 -560
rect 2580 -580 2600 -560
rect 2620 -580 2640 -560
rect 2660 -580 2680 -560
rect 2700 -580 2720 -560
rect 2740 -580 2760 -560
rect 2780 -580 2800 -560
rect 2820 -580 2840 -560
rect 2860 -580 2880 -560
rect 2900 -580 2920 -560
rect 2940 -580 2960 -560
rect 2980 -580 3000 -560
rect 3020 -580 3040 -560
rect 3060 -580 3080 -560
rect 3100 -580 3120 -560
rect 3140 -580 3160 -560
rect 3180 -580 3200 -560
rect 3220 -580 3240 -560
rect 3645 -635 3665 -605
rect 3685 -635 3705 -605
rect 3725 -635 3745 -605
rect 3765 -635 3785 -605
rect -1040 -680 -1020 -660
rect -1000 -680 -980 -660
rect -960 -680 -940 -660
rect -920 -680 -900 -660
rect -880 -680 -860 -660
rect -840 -680 -820 -660
rect -800 -680 -780 -660
rect -760 -680 -740 -660
rect -720 -680 -700 -660
rect -680 -680 -660 -660
rect -640 -680 -620 -660
rect -600 -680 -580 -660
rect -560 -680 -540 -660
rect -520 -680 -500 -660
rect -480 -680 -460 -660
rect -440 -680 -420 -660
rect -400 -680 -380 -660
rect -360 -680 -340 -660
rect -320 -680 -300 -660
rect -280 -680 -260 -660
rect 390 -680 410 -660
rect 430 -680 450 -660
rect 470 -680 490 -660
rect 510 -680 530 -660
rect 550 -680 570 -660
rect 590 -680 610 -660
rect 630 -680 650 -660
rect 670 -680 690 -660
rect 710 -680 730 -660
rect 750 -680 770 -660
rect 790 -680 810 -660
rect 830 -680 850 -660
rect 870 -680 890 -660
rect 910 -680 930 -660
rect 950 -680 970 -660
rect 990 -680 1010 -660
rect 1030 -680 1050 -660
rect 1070 -680 1090 -660
rect 1110 -680 1130 -660
rect 1150 -680 1170 -660
rect 3645 -735 3665 -705
rect 3685 -735 3705 -705
rect 3725 -735 3745 -705
rect 3765 -735 3785 -705
rect -3110 -780 -3090 -760
rect -3070 -780 -3050 -760
rect -3030 -780 -3010 -760
rect -2990 -780 -2970 -760
rect -2950 -780 -2930 -760
rect -2910 -780 -2890 -760
rect -2870 -780 -2850 -760
rect -2830 -780 -2810 -760
rect -2790 -780 -2770 -760
rect -2750 -780 -2730 -760
rect -2710 -780 -2690 -760
rect -2670 -780 -2650 -760
rect -2630 -780 -2610 -760
rect -2590 -780 -2570 -760
rect -2550 -780 -2530 -760
rect -2510 -780 -2490 -760
rect -2470 -780 -2450 -760
rect -2430 -780 -2410 -760
rect -2390 -780 -2370 -760
rect -2350 -780 -2330 -760
rect 2460 -780 2480 -760
rect 2500 -780 2520 -760
rect 2540 -780 2560 -760
rect 2580 -780 2600 -760
rect 2620 -780 2640 -760
rect 2660 -780 2680 -760
rect 2700 -780 2720 -760
rect 2740 -780 2760 -760
rect 2780 -780 2800 -760
rect 2820 -780 2840 -760
rect 2860 -780 2880 -760
rect 2900 -780 2920 -760
rect 2940 -780 2960 -760
rect 2980 -780 3000 -760
rect 3020 -780 3040 -760
rect 3060 -780 3080 -760
rect 3100 -780 3120 -760
rect 3140 -780 3160 -760
rect 3180 -780 3200 -760
rect 3220 -780 3240 -760
rect 3645 -835 3665 -805
rect 3685 -835 3705 -805
rect 3725 -835 3745 -805
rect 3765 -835 3785 -805
rect -1040 -880 -1020 -860
rect -1000 -880 -980 -860
rect -960 -880 -940 -860
rect -920 -880 -900 -860
rect -880 -880 -860 -860
rect -840 -880 -820 -860
rect -800 -880 -780 -860
rect -760 -880 -740 -860
rect -720 -880 -700 -860
rect -680 -880 -660 -860
rect -640 -880 -620 -860
rect -600 -880 -580 -860
rect -560 -880 -540 -860
rect -520 -880 -500 -860
rect -480 -880 -460 -860
rect -440 -880 -420 -860
rect -400 -880 -380 -860
rect -360 -880 -340 -860
rect -320 -880 -300 -860
rect -280 -880 -260 -860
rect 390 -880 410 -860
rect 430 -880 450 -860
rect 470 -880 490 -860
rect 510 -880 530 -860
rect 550 -880 570 -860
rect 590 -880 610 -860
rect 630 -880 650 -860
rect 670 -880 690 -860
rect 710 -880 730 -860
rect 750 -880 770 -860
rect 790 -880 810 -860
rect 830 -880 850 -860
rect 870 -880 890 -860
rect 910 -880 930 -860
rect 950 -880 970 -860
rect 990 -880 1010 -860
rect 1030 -880 1050 -860
rect 1070 -880 1090 -860
rect 1110 -880 1130 -860
rect 1150 -880 1170 -860
rect 3645 -935 3665 -905
rect 3685 -935 3705 -905
rect 3725 -935 3745 -905
rect 3765 -935 3785 -905
rect -3110 -980 -3090 -960
rect -3070 -980 -3050 -960
rect -3030 -980 -3010 -960
rect -2990 -980 -2970 -960
rect -2950 -980 -2930 -960
rect -2910 -980 -2890 -960
rect -2870 -980 -2850 -960
rect -2830 -980 -2810 -960
rect -2790 -980 -2770 -960
rect -2750 -980 -2730 -960
rect -2710 -980 -2690 -960
rect -2670 -980 -2650 -960
rect -2630 -980 -2610 -960
rect -2590 -980 -2570 -960
rect -2550 -980 -2530 -960
rect -2510 -980 -2490 -960
rect -2470 -980 -2450 -960
rect -2430 -980 -2410 -960
rect -2390 -980 -2370 -960
rect -2350 -980 -2330 -960
rect 2460 -980 2480 -960
rect 2500 -980 2520 -960
rect 2540 -980 2560 -960
rect 2580 -980 2600 -960
rect 2620 -980 2640 -960
rect 2660 -980 2680 -960
rect 2700 -980 2720 -960
rect 2740 -980 2760 -960
rect 2780 -980 2800 -960
rect 2820 -980 2840 -960
rect 2860 -980 2880 -960
rect 2900 -980 2920 -960
rect 2940 -980 2960 -960
rect 2980 -980 3000 -960
rect 3020 -980 3040 -960
rect 3060 -980 3080 -960
rect 3100 -980 3120 -960
rect 3140 -980 3160 -960
rect 3180 -980 3200 -960
rect 3220 -980 3240 -960
rect 3645 -1035 3665 -1005
rect 3685 -1035 3705 -1005
rect 3725 -1035 3745 -1005
rect 3765 -1035 3785 -1005
rect -1040 -1080 -1020 -1060
rect -1000 -1080 -980 -1060
rect -960 -1080 -940 -1060
rect -920 -1080 -900 -1060
rect -880 -1080 -860 -1060
rect -840 -1080 -820 -1060
rect -800 -1080 -780 -1060
rect -760 -1080 -740 -1060
rect -720 -1080 -700 -1060
rect -680 -1080 -660 -1060
rect -640 -1080 -620 -1060
rect -600 -1080 -580 -1060
rect -560 -1080 -540 -1060
rect -520 -1080 -500 -1060
rect -480 -1080 -460 -1060
rect -440 -1080 -420 -1060
rect -400 -1080 -380 -1060
rect -360 -1080 -340 -1060
rect -320 -1080 -300 -1060
rect -280 -1080 -260 -1060
rect 390 -1080 410 -1060
rect 430 -1080 450 -1060
rect 470 -1080 490 -1060
rect 510 -1080 530 -1060
rect 550 -1080 570 -1060
rect 590 -1080 610 -1060
rect 630 -1080 650 -1060
rect 670 -1080 690 -1060
rect 710 -1080 730 -1060
rect 750 -1080 770 -1060
rect 790 -1080 810 -1060
rect 830 -1080 850 -1060
rect 870 -1080 890 -1060
rect 910 -1080 930 -1060
rect 950 -1080 970 -1060
rect 990 -1080 1010 -1060
rect 1030 -1080 1050 -1060
rect 1070 -1080 1090 -1060
rect 1110 -1080 1130 -1060
rect 1150 -1080 1170 -1060
rect 3645 -1135 3665 -1105
rect 3685 -1135 3705 -1105
rect 3725 -1135 3745 -1105
rect 3765 -1135 3785 -1105
rect -3110 -1180 -3090 -1160
rect -3070 -1180 -3050 -1160
rect -3030 -1180 -3010 -1160
rect -2990 -1180 -2970 -1160
rect -2950 -1180 -2930 -1160
rect -2910 -1180 -2890 -1160
rect -2870 -1180 -2850 -1160
rect -2830 -1180 -2810 -1160
rect -2790 -1180 -2770 -1160
rect -2750 -1180 -2730 -1160
rect -2710 -1180 -2690 -1160
rect -2670 -1180 -2650 -1160
rect -2630 -1180 -2610 -1160
rect -2590 -1180 -2570 -1160
rect -2550 -1180 -2530 -1160
rect -2510 -1180 -2490 -1160
rect -2470 -1180 -2450 -1160
rect -2430 -1180 -2410 -1160
rect -2390 -1180 -2370 -1160
rect -2350 -1180 -2330 -1160
rect 2460 -1180 2480 -1160
rect 2500 -1180 2520 -1160
rect 2540 -1180 2560 -1160
rect 2580 -1180 2600 -1160
rect 2620 -1180 2640 -1160
rect 2660 -1180 2680 -1160
rect 2700 -1180 2720 -1160
rect 2740 -1180 2760 -1160
rect 2780 -1180 2800 -1160
rect 2820 -1180 2840 -1160
rect 2860 -1180 2880 -1160
rect 2900 -1180 2920 -1160
rect 2940 -1180 2960 -1160
rect 2980 -1180 3000 -1160
rect 3020 -1180 3040 -1160
rect 3060 -1180 3080 -1160
rect 3100 -1180 3120 -1160
rect 3140 -1180 3160 -1160
rect 3180 -1180 3200 -1160
rect 3220 -1180 3240 -1160
rect -3110 -1220 -3090 -1200
rect -3070 -1220 -3050 -1200
rect -3030 -1220 -3010 -1200
rect -2990 -1220 -2970 -1200
rect -2950 -1220 -2930 -1200
rect -2910 -1220 -2890 -1200
rect -2870 -1220 -2850 -1200
rect -2830 -1220 -2810 -1200
rect -2790 -1220 -2770 -1200
rect -2750 -1220 -2730 -1200
rect -2710 -1220 -2690 -1200
rect -2670 -1220 -2650 -1200
rect -2630 -1220 -2610 -1200
rect -2590 -1220 -2570 -1200
rect -2550 -1220 -2530 -1200
rect -2510 -1220 -2490 -1200
rect -2470 -1220 -2450 -1200
rect -2430 -1220 -2410 -1200
rect -2390 -1220 -2370 -1200
rect -2350 -1220 -2330 -1200
rect 2460 -1220 2480 -1200
rect 2500 -1220 2520 -1200
rect 2540 -1220 2560 -1200
rect 2580 -1220 2600 -1200
rect 2620 -1220 2640 -1200
rect 2660 -1220 2680 -1200
rect 2700 -1220 2720 -1200
rect 2740 -1220 2760 -1200
rect 2780 -1220 2800 -1200
rect 2820 -1220 2840 -1200
rect 2860 -1220 2880 -1200
rect 2900 -1220 2920 -1200
rect 2940 -1220 2960 -1200
rect 2980 -1220 3000 -1200
rect 3020 -1220 3040 -1200
rect 3060 -1220 3080 -1200
rect 3100 -1220 3120 -1200
rect 3140 -1220 3160 -1200
rect 3180 -1220 3200 -1200
rect 3220 -1220 3240 -1200
<< metal1 >>
rect -2575 2005 -2395 2020
rect 2220 2005 3020 2020
rect 15 1690 115 1930
rect 15 600 115 1660
rect -2490 -110 -2370 490
rect -1930 485 -1130 525
rect 1260 485 2060 525
rect -145 20 10 390
rect 120 20 275 390
rect -3120 -120 -2320 -110
rect -3120 -140 -3110 -120
rect -3090 -140 -3070 -120
rect -3050 -140 -3030 -120
rect -3010 -140 -2990 -120
rect -2970 -140 -2950 -120
rect -2930 -140 -2910 -120
rect -2890 -140 -2870 -120
rect -2850 -140 -2830 -120
rect -2810 -140 -2790 -120
rect -2770 -140 -2750 -120
rect -2730 -140 -2710 -120
rect -2690 -140 -2670 -120
rect -2650 -140 -2630 -120
rect -2610 -140 -2590 -120
rect -2570 -140 -2550 -120
rect -2530 -140 -2510 -120
rect -2490 -140 -2470 -120
rect -2450 -140 -2430 -120
rect -2410 -140 -2390 -120
rect -2370 -140 -2350 -120
rect -2330 -140 -2320 -120
rect -3120 -160 -2320 -140
rect -3120 -180 -3110 -160
rect -3090 -180 -3070 -160
rect -3050 -180 -3030 -160
rect -3010 -180 -2990 -160
rect -2970 -180 -2950 -160
rect -2930 -180 -2910 -160
rect -2890 -180 -2870 -160
rect -2850 -180 -2830 -160
rect -2810 -180 -2790 -160
rect -2770 -180 -2750 -160
rect -2730 -180 -2710 -160
rect -2690 -180 -2670 -160
rect -2650 -180 -2630 -160
rect -2610 -180 -2590 -160
rect -2570 -180 -2550 -160
rect -2530 -180 -2510 -160
rect -2490 -180 -2470 -160
rect -2450 -180 -2430 -160
rect -2410 -180 -2390 -160
rect -2370 -180 -2350 -160
rect -2330 -180 -2320 -160
rect -3120 -360 -2320 -180
rect -3120 -380 -3110 -360
rect -3090 -380 -3070 -360
rect -3050 -380 -3030 -360
rect -3010 -380 -2990 -360
rect -2970 -380 -2950 -360
rect -2930 -380 -2910 -360
rect -2890 -380 -2870 -360
rect -2850 -380 -2830 -360
rect -2810 -380 -2790 -360
rect -2770 -380 -2750 -360
rect -2730 -380 -2710 -360
rect -2690 -380 -2670 -360
rect -2650 -380 -2630 -360
rect -2610 -380 -2590 -360
rect -2570 -380 -2550 -360
rect -2530 -380 -2510 -360
rect -2490 -380 -2470 -360
rect -2450 -380 -2430 -360
rect -2410 -380 -2390 -360
rect -2370 -380 -2350 -360
rect -2330 -380 -2320 -360
rect -3120 -560 -2320 -380
rect -3120 -580 -3110 -560
rect -3090 -580 -3070 -560
rect -3050 -580 -3030 -560
rect -3010 -580 -2990 -560
rect -2970 -580 -2950 -560
rect -2930 -580 -2910 -560
rect -2890 -580 -2870 -560
rect -2850 -580 -2830 -560
rect -2810 -580 -2790 -560
rect -2770 -580 -2750 -560
rect -2730 -580 -2710 -560
rect -2690 -580 -2670 -560
rect -2650 -580 -2630 -560
rect -2610 -580 -2590 -560
rect -2570 -580 -2550 -560
rect -2530 -580 -2510 -560
rect -2490 -580 -2470 -560
rect -2450 -580 -2430 -560
rect -2410 -580 -2390 -560
rect -2370 -580 -2350 -560
rect -2330 -580 -2320 -560
rect -3120 -760 -2320 -580
rect -3120 -780 -3110 -760
rect -3090 -780 -3070 -760
rect -3050 -780 -3030 -760
rect -3010 -780 -2990 -760
rect -2970 -780 -2950 -760
rect -2930 -780 -2910 -760
rect -2890 -780 -2870 -760
rect -2850 -780 -2830 -760
rect -2810 -780 -2790 -760
rect -2770 -780 -2750 -760
rect -2730 -780 -2710 -760
rect -2690 -780 -2670 -760
rect -2650 -780 -2630 -760
rect -2610 -780 -2590 -760
rect -2570 -780 -2550 -760
rect -2530 -780 -2510 -760
rect -2490 -780 -2470 -760
rect -2450 -780 -2430 -760
rect -2410 -780 -2390 -760
rect -2370 -780 -2350 -760
rect -2330 -780 -2320 -760
rect -3120 -960 -2320 -780
rect -3120 -980 -3110 -960
rect -3090 -980 -3070 -960
rect -3050 -980 -3030 -960
rect -3010 -980 -2990 -960
rect -2970 -980 -2950 -960
rect -2930 -980 -2910 -960
rect -2890 -980 -2870 -960
rect -2850 -980 -2830 -960
rect -2810 -980 -2790 -960
rect -2770 -980 -2750 -960
rect -2730 -980 -2710 -960
rect -2690 -980 -2670 -960
rect -2650 -980 -2630 -960
rect -2610 -980 -2590 -960
rect -2570 -980 -2550 -960
rect -2530 -980 -2510 -960
rect -2490 -980 -2470 -960
rect -2450 -980 -2430 -960
rect -2410 -980 -2390 -960
rect -2370 -980 -2350 -960
rect -2330 -980 -2320 -960
rect -3120 -1160 -2320 -980
rect -1050 -260 -250 -95
rect -1050 -280 -1040 -260
rect -1020 -280 -1000 -260
rect -980 -280 -960 -260
rect -940 -280 -920 -260
rect -900 -280 -880 -260
rect -860 -280 -840 -260
rect -820 -280 -800 -260
rect -780 -280 -760 -260
rect -740 -280 -720 -260
rect -700 -280 -680 -260
rect -660 -280 -640 -260
rect -620 -280 -600 -260
rect -580 -280 -560 -260
rect -540 -280 -520 -260
rect -500 -280 -480 -260
rect -460 -280 -440 -260
rect -420 -280 -400 -260
rect -380 -280 -360 -260
rect -340 -280 -320 -260
rect -300 -280 -280 -260
rect -260 -280 -250 -260
rect -1050 -460 -250 -280
rect -1050 -480 -1040 -460
rect -1020 -480 -1000 -460
rect -980 -480 -960 -460
rect -940 -480 -920 -460
rect -900 -480 -880 -460
rect -860 -480 -840 -460
rect -820 -480 -800 -460
rect -780 -480 -760 -460
rect -740 -480 -720 -460
rect -700 -480 -680 -460
rect -660 -480 -640 -460
rect -620 -480 -600 -460
rect -580 -480 -560 -460
rect -540 -480 -520 -460
rect -500 -480 -480 -460
rect -460 -480 -440 -460
rect -420 -480 -400 -460
rect -380 -480 -360 -460
rect -340 -480 -320 -460
rect -300 -480 -280 -460
rect -260 -480 -250 -460
rect -1050 -660 -250 -480
rect -1050 -680 -1040 -660
rect -1020 -680 -1000 -660
rect -980 -680 -960 -660
rect -940 -680 -920 -660
rect -900 -680 -880 -660
rect -860 -680 -840 -660
rect -820 -680 -800 -660
rect -780 -680 -760 -660
rect -740 -680 -720 -660
rect -700 -680 -680 -660
rect -660 -680 -640 -660
rect -620 -680 -600 -660
rect -580 -680 -560 -660
rect -540 -680 -520 -660
rect -500 -680 -480 -660
rect -460 -680 -440 -660
rect -420 -680 -400 -660
rect -380 -680 -360 -660
rect -340 -680 -320 -660
rect -300 -680 -280 -660
rect -260 -680 -250 -660
rect -1050 -860 -250 -680
rect -1050 -880 -1040 -860
rect -1020 -880 -1000 -860
rect -980 -880 -960 -860
rect -940 -880 -920 -860
rect -900 -880 -880 -860
rect -860 -880 -840 -860
rect -820 -880 -800 -860
rect -780 -880 -760 -860
rect -740 -880 -720 -860
rect -700 -880 -680 -860
rect -660 -880 -640 -860
rect -620 -880 -600 -860
rect -580 -880 -560 -860
rect -540 -880 -520 -860
rect -500 -880 -480 -860
rect -460 -880 -440 -860
rect -420 -880 -400 -860
rect -380 -880 -360 -860
rect -340 -880 -320 -860
rect -300 -880 -280 -860
rect -260 -880 -250 -860
rect -1050 -1060 -250 -880
rect -1050 -1080 -1040 -1060
rect -1020 -1080 -1000 -1060
rect -980 -1080 -960 -1060
rect -940 -1080 -920 -1060
rect -900 -1080 -880 -1060
rect -860 -1080 -840 -1060
rect -820 -1080 -800 -1060
rect -780 -1080 -760 -1060
rect -740 -1080 -720 -1060
rect -700 -1080 -680 -1060
rect -660 -1080 -640 -1060
rect -620 -1080 -600 -1060
rect -580 -1080 -560 -1060
rect -540 -1080 -520 -1060
rect -500 -1080 -480 -1060
rect -460 -1080 -440 -1060
rect -420 -1080 -400 -1060
rect -380 -1080 -360 -1060
rect -340 -1080 -320 -1060
rect -300 -1080 -280 -1060
rect -260 -1080 -250 -1060
rect -1050 -1150 -250 -1080
rect 380 -260 1180 -95
rect 2500 -110 2620 490
rect 380 -280 390 -260
rect 410 -280 430 -260
rect 450 -280 470 -260
rect 490 -280 510 -260
rect 530 -280 550 -260
rect 570 -280 590 -260
rect 610 -280 630 -260
rect 650 -280 670 -260
rect 690 -280 710 -260
rect 730 -280 750 -260
rect 770 -280 790 -260
rect 810 -280 830 -260
rect 850 -280 870 -260
rect 890 -280 910 -260
rect 930 -280 950 -260
rect 970 -280 990 -260
rect 1010 -280 1030 -260
rect 1050 -280 1070 -260
rect 1090 -280 1110 -260
rect 1130 -280 1150 -260
rect 1170 -280 1180 -260
rect 380 -460 1180 -280
rect 380 -480 390 -460
rect 410 -480 430 -460
rect 450 -480 470 -460
rect 490 -480 510 -460
rect 530 -480 550 -460
rect 570 -480 590 -460
rect 610 -480 630 -460
rect 650 -480 670 -460
rect 690 -480 710 -460
rect 730 -480 750 -460
rect 770 -480 790 -460
rect 810 -480 830 -460
rect 850 -480 870 -460
rect 890 -480 910 -460
rect 930 -480 950 -460
rect 970 -480 990 -460
rect 1010 -480 1030 -460
rect 1050 -480 1070 -460
rect 1090 -480 1110 -460
rect 1130 -480 1150 -460
rect 1170 -480 1180 -460
rect 380 -660 1180 -480
rect 380 -680 390 -660
rect 410 -680 430 -660
rect 450 -680 470 -660
rect 490 -680 510 -660
rect 530 -680 550 -660
rect 570 -680 590 -660
rect 610 -680 630 -660
rect 650 -680 670 -660
rect 690 -680 710 -660
rect 730 -680 750 -660
rect 770 -680 790 -660
rect 810 -680 830 -660
rect 850 -680 870 -660
rect 890 -680 910 -660
rect 930 -680 950 -660
rect 970 -680 990 -660
rect 1010 -680 1030 -660
rect 1050 -680 1070 -660
rect 1090 -680 1110 -660
rect 1130 -680 1150 -660
rect 1170 -680 1180 -660
rect 380 -860 1180 -680
rect 380 -880 390 -860
rect 410 -880 430 -860
rect 450 -880 470 -860
rect 490 -880 510 -860
rect 530 -880 550 -860
rect 570 -880 590 -860
rect 610 -880 630 -860
rect 650 -880 670 -860
rect 690 -880 710 -860
rect 730 -880 750 -860
rect 770 -880 790 -860
rect 810 -880 830 -860
rect 850 -880 870 -860
rect 890 -880 910 -860
rect 930 -880 950 -860
rect 970 -880 990 -860
rect 1010 -880 1030 -860
rect 1050 -880 1070 -860
rect 1090 -880 1110 -860
rect 1130 -880 1150 -860
rect 1170 -880 1180 -860
rect 380 -1060 1180 -880
rect 380 -1080 390 -1060
rect 410 -1080 430 -1060
rect 450 -1080 470 -1060
rect 490 -1080 510 -1060
rect 530 -1080 550 -1060
rect 570 -1080 590 -1060
rect 610 -1080 630 -1060
rect 650 -1080 670 -1060
rect 690 -1080 710 -1060
rect 730 -1080 750 -1060
rect 770 -1080 790 -1060
rect 810 -1080 830 -1060
rect 850 -1080 870 -1060
rect 890 -1080 910 -1060
rect 930 -1080 950 -1060
rect 970 -1080 990 -1060
rect 1010 -1080 1030 -1060
rect 1050 -1080 1070 -1060
rect 1090 -1080 1110 -1060
rect 1130 -1080 1150 -1060
rect 1170 -1080 1180 -1060
rect 380 -1150 1180 -1080
rect 2450 -120 3250 -110
rect 2450 -140 2460 -120
rect 2480 -140 2500 -120
rect 2520 -140 2540 -120
rect 2560 -140 2580 -120
rect 2600 -140 2620 -120
rect 2640 -140 2660 -120
rect 2680 -140 2700 -120
rect 2720 -140 2740 -120
rect 2760 -140 2780 -120
rect 2800 -140 2820 -120
rect 2840 -140 2860 -120
rect 2880 -140 2900 -120
rect 2920 -140 2940 -120
rect 2960 -140 2980 -120
rect 3000 -140 3020 -120
rect 3040 -140 3060 -120
rect 3080 -140 3100 -120
rect 3120 -140 3140 -120
rect 3160 -140 3180 -120
rect 3200 -140 3220 -120
rect 3240 -140 3250 -120
rect 2450 -160 3250 -140
rect 2450 -180 2460 -160
rect 2480 -180 2500 -160
rect 2520 -180 2540 -160
rect 2560 -180 2580 -160
rect 2600 -180 2620 -160
rect 2640 -180 2660 -160
rect 2680 -180 2700 -160
rect 2720 -180 2740 -160
rect 2760 -180 2780 -160
rect 2800 -180 2820 -160
rect 2840 -180 2860 -160
rect 2880 -180 2900 -160
rect 2920 -180 2940 -160
rect 2960 -180 2980 -160
rect 3000 -180 3020 -160
rect 3040 -180 3060 -160
rect 3080 -180 3100 -160
rect 3120 -180 3140 -160
rect 3160 -180 3180 -160
rect 3200 -180 3220 -160
rect 3240 -180 3250 -160
rect 2450 -360 3250 -180
rect 2450 -380 2460 -360
rect 2480 -380 2500 -360
rect 2520 -380 2540 -360
rect 2560 -380 2580 -360
rect 2600 -380 2620 -360
rect 2640 -380 2660 -360
rect 2680 -380 2700 -360
rect 2720 -380 2740 -360
rect 2760 -380 2780 -360
rect 2800 -380 2820 -360
rect 2840 -380 2860 -360
rect 2880 -380 2900 -360
rect 2920 -380 2940 -360
rect 2960 -380 2980 -360
rect 3000 -380 3020 -360
rect 3040 -380 3060 -360
rect 3080 -380 3100 -360
rect 3120 -380 3140 -360
rect 3160 -380 3180 -360
rect 3200 -380 3220 -360
rect 3240 -380 3250 -360
rect 2450 -560 3250 -380
rect 2450 -580 2460 -560
rect 2480 -580 2500 -560
rect 2520 -580 2540 -560
rect 2560 -580 2580 -560
rect 2600 -580 2620 -560
rect 2640 -580 2660 -560
rect 2680 -580 2700 -560
rect 2720 -580 2740 -560
rect 2760 -580 2780 -560
rect 2800 -580 2820 -560
rect 2840 -580 2860 -560
rect 2880 -580 2900 -560
rect 2920 -580 2940 -560
rect 2960 -580 2980 -560
rect 3000 -580 3020 -560
rect 3040 -580 3060 -560
rect 3080 -580 3100 -560
rect 3120 -580 3140 -560
rect 3160 -580 3180 -560
rect 3200 -580 3220 -560
rect 3240 -580 3250 -560
rect 2450 -760 3250 -580
rect 2450 -780 2460 -760
rect 2480 -780 2500 -760
rect 2520 -780 2540 -760
rect 2560 -780 2580 -760
rect 2600 -780 2620 -760
rect 2640 -780 2660 -760
rect 2680 -780 2700 -760
rect 2720 -780 2740 -760
rect 2760 -780 2780 -760
rect 2800 -780 2820 -760
rect 2840 -780 2860 -760
rect 2880 -780 2900 -760
rect 2920 -780 2940 -760
rect 2960 -780 2980 -760
rect 3000 -780 3020 -760
rect 3040 -780 3060 -760
rect 3080 -780 3100 -760
rect 3120 -780 3140 -760
rect 3160 -780 3180 -760
rect 3200 -780 3220 -760
rect 3240 -780 3250 -760
rect 2450 -960 3250 -780
rect 2450 -980 2460 -960
rect 2480 -980 2500 -960
rect 2520 -980 2540 -960
rect 2560 -980 2580 -960
rect 2600 -980 2620 -960
rect 2640 -980 2660 -960
rect 2680 -980 2700 -960
rect 2720 -980 2740 -960
rect 2760 -980 2780 -960
rect 2800 -980 2820 -960
rect 2840 -980 2860 -960
rect 2880 -980 2900 -960
rect 2920 -980 2940 -960
rect 2960 -980 2980 -960
rect 3000 -980 3020 -960
rect 3040 -980 3060 -960
rect 3080 -980 3100 -960
rect 3120 -980 3140 -960
rect 3160 -980 3180 -960
rect 3200 -980 3220 -960
rect 3240 -980 3250 -960
rect -3120 -1180 -3110 -1160
rect -3090 -1180 -3070 -1160
rect -3050 -1180 -3030 -1160
rect -3010 -1180 -2990 -1160
rect -2970 -1180 -2950 -1160
rect -2930 -1180 -2910 -1160
rect -2890 -1180 -2870 -1160
rect -2850 -1180 -2830 -1160
rect -2810 -1180 -2790 -1160
rect -2770 -1180 -2750 -1160
rect -2730 -1180 -2710 -1160
rect -2690 -1180 -2670 -1160
rect -2650 -1180 -2630 -1160
rect -2610 -1180 -2590 -1160
rect -2570 -1180 -2550 -1160
rect -2530 -1180 -2510 -1160
rect -2490 -1180 -2470 -1160
rect -2450 -1180 -2430 -1160
rect -2410 -1180 -2390 -1160
rect -2370 -1180 -2350 -1160
rect -2330 -1180 -2320 -1160
rect -3120 -1200 -2320 -1180
rect -3120 -1220 -3110 -1200
rect -3090 -1220 -3070 -1200
rect -3050 -1220 -3030 -1200
rect -3010 -1220 -2990 -1200
rect -2970 -1220 -2950 -1200
rect -2930 -1220 -2910 -1200
rect -2890 -1220 -2870 -1200
rect -2850 -1220 -2830 -1200
rect -2810 -1220 -2790 -1200
rect -2770 -1220 -2750 -1200
rect -2730 -1220 -2710 -1200
rect -2690 -1220 -2670 -1200
rect -2650 -1220 -2630 -1200
rect -2610 -1220 -2590 -1200
rect -2570 -1220 -2550 -1200
rect -2530 -1220 -2510 -1200
rect -2490 -1220 -2470 -1200
rect -2450 -1220 -2430 -1200
rect -2410 -1220 -2390 -1200
rect -2370 -1220 -2350 -1200
rect -2330 -1220 -2320 -1200
rect -3120 -1245 -2320 -1220
rect 2450 -1160 3250 -980
rect 3635 -205 3790 -195
rect 3635 -235 3645 -205
rect 3665 -235 3685 -205
rect 3705 -235 3725 -205
rect 3745 -235 3765 -205
rect 3785 -235 3790 -205
rect 3635 -305 3790 -235
rect 3635 -335 3645 -305
rect 3665 -335 3685 -305
rect 3705 -335 3725 -305
rect 3745 -335 3765 -305
rect 3785 -335 3790 -305
rect 3635 -405 3790 -335
rect 3635 -435 3645 -405
rect 3665 -435 3685 -405
rect 3705 -435 3725 -405
rect 3745 -435 3765 -405
rect 3785 -435 3790 -405
rect 3635 -505 3790 -435
rect 3635 -535 3645 -505
rect 3665 -535 3685 -505
rect 3705 -535 3725 -505
rect 3745 -535 3765 -505
rect 3785 -535 3790 -505
rect 3635 -605 3790 -535
rect 3635 -635 3645 -605
rect 3665 -635 3685 -605
rect 3705 -635 3725 -605
rect 3745 -635 3765 -605
rect 3785 -635 3790 -605
rect 3635 -705 3790 -635
rect 3635 -735 3645 -705
rect 3665 -735 3685 -705
rect 3705 -735 3725 -705
rect 3745 -735 3765 -705
rect 3785 -735 3790 -705
rect 3635 -805 3790 -735
rect 3635 -835 3645 -805
rect 3665 -835 3685 -805
rect 3705 -835 3725 -805
rect 3745 -835 3765 -805
rect 3785 -835 3790 -805
rect 3635 -905 3790 -835
rect 3635 -935 3645 -905
rect 3665 -935 3685 -905
rect 3705 -935 3725 -905
rect 3745 -935 3765 -905
rect 3785 -935 3790 -905
rect 3635 -1005 3790 -935
rect 3635 -1035 3645 -1005
rect 3665 -1035 3685 -1005
rect 3705 -1035 3725 -1005
rect 3745 -1035 3765 -1005
rect 3785 -1035 3790 -1005
rect 3635 -1105 3790 -1035
rect 3635 -1135 3645 -1105
rect 3665 -1135 3685 -1105
rect 3705 -1135 3725 -1105
rect 3745 -1135 3765 -1105
rect 3785 -1135 3790 -1105
rect 3635 -1150 3790 -1135
rect 2450 -1180 2460 -1160
rect 2480 -1180 2500 -1160
rect 2520 -1180 2540 -1160
rect 2560 -1180 2580 -1160
rect 2600 -1180 2620 -1160
rect 2640 -1180 2660 -1160
rect 2680 -1180 2700 -1160
rect 2720 -1180 2740 -1160
rect 2760 -1180 2780 -1160
rect 2800 -1180 2820 -1160
rect 2840 -1180 2860 -1160
rect 2880 -1180 2900 -1160
rect 2920 -1180 2940 -1160
rect 2960 -1180 2980 -1160
rect 3000 -1180 3020 -1160
rect 3040 -1180 3060 -1160
rect 3080 -1180 3100 -1160
rect 3120 -1180 3140 -1160
rect 3160 -1180 3180 -1160
rect 3200 -1180 3220 -1160
rect 3240 -1180 3250 -1160
rect 2450 -1200 3250 -1180
rect 2450 -1220 2460 -1200
rect 2480 -1220 2500 -1200
rect 2520 -1220 2540 -1200
rect 2560 -1220 2580 -1200
rect 2600 -1220 2620 -1200
rect 2640 -1220 2660 -1200
rect 2680 -1220 2700 -1200
rect 2720 -1220 2740 -1200
rect 2760 -1220 2780 -1200
rect 2800 -1220 2820 -1200
rect 2840 -1220 2860 -1200
rect 2880 -1220 2900 -1200
rect 2920 -1220 2940 -1200
rect 2960 -1220 2980 -1200
rect 3000 -1220 3020 -1200
rect 3040 -1220 3060 -1200
rect 3080 -1220 3100 -1200
rect 3120 -1220 3140 -1200
rect 3160 -1220 3180 -1200
rect 3200 -1220 3220 -1200
rect 3240 -1220 3250 -1200
rect 2450 -1245 3250 -1220
use core_half  core_half_0
timestamp 1636159292
transform -1 0 -3650 0 1 560
box -3670 -655 -660 1470
use core_half  core_half_1
timestamp 1636159292
transform 1 0 3780 0 1 560
box -3670 -655 -660 1470
<< labels >>
rlabel metal1 2840 -1240 2840 -1240 1 GND
port 7 n
rlabel metal1 3650 -475 3650 -475 1 Vb1
port 15 n
rlabel metal1 -2740 -1240 -2740 -1240 1 GND
port 7 n
rlabel metal1 -30 205 -30 205 1 Vin_p
port 4 n
rlabel metal1 190 205 190 205 1 Vin_n
port 2 n
rlabel metal1 60 1825 60 1825 1 Vcmfb
port 14 n
rlabel metal1 60 1335 60 1335 1 Vb2
port 13 n
rlabel metal1 2590 2015 2590 2015 1 VDD#1
port 10 n
rlabel metal1 -2495 2015 -2495 2015 1 VDD
port 9 n
rlabel metal1 -1590 500 -1590 500 1 Vout_n
port 5 n
rlabel metal1 1660 495 1660 495 1 Vout_p
port 3 n
<< end >>
