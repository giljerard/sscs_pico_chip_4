magic
tech sky130A
magscale 1 2
timestamp 1637733805
<< xpolycontact >>
rect -1740 4130 -1600 4610
rect 16380 4130 16520 4610
rect -330 -380 150 -98
rect 7150 -380 7630 -98
rect 14630 -380 15110 -98
rect -1350 -4552 -870 -4270
rect -588 -4552 -110 -4270
rect 14890 -4552 15368 -4270
rect 15650 -4552 16130 -4270
rect -1740 -6950 -1600 -6470
rect 16380 -6950 16520 -6470
rect -270 -9900 210 -9618
rect 7210 -9900 7690 -9618
rect 14690 -9900 15170 -9618
<< xpolyres >>
rect -1740 -6470 -1600 4130
rect 150 -380 7150 -98
rect 7630 -380 14630 -98
rect -870 -4552 -588 -4270
rect 15368 -4552 15650 -4270
rect 16380 -6470 16520 4130
rect 210 -9900 7210 -9618
rect 7690 -9900 14690 -9618
<< viali >>
rect -1700 4550 -1640 4590
rect -1700 4470 -1640 4510
rect -1700 4390 -1640 4430
rect -1700 4310 -1640 4350
rect -1700 4230 -1640 4270
rect -1700 4150 -1640 4190
rect 16420 4550 16480 4590
rect 16420 4470 16480 4510
rect 16420 4390 16480 4430
rect 16420 4310 16480 4350
rect 16420 4230 16480 4270
rect 16420 4150 16480 4190
rect -310 -180 -270 -140
rect -230 -180 -190 -140
rect -150 -180 -110 -140
rect -70 -180 -30 -140
rect 10 -180 50 -140
rect 90 -180 130 -140
rect -310 -260 -270 -220
rect -230 -260 -190 -220
rect -150 -260 -110 -220
rect -70 -260 -30 -220
rect 10 -260 50 -220
rect 90 -260 130 -220
rect -310 -340 -270 -300
rect -230 -340 -190 -300
rect -150 -340 -110 -300
rect -70 -340 -30 -300
rect 10 -340 50 -300
rect 90 -340 130 -300
rect 7170 -180 7210 -140
rect 7250 -180 7290 -140
rect 7330 -180 7370 -140
rect 7410 -180 7450 -140
rect 7490 -180 7530 -140
rect 7570 -180 7610 -140
rect 7170 -260 7210 -220
rect 7250 -260 7290 -220
rect 7330 -260 7370 -220
rect 7410 -260 7450 -220
rect 7490 -260 7530 -220
rect 7570 -260 7610 -220
rect 7170 -340 7210 -300
rect 7250 -340 7290 -300
rect 7330 -340 7370 -300
rect 7410 -340 7450 -300
rect 7490 -340 7530 -300
rect 7570 -340 7610 -300
rect 14650 -180 14690 -140
rect 14730 -180 14770 -140
rect 14810 -180 14850 -140
rect 14890 -180 14930 -140
rect 14970 -180 15010 -140
rect 15050 -180 15090 -140
rect 14650 -260 14690 -220
rect 14730 -260 14770 -220
rect 14810 -260 14850 -220
rect 14890 -260 14930 -220
rect 14970 -260 15010 -220
rect 15050 -260 15090 -220
rect 14650 -340 14690 -300
rect 14730 -340 14770 -300
rect 14810 -340 14850 -300
rect 14890 -340 14930 -300
rect 14970 -340 15010 -300
rect 15050 -340 15090 -300
rect -1330 -4352 -1290 -4312
rect -1250 -4352 -1210 -4312
rect -1170 -4352 -1130 -4312
rect -1090 -4352 -1050 -4312
rect -1010 -4352 -970 -4312
rect -930 -4352 -890 -4312
rect -1330 -4432 -1290 -4392
rect -1250 -4432 -1210 -4392
rect -1170 -4432 -1130 -4392
rect -1090 -4432 -1050 -4392
rect -1010 -4432 -970 -4392
rect -930 -4432 -890 -4392
rect -1330 -4512 -1290 -4472
rect -1250 -4512 -1210 -4472
rect -1170 -4512 -1130 -4472
rect -1090 -4512 -1050 -4472
rect -1010 -4512 -970 -4472
rect -930 -4512 -890 -4472
rect -570 -4352 -530 -4312
rect -490 -4352 -450 -4312
rect -410 -4352 -370 -4312
rect -330 -4352 -290 -4312
rect -250 -4352 -210 -4312
rect -170 -4352 -130 -4312
rect -570 -4432 -530 -4392
rect -490 -4432 -450 -4392
rect -410 -4432 -370 -4392
rect -330 -4432 -290 -4392
rect -250 -4432 -210 -4392
rect -170 -4432 -130 -4392
rect -570 -4512 -530 -4472
rect -490 -4512 -450 -4472
rect -410 -4512 -370 -4472
rect -330 -4512 -290 -4472
rect -250 -4512 -210 -4472
rect -170 -4512 -130 -4472
rect 14910 -4352 14950 -4312
rect 14990 -4352 15030 -4312
rect 15070 -4352 15110 -4312
rect 15150 -4352 15190 -4312
rect 15230 -4352 15270 -4312
rect 15310 -4352 15350 -4312
rect 14910 -4432 14950 -4392
rect 14990 -4432 15030 -4392
rect 15070 -4432 15110 -4392
rect 15150 -4432 15190 -4392
rect 15230 -4432 15270 -4392
rect 15310 -4432 15350 -4392
rect 14910 -4512 14950 -4472
rect 14990 -4512 15030 -4472
rect 15070 -4512 15110 -4472
rect 15150 -4512 15190 -4472
rect 15230 -4512 15270 -4472
rect 15310 -4512 15350 -4472
rect 15670 -4352 15710 -4312
rect 15750 -4352 15790 -4312
rect 15830 -4352 15870 -4312
rect 15910 -4352 15950 -4312
rect 15990 -4352 16030 -4312
rect 16070 -4352 16110 -4312
rect 15670 -4432 15710 -4392
rect 15750 -4432 15790 -4392
rect 15830 -4432 15870 -4392
rect 15910 -4432 15950 -4392
rect 15990 -4432 16030 -4392
rect 16070 -4432 16110 -4392
rect 15670 -4512 15710 -4472
rect 15750 -4512 15790 -4472
rect 15830 -4512 15870 -4472
rect 15910 -4512 15950 -4472
rect 15990 -4512 16030 -4472
rect 16070 -4512 16110 -4472
rect -1700 -6530 -1640 -6490
rect -1700 -6610 -1640 -6570
rect -1700 -6690 -1640 -6650
rect -1700 -6770 -1640 -6730
rect -1700 -6850 -1640 -6810
rect -1700 -6930 -1640 -6890
rect 16420 -6530 16480 -6490
rect 16420 -6610 16480 -6570
rect 16420 -6690 16480 -6650
rect 16420 -6770 16480 -6730
rect 16420 -6850 16480 -6810
rect 16420 -6930 16480 -6890
rect -250 -9700 -210 -9660
rect -170 -9700 -130 -9660
rect -90 -9700 -50 -9660
rect -10 -9700 30 -9660
rect 70 -9700 110 -9660
rect 150 -9700 190 -9660
rect -250 -9780 -210 -9740
rect -170 -9780 -130 -9740
rect -90 -9780 -50 -9740
rect -10 -9780 30 -9740
rect 70 -9780 110 -9740
rect 150 -9780 190 -9740
rect -250 -9860 -210 -9820
rect -170 -9860 -130 -9820
rect -90 -9860 -50 -9820
rect -10 -9860 30 -9820
rect 70 -9860 110 -9820
rect 150 -9860 190 -9820
rect 7230 -9700 7270 -9660
rect 7310 -9700 7350 -9660
rect 7390 -9700 7430 -9660
rect 7470 -9700 7510 -9660
rect 7550 -9700 7590 -9660
rect 7630 -9700 7670 -9660
rect 7230 -9780 7270 -9740
rect 7310 -9780 7350 -9740
rect 7390 -9780 7430 -9740
rect 7470 -9780 7510 -9740
rect 7550 -9780 7590 -9740
rect 7630 -9780 7670 -9740
rect 7230 -9860 7270 -9820
rect 7310 -9860 7350 -9820
rect 7390 -9860 7430 -9820
rect 7470 -9860 7510 -9820
rect 7550 -9860 7590 -9820
rect 7630 -9860 7670 -9820
rect 14710 -9700 14750 -9660
rect 14790 -9700 14830 -9660
rect 14870 -9700 14910 -9660
rect 14950 -9700 14990 -9660
rect 15030 -9700 15070 -9660
rect 15110 -9700 15150 -9660
rect 14710 -9780 14750 -9740
rect 14790 -9780 14830 -9740
rect 14870 -9780 14910 -9740
rect 14950 -9780 14990 -9740
rect 15030 -9780 15070 -9740
rect 15110 -9780 15150 -9740
rect 14710 -9860 14750 -9820
rect 14790 -9860 14830 -9820
rect 14870 -9860 14910 -9820
rect 14950 -9860 14990 -9820
rect 15030 -9860 15070 -9820
rect 15110 -9860 15150 -9820
<< metal1 >>
rect 23460 7210 23940 7230
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 6920 23940 7030
rect 25860 7210 26340 7230
rect 25860 7140 25890 7210
rect 25960 7140 26000 7210
rect 26070 7140 26110 7210
rect 26180 7140 26220 7210
rect 26290 7140 26340 7210
rect 25860 7100 26340 7140
rect 25860 7030 25890 7100
rect 25960 7030 26000 7100
rect 26070 7030 26110 7100
rect 26180 7030 26220 7100
rect 26290 7030 26340 7100
rect 25860 6950 26340 7030
rect 11760 6880 13360 6900
rect 1540 6850 3140 6870
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 1540 6520 3140 6670
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6550 13360 6700
rect 21800 5670 22120 5690
rect 21800 5600 21820 5670
rect 21890 5600 21930 5670
rect 22000 5600 22120 5670
rect 21800 5560 22120 5600
rect 21800 5490 21820 5560
rect 21890 5490 21930 5560
rect 22000 5490 22120 5560
rect 21800 5450 22120 5490
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 21800 5380 21820 5450
rect 21890 5380 21930 5450
rect 22000 5380 22120 5450
rect 21800 5340 22120 5380
rect 21800 5270 21820 5340
rect 21890 5270 21930 5340
rect 22000 5270 22120 5340
rect 21800 5230 22120 5270
rect 21800 5160 21820 5230
rect 21890 5160 21930 5230
rect 22000 5160 22120 5230
rect 21800 5120 22120 5160
rect 21800 5050 21820 5120
rect 21890 5050 21930 5120
rect 22000 5050 22120 5120
rect 21800 5010 22120 5050
rect 21800 4940 21820 5010
rect 21890 4940 21930 5010
rect 22000 4940 22120 5010
rect 21800 4900 22120 4940
rect 21800 4830 21820 4900
rect 21890 4830 21930 4900
rect 22000 4830 22120 4900
rect 21800 4790 22120 4830
rect 21800 4720 21820 4790
rect 21890 4720 21930 4790
rect 22000 4720 22120 4790
rect 21800 4680 22120 4720
rect 21800 4610 21820 4680
rect 21890 4610 21930 4680
rect 22000 4610 22120 4680
rect -1740 4590 -1600 4610
rect -1740 4580 -1700 4590
rect -1740 4510 -1710 4580
rect -1740 4470 -1700 4510
rect -1740 4400 -1710 4470
rect -1740 4390 -1700 4400
rect -1640 4390 -1600 4590
rect -1740 4360 -1600 4390
rect -1740 4290 -1710 4360
rect -1640 4290 -1600 4360
rect -1740 4270 -1600 4290
rect -1740 4250 -1700 4270
rect -1740 4180 -1710 4250
rect -1740 4150 -1700 4180
rect -1640 4150 -1600 4270
rect -1740 4130 -1600 4150
rect 16380 4590 16520 4610
rect 16380 4390 16420 4590
rect 16480 4580 16520 4590
rect 16490 4510 16520 4580
rect 16480 4470 16520 4510
rect 16490 4400 16520 4470
rect 16480 4390 16520 4400
rect 16380 4360 16520 4390
rect 16380 4290 16420 4360
rect 16490 4290 16520 4360
rect 16380 4270 16520 4290
rect 16380 4150 16420 4270
rect 16480 4250 16520 4270
rect 16490 4180 16520 4250
rect 16480 4150 16520 4180
rect 16380 4130 16520 4150
rect 21800 4570 22120 4610
rect 21800 4500 21820 4570
rect 21890 4500 21930 4570
rect 22000 4500 22120 4570
rect 21800 3990 22120 4500
rect 24700 3360 25030 3380
rect 24700 3290 24720 3360
rect 24790 3290 24830 3360
rect 24900 3290 24940 3360
rect 25010 3290 25030 3360
rect 24700 3250 25030 3290
rect 24700 3180 24720 3250
rect 24790 3180 24830 3250
rect 24900 3180 24940 3250
rect 25010 3180 25030 3250
rect 24700 3140 25030 3180
rect 24700 3070 24720 3140
rect 24790 3070 24830 3140
rect 24900 3070 24940 3140
rect 25010 3070 25030 3140
rect 24700 3050 25030 3070
rect 22420 2600 22900 2670
rect 22420 2530 22470 2600
rect 22540 2530 22580 2600
rect 22650 2530 22690 2600
rect 22760 2530 22800 2600
rect 22870 2530 22900 2600
rect 22420 2490 22900 2530
rect 22420 2420 22470 2490
rect 22540 2420 22580 2490
rect 22650 2420 22690 2490
rect 22760 2420 22800 2490
rect 22870 2420 22900 2490
rect 22420 2400 22900 2420
rect 26900 2600 27380 2660
rect 26900 2530 26950 2600
rect 27020 2530 27060 2600
rect 27130 2530 27170 2600
rect 27240 2530 27280 2600
rect 27350 2530 27380 2600
rect 26900 2490 27380 2530
rect 26900 2420 26950 2490
rect 27020 2420 27060 2490
rect 27130 2420 27170 2490
rect 27240 2420 27280 2490
rect 27350 2420 27380 2490
rect 26900 2400 27380 2420
rect 14590 1160 14900 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 14900 1160
rect 14590 1050 14900 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 14900 1050
rect 14590 940 14900 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 14900 940
rect 14590 850 14900 870
rect 23460 920 23940 940
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 640 23940 740
rect 25860 920 26340 940
rect 25860 850 25890 920
rect 25960 850 26000 920
rect 26070 850 26110 920
rect 26180 850 26220 920
rect 26290 850 26340 920
rect 25860 810 26340 850
rect 25860 740 25890 810
rect 25960 740 26000 810
rect 26070 740 26110 810
rect 26180 740 26220 810
rect 26290 740 26340 810
rect 25860 650 26340 740
rect -330 -140 150 -98
rect -330 -180 -310 -140
rect -110 -180 -80 -140
rect -10 -180 10 -140
rect 130 -180 150 -140
rect -330 -210 -300 -180
rect -230 -210 -190 -180
rect -120 -210 -80 -180
rect -10 -210 30 -180
rect 100 -210 150 -180
rect -330 -220 150 -210
rect -330 -260 -310 -220
rect -270 -260 -230 -220
rect -190 -260 -150 -220
rect -110 -260 -70 -220
rect -30 -260 10 -220
rect 50 -260 90 -220
rect 130 -260 150 -220
rect -330 -270 150 -260
rect -330 -300 -300 -270
rect -230 -300 -190 -270
rect -120 -300 -80 -270
rect -10 -300 30 -270
rect 100 -300 150 -270
rect -330 -340 -310 -300
rect -110 -340 -80 -300
rect -10 -340 10 -300
rect 130 -340 150 -300
rect -330 -380 150 -340
rect 1080 -790 2680 40
rect 7150 -120 7630 -98
rect 7150 -140 7180 -120
rect 7240 -140 7280 -120
rect 7340 -140 7440 -120
rect 7500 -140 7540 -120
rect 7600 -140 7630 -120
rect 7150 -180 7170 -140
rect 7240 -180 7250 -140
rect 7370 -180 7410 -140
rect 7530 -180 7540 -140
rect 7610 -180 7630 -140
rect 7150 -210 7630 -180
rect 7150 -220 7180 -210
rect 7240 -220 7280 -210
rect 7340 -220 7440 -210
rect 7500 -220 7540 -210
rect 7600 -220 7630 -210
rect 7150 -260 7170 -220
rect 7240 -260 7250 -220
rect 7370 -260 7410 -220
rect 7530 -260 7540 -220
rect 7610 -260 7630 -220
rect 7150 -270 7180 -260
rect 7240 -270 7280 -260
rect 7340 -270 7440 -260
rect 7500 -270 7540 -260
rect 7600 -270 7630 -260
rect 7150 -300 7630 -270
rect 7150 -340 7170 -300
rect 7240 -340 7250 -300
rect 7370 -340 7410 -300
rect 7530 -340 7540 -300
rect 7610 -340 7630 -300
rect 7150 -360 7180 -340
rect 7240 -360 7280 -340
rect 7340 -360 7440 -340
rect 7500 -360 7540 -340
rect 7600 -360 7630 -340
rect 7150 -380 7630 -360
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -990 2680 -970
rect 12220 -790 13820 40
rect 14630 -140 15110 -98
rect 14630 -180 14650 -140
rect 14850 -180 14880 -140
rect 14950 -180 14970 -140
rect 15090 -180 15110 -140
rect 14630 -210 14660 -180
rect 14730 -210 14770 -180
rect 14840 -210 14880 -180
rect 14950 -210 14990 -180
rect 15060 -210 15110 -180
rect 14630 -220 15110 -210
rect 14630 -260 14650 -220
rect 14690 -260 14730 -220
rect 14770 -260 14810 -220
rect 14850 -260 14890 -220
rect 14930 -260 14970 -220
rect 15010 -260 15050 -220
rect 15090 -260 15110 -220
rect 14630 -270 15110 -260
rect 14630 -300 14660 -270
rect 14730 -300 14770 -270
rect 14840 -300 14880 -270
rect 14950 -300 14990 -270
rect 15060 -300 15110 -270
rect 14630 -340 14650 -300
rect 14850 -340 14880 -300
rect 14950 -340 14970 -300
rect 15090 -340 15110 -300
rect 14630 -380 15110 -340
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -990 13820 -970
rect 21800 -850 22060 -820
rect 21800 -920 21820 -850
rect 21890 -920 21930 -850
rect 22000 -920 22060 -850
rect 21800 -960 22060 -920
rect 21800 -1030 21820 -960
rect 21890 -1030 21930 -960
rect 22000 -1030 22060 -960
rect 21800 -1070 22060 -1030
rect 21800 -1140 21820 -1070
rect 21890 -1140 21930 -1070
rect 22000 -1140 22060 -1070
rect 21800 -1180 22060 -1140
rect 21800 -1250 21820 -1180
rect 21890 -1250 21930 -1180
rect 22000 -1250 22060 -1180
rect 21800 -1290 22060 -1250
rect 21800 -1360 21820 -1290
rect 21890 -1360 21930 -1290
rect 22000 -1360 22060 -1290
rect 21800 -1400 22060 -1360
rect 21800 -1470 21820 -1400
rect 21890 -1470 21930 -1400
rect 22000 -1470 22060 -1400
rect 21800 -1510 22060 -1470
rect 21800 -1580 21820 -1510
rect 21890 -1580 21930 -1510
rect 22000 -1580 22060 -1510
rect 21800 -1620 22060 -1580
rect 21800 -1690 21820 -1620
rect 21890 -1690 21930 -1620
rect 22000 -1690 22060 -1620
rect 21800 -1730 22060 -1690
rect 21800 -1800 21820 -1730
rect 21890 -1800 21930 -1730
rect 22000 -1800 22060 -1730
rect 21800 -1840 22060 -1800
rect 21800 -1910 21820 -1840
rect 21890 -1910 21930 -1840
rect 22000 -1910 22060 -1840
rect 21800 -1950 22060 -1910
rect 21800 -2020 21820 -1950
rect 21890 -2020 21930 -1950
rect 22000 -2020 22060 -1950
rect 21800 -2040 22060 -2020
rect 1540 -2780 3140 -2760
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -3020 3140 -2960
rect 11760 -2780 13360 -2760
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -3020 13360 -2960
rect 24720 -3050 25050 -3030
rect 24720 -3120 24740 -3050
rect 24810 -3120 24850 -3050
rect 24920 -3120 24960 -3050
rect 25030 -3120 25050 -3050
rect 24720 -3160 25050 -3120
rect 24720 -3230 24740 -3160
rect 24810 -3230 24850 -3160
rect 24920 -3230 24960 -3160
rect 25030 -3230 25050 -3160
rect 24720 -3270 25050 -3230
rect 24720 -3340 24740 -3270
rect 24810 -3340 24850 -3270
rect 24920 -3340 24960 -3270
rect 25030 -3340 25050 -3270
rect 24720 -3360 25050 -3340
rect 22420 -3690 22900 -3630
rect 22420 -3760 22470 -3690
rect 22540 -3760 22580 -3690
rect 22650 -3760 22690 -3690
rect 22760 -3760 22800 -3690
rect 22870 -3760 22900 -3690
rect 22420 -3800 22900 -3760
rect 7290 -3880 7620 -3860
rect 7290 -3950 7310 -3880
rect 7380 -3950 7420 -3880
rect 7490 -3950 7530 -3880
rect 7600 -3950 7620 -3880
rect 22420 -3870 22470 -3800
rect 22540 -3870 22580 -3800
rect 22650 -3870 22690 -3800
rect 22760 -3870 22800 -3800
rect 22870 -3870 22900 -3800
rect 22420 -3890 22900 -3870
rect 26900 -3690 27380 -3630
rect 26900 -3760 26950 -3690
rect 27020 -3760 27060 -3690
rect 27130 -3760 27170 -3690
rect 27240 -3760 27280 -3690
rect 27350 -3760 27380 -3690
rect 26900 -3800 27380 -3760
rect 26900 -3870 26950 -3800
rect 27020 -3870 27060 -3800
rect 27130 -3870 27170 -3800
rect 27240 -3870 27280 -3800
rect 27350 -3870 27380 -3800
rect 26900 -3890 27380 -3870
rect 7290 -3990 7620 -3950
rect 7290 -4060 7310 -3990
rect 7380 -4060 7420 -3990
rect 7490 -4060 7530 -3990
rect 7600 -4060 7620 -3990
rect 7290 -4100 7620 -4060
rect 7290 -4170 7310 -4100
rect 7380 -4170 7420 -4100
rect 7490 -4170 7530 -4100
rect 7600 -4170 7620 -4100
rect 7290 -4190 7620 -4170
rect -1350 -4312 -870 -4270
rect -1350 -4432 -1330 -4312
rect -1290 -4350 -1250 -4312
rect -1210 -4350 -1170 -4312
rect -1130 -4350 -1090 -4312
rect -1050 -4350 -1010 -4312
rect -970 -4350 -930 -4312
rect -1260 -4352 -1250 -4350
rect -1130 -4352 -1110 -4350
rect -1040 -4352 -1010 -4350
rect -890 -4352 -870 -4312
rect -1260 -4392 -1220 -4352
rect -1150 -4392 -1110 -4352
rect -1040 -4392 -1000 -4352
rect -930 -4392 -870 -4352
rect -1260 -4420 -1250 -4392
rect -1130 -4420 -1110 -4392
rect -1040 -4420 -1010 -4392
rect -1290 -4432 -1250 -4420
rect -1210 -4432 -1170 -4420
rect -1130 -4432 -1090 -4420
rect -1050 -4432 -1010 -4420
rect -970 -4432 -930 -4420
rect -890 -4432 -870 -4392
rect -1350 -4460 -870 -4432
rect -1350 -4530 -1330 -4460
rect -1260 -4472 -1220 -4460
rect -1150 -4472 -1110 -4460
rect -1040 -4472 -1000 -4460
rect -930 -4472 -870 -4460
rect -1260 -4512 -1250 -4472
rect -1130 -4512 -1110 -4472
rect -1040 -4512 -1010 -4472
rect -890 -4512 -870 -4472
rect -1260 -4530 -1220 -4512
rect -1150 -4530 -1110 -4512
rect -1040 -4530 -1000 -4512
rect -930 -4530 -870 -4512
rect -1350 -4552 -870 -4530
rect -588 -4290 -110 -4270
rect -588 -4312 -560 -4290
rect -490 -4312 -450 -4290
rect -380 -4312 -340 -4290
rect -270 -4312 -230 -4290
rect -160 -4312 -110 -4290
rect -588 -4352 -570 -4312
rect -370 -4352 -340 -4312
rect -270 -4352 -250 -4312
rect -130 -4352 -110 -4312
rect -588 -4360 -560 -4352
rect -490 -4360 -450 -4352
rect -380 -4360 -340 -4352
rect -270 -4360 -230 -4352
rect -160 -4360 -110 -4352
rect -588 -4392 -110 -4360
rect -588 -4432 -570 -4392
rect -530 -4400 -490 -4392
rect -450 -4400 -410 -4392
rect -370 -4400 -330 -4392
rect -290 -4400 -250 -4392
rect -210 -4400 -170 -4392
rect -370 -4432 -340 -4400
rect -270 -4432 -250 -4400
rect -130 -4432 -110 -4392
rect -588 -4470 -560 -4432
rect -490 -4470 -450 -4432
rect -380 -4470 -340 -4432
rect -270 -4470 -230 -4432
rect -160 -4470 -110 -4432
rect -588 -4472 -110 -4470
rect -588 -4512 -570 -4472
rect -530 -4512 -490 -4472
rect -450 -4512 -410 -4472
rect -370 -4512 -330 -4472
rect -290 -4512 -250 -4472
rect -210 -4512 -170 -4472
rect -130 -4512 -110 -4472
rect -588 -4552 -110 -4512
rect 14890 -4290 15368 -4270
rect 14890 -4312 14940 -4290
rect 15010 -4312 15050 -4290
rect 15120 -4312 15160 -4290
rect 15230 -4312 15270 -4290
rect 15340 -4312 15368 -4290
rect 14890 -4352 14910 -4312
rect 15030 -4352 15050 -4312
rect 15120 -4352 15150 -4312
rect 15350 -4352 15368 -4312
rect 14890 -4360 14940 -4352
rect 15010 -4360 15050 -4352
rect 15120 -4360 15160 -4352
rect 15230 -4360 15270 -4352
rect 15340 -4360 15368 -4352
rect 14890 -4392 15368 -4360
rect 14890 -4432 14910 -4392
rect 14950 -4400 14990 -4392
rect 15030 -4400 15070 -4392
rect 15110 -4400 15150 -4392
rect 15190 -4400 15230 -4392
rect 15030 -4432 15050 -4400
rect 15120 -4432 15150 -4400
rect 15270 -4400 15310 -4392
rect 15350 -4432 15368 -4392
rect 14890 -4470 14940 -4432
rect 15010 -4470 15050 -4432
rect 15120 -4470 15160 -4432
rect 15230 -4470 15270 -4432
rect 15340 -4470 15368 -4432
rect 14890 -4472 15368 -4470
rect 14890 -4512 14910 -4472
rect 14950 -4512 14990 -4472
rect 15030 -4512 15070 -4472
rect 15110 -4512 15150 -4472
rect 15190 -4512 15230 -4472
rect 15270 -4512 15310 -4472
rect 15350 -4512 15368 -4472
rect 14890 -4552 15368 -4512
rect 15650 -4312 16130 -4270
rect 15650 -4352 15670 -4312
rect 15710 -4350 15750 -4312
rect 15790 -4350 15830 -4312
rect 15870 -4350 15910 -4312
rect 15950 -4350 15990 -4312
rect 16030 -4350 16070 -4312
rect 15790 -4352 15820 -4350
rect 15890 -4352 15910 -4350
rect 16030 -4352 16040 -4350
rect 15650 -4392 15710 -4352
rect 15780 -4392 15820 -4352
rect 15890 -4392 15930 -4352
rect 16000 -4392 16040 -4352
rect 15650 -4432 15670 -4392
rect 15790 -4420 15820 -4392
rect 15890 -4420 15910 -4392
rect 16030 -4420 16040 -4392
rect 15710 -4432 15750 -4420
rect 15790 -4432 15830 -4420
rect 15870 -4432 15910 -4420
rect 15950 -4432 15990 -4420
rect 16030 -4432 16070 -4420
rect 16110 -4432 16130 -4312
rect 15650 -4460 16130 -4432
rect 15650 -4472 15710 -4460
rect 15780 -4472 15820 -4460
rect 15890 -4472 15930 -4460
rect 16000 -4472 16040 -4460
rect 15650 -4512 15670 -4472
rect 15790 -4512 15820 -4472
rect 15890 -4512 15910 -4472
rect 16030 -4512 16040 -4472
rect 15650 -4530 15710 -4512
rect 15780 -4530 15820 -4512
rect 15890 -4530 15930 -4512
rect 16000 -4530 16040 -4512
rect 16110 -4530 16130 -4460
rect 15650 -4552 16130 -4530
rect 7570 -6460 7870 -6420
rect -1740 -6490 -1600 -6470
rect -1740 -6520 -1700 -6490
rect -1740 -6590 -1710 -6520
rect -1740 -6610 -1700 -6590
rect -1640 -6610 -1600 -6490
rect 7570 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 7870 -6460
rect 7570 -6560 7870 -6520
rect -1740 -6630 -1600 -6610
rect 7570 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 7870 -6560
rect -1740 -6700 -1710 -6630
rect -1640 -6700 -1600 -6630
rect 7570 -6660 7870 -6620
rect -1740 -6730 -1600 -6700
rect 7570 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 7870 -6660
rect 16380 -6490 16520 -6470
rect 16380 -6610 16420 -6490
rect 16480 -6520 16520 -6490
rect 16490 -6590 16520 -6520
rect 16480 -6610 16520 -6590
rect 16380 -6630 16520 -6610
rect -1740 -6740 -1700 -6730
rect -1740 -6810 -1710 -6740
rect -1740 -6850 -1700 -6810
rect -1740 -6920 -1710 -6850
rect -1740 -6930 -1700 -6920
rect -1640 -6930 -1600 -6730
rect 7570 -6760 7870 -6720
rect 16380 -6700 16420 -6630
rect 16490 -6700 16520 -6630
rect 16380 -6730 16520 -6700
rect 7570 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 7870 -6760
rect 7570 -6850 7870 -6820
rect 16380 -6930 16420 -6730
rect 16480 -6740 16520 -6730
rect 16490 -6810 16520 -6740
rect 16480 -6850 16520 -6810
rect 16490 -6920 16520 -6850
rect 16480 -6930 16520 -6920
rect -1740 -6950 -1600 -6930
rect 16380 -6950 16520 -6930
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 21610 -8360 22540 -8330
rect 21610 -8430 21630 -8360
rect 21700 -8430 21730 -8360
rect 21800 -8430 21830 -8360
rect 21900 -8430 22540 -8360
rect 21610 -8460 22540 -8430
rect 21610 -8530 21630 -8460
rect 21700 -8530 21730 -8460
rect 21800 -8530 21830 -8460
rect 21900 -8530 22540 -8460
rect 21610 -8560 22540 -8530
rect 21610 -8630 21630 -8560
rect 21700 -8630 21730 -8560
rect 21800 -8630 21830 -8560
rect 21900 -8630 22540 -8560
rect 21610 -8650 22540 -8630
rect 22630 -9010 22950 -8980
rect 22630 -9080 22650 -9010
rect 22720 -9080 22750 -9010
rect 22820 -9080 22850 -9010
rect 22920 -9080 22950 -9010
rect 22630 -9110 22950 -9080
rect 22630 -9180 22650 -9110
rect 22720 -9180 22750 -9110
rect 22820 -9180 22850 -9110
rect 22920 -9180 22950 -9110
rect 22630 -9210 22950 -9180
rect 22630 -9280 22650 -9210
rect 22720 -9280 22750 -9210
rect 22820 -9280 22850 -9210
rect 22920 -9280 22950 -9210
rect 22630 -9300 22950 -9280
rect -270 -9660 210 -9618
rect -270 -9700 -250 -9660
rect -50 -9700 -20 -9660
rect 50 -9700 70 -9660
rect 190 -9700 210 -9660
rect -270 -9730 -240 -9700
rect -170 -9730 -130 -9700
rect -60 -9730 -20 -9700
rect 50 -9730 90 -9700
rect 160 -9730 210 -9700
rect -270 -9740 210 -9730
rect -270 -9780 -250 -9740
rect -210 -9780 -170 -9740
rect -130 -9780 -90 -9740
rect -50 -9780 -10 -9740
rect 30 -9780 70 -9740
rect 110 -9780 150 -9740
rect 190 -9780 210 -9740
rect -270 -9790 210 -9780
rect -270 -9820 -240 -9790
rect -170 -9820 -130 -9790
rect -60 -9820 -20 -9790
rect 50 -9820 90 -9790
rect 160 -9820 210 -9790
rect -270 -9860 -250 -9820
rect -50 -9860 -20 -9820
rect 50 -9860 70 -9820
rect 190 -9860 210 -9820
rect -270 -9900 210 -9860
rect 1080 -10340 2680 -9500
rect 7210 -9640 7690 -9618
rect 7210 -9660 7240 -9640
rect 7300 -9660 7340 -9640
rect 7400 -9660 7500 -9640
rect 7560 -9660 7600 -9640
rect 7660 -9660 7690 -9640
rect 7210 -9700 7230 -9660
rect 7300 -9700 7310 -9660
rect 7430 -9700 7470 -9660
rect 7590 -9700 7600 -9660
rect 7670 -9700 7690 -9660
rect 7210 -9730 7690 -9700
rect 7210 -9740 7240 -9730
rect 7300 -9740 7340 -9730
rect 7400 -9740 7500 -9730
rect 7560 -9740 7600 -9730
rect 7660 -9740 7690 -9730
rect 7210 -9780 7230 -9740
rect 7300 -9780 7310 -9740
rect 7430 -9780 7470 -9740
rect 7590 -9780 7600 -9740
rect 7670 -9780 7690 -9740
rect 7210 -9790 7240 -9780
rect 7300 -9790 7340 -9780
rect 7400 -9790 7500 -9780
rect 7560 -9790 7600 -9780
rect 7660 -9790 7690 -9780
rect 7210 -9820 7690 -9790
rect 7210 -9860 7230 -9820
rect 7300 -9860 7310 -9820
rect 7430 -9860 7470 -9820
rect 7590 -9860 7600 -9820
rect 7670 -9860 7690 -9820
rect 7210 -9880 7240 -9860
rect 7300 -9880 7340 -9860
rect 7400 -9880 7500 -9860
rect 7560 -9880 7600 -9860
rect 7660 -9880 7690 -9860
rect 7210 -9900 7690 -9880
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10540 2680 -10520
rect 12220 -10370 13820 -9520
rect 14690 -9660 15170 -9618
rect 14690 -9700 14710 -9660
rect 14910 -9700 14940 -9660
rect 15010 -9700 15030 -9660
rect 15150 -9700 15170 -9660
rect 14690 -9730 14720 -9700
rect 14790 -9730 14830 -9700
rect 14900 -9730 14940 -9700
rect 15010 -9730 15050 -9700
rect 15120 -9730 15170 -9700
rect 14690 -9740 15170 -9730
rect 14690 -9780 14710 -9740
rect 14750 -9780 14790 -9740
rect 14830 -9780 14870 -9740
rect 14910 -9780 14950 -9740
rect 14990 -9780 15030 -9740
rect 15070 -9780 15110 -9740
rect 15150 -9780 15170 -9740
rect 14690 -9790 15170 -9780
rect 14690 -9820 14720 -9790
rect 14790 -9820 14830 -9790
rect 14900 -9820 14940 -9790
rect 15010 -9820 15050 -9790
rect 15120 -9820 15170 -9790
rect 14690 -9860 14710 -9820
rect 14910 -9860 14940 -9820
rect 15010 -9860 15030 -9820
rect 15150 -9860 15170 -9820
rect 14690 -9900 15170 -9860
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10570 13820 -10550
rect 2210 -12300 3810 -12280
rect 2210 -12370 2240 -12300
rect 2310 -12370 2350 -12300
rect 2420 -12370 2460 -12300
rect 2530 -12370 2570 -12300
rect 2640 -12370 2680 -12300
rect 2750 -12370 2790 -12300
rect 2860 -12370 2900 -12300
rect 2970 -12370 3010 -12300
rect 3080 -12370 3120 -12300
rect 3190 -12370 3230 -12300
rect 3300 -12370 3340 -12300
rect 3410 -12370 3450 -12300
rect 3520 -12370 3560 -12300
rect 3630 -12370 3670 -12300
rect 3740 -12370 3810 -12300
rect 2210 -12410 3810 -12370
rect 2210 -12480 2240 -12410
rect 2310 -12480 2350 -12410
rect 2420 -12480 2460 -12410
rect 2530 -12480 2570 -12410
rect 2640 -12480 2680 -12410
rect 2750 -12480 2790 -12410
rect 2860 -12480 2900 -12410
rect 2970 -12480 3010 -12410
rect 3080 -12480 3120 -12410
rect 3190 -12480 3230 -12410
rect 3300 -12480 3340 -12410
rect 3410 -12480 3450 -12410
rect 3520 -12480 3560 -12410
rect 3630 -12480 3670 -12410
rect 3740 -12480 3810 -12410
rect 2210 -12550 3810 -12480
rect 11090 -12300 12690 -12280
rect 11090 -12370 11120 -12300
rect 11190 -12370 11230 -12300
rect 11300 -12370 11340 -12300
rect 11410 -12370 11450 -12300
rect 11520 -12370 11560 -12300
rect 11630 -12370 11670 -12300
rect 11740 -12370 11780 -12300
rect 11850 -12370 11890 -12300
rect 11960 -12370 12000 -12300
rect 12070 -12370 12110 -12300
rect 12180 -12370 12220 -12300
rect 12290 -12370 12330 -12300
rect 12400 -12370 12440 -12300
rect 12510 -12370 12550 -12300
rect 12620 -12370 12690 -12300
rect 11090 -12410 12690 -12370
rect 11090 -12480 11120 -12410
rect 11190 -12480 11230 -12410
rect 11300 -12480 11340 -12410
rect 11410 -12480 11450 -12410
rect 11520 -12480 11560 -12410
rect 11630 -12480 11670 -12410
rect 11740 -12480 11780 -12410
rect 11850 -12480 11890 -12410
rect 11960 -12480 12000 -12410
rect 12070 -12480 12110 -12410
rect 12180 -12480 12220 -12410
rect 12290 -12480 12330 -12410
rect 12400 -12480 12440 -12410
rect 12510 -12480 12550 -12410
rect 12620 -12480 12690 -12410
rect 11090 -12550 12690 -12480
rect 21610 -14020 22820 -13990
rect 21610 -14090 21630 -14020
rect 21700 -14090 21730 -14020
rect 21800 -14090 21830 -14020
rect 21900 -14090 22820 -14020
rect 21610 -14120 22820 -14090
rect 21610 -14190 21630 -14120
rect 21700 -14190 21730 -14120
rect 21800 -14190 21830 -14120
rect 21900 -14190 22820 -14120
rect 21610 -14220 22820 -14190
rect 21610 -14290 21630 -14220
rect 21700 -14290 21730 -14220
rect 21800 -14290 21830 -14220
rect 21900 -14290 22820 -14220
rect 21610 -14310 22820 -14290
rect 22900 -14870 23220 -14840
rect 22900 -14940 22920 -14870
rect 22990 -14940 23020 -14870
rect 23090 -14940 23120 -14870
rect 23190 -14940 23220 -14870
rect 22900 -14970 23220 -14940
rect 22900 -15040 22920 -14970
rect 22990 -15040 23020 -14970
rect 23090 -15040 23120 -14970
rect 23190 -15040 23220 -14970
rect 22900 -15070 23220 -15040
rect 22900 -15140 22920 -15070
rect 22990 -15140 23020 -15070
rect 23090 -15140 23120 -15070
rect 23190 -15140 23220 -15070
rect 22900 -15160 23220 -15140
rect 7210 -17600 7650 -17580
rect 7210 -17670 7230 -17600
rect 7300 -17670 7340 -17600
rect 7410 -17670 7450 -17600
rect 7520 -17670 7560 -17600
rect 7630 -17670 7650 -17600
rect 7210 -17710 7650 -17670
rect 7210 -17780 7230 -17710
rect 7300 -17780 7340 -17710
rect 7410 -17780 7450 -17710
rect 7520 -17780 7560 -17710
rect 7630 -17780 7650 -17710
rect 7210 -17820 7650 -17780
rect 7210 -17890 7230 -17820
rect 7300 -17890 7340 -17820
rect 7410 -17890 7450 -17820
rect 7520 -17890 7560 -17820
rect 7630 -17890 7650 -17820
rect 7210 -17930 7650 -17890
rect 7210 -18000 7230 -17930
rect 7300 -18000 7340 -17930
rect 7410 -18000 7450 -17930
rect 7520 -18000 7560 -17930
rect 7630 -18000 7650 -17930
rect 7210 -18020 7650 -18000
rect 21610 -20100 22620 -20070
rect 21610 -20170 21630 -20100
rect 21700 -20170 21730 -20100
rect 21800 -20170 21830 -20100
rect 21900 -20170 22620 -20100
rect 21610 -20200 22620 -20170
rect 21610 -20270 21630 -20200
rect 21700 -20270 21730 -20200
rect 21800 -20270 21830 -20200
rect 21900 -20270 22620 -20200
rect 21610 -20300 22620 -20270
rect 21610 -20370 21630 -20300
rect 21700 -20370 21730 -20300
rect 21800 -20370 21830 -20300
rect 21900 -20370 22620 -20300
rect 21610 -20390 22620 -20370
rect 22680 -20730 23000 -20700
rect 22680 -20800 22700 -20730
rect 22770 -20800 22800 -20730
rect 22870 -20800 22900 -20730
rect 22970 -20800 23000 -20730
rect 22680 -20830 23000 -20800
rect 22680 -20900 22700 -20830
rect 22770 -20900 22800 -20830
rect 22870 -20900 22900 -20830
rect 22970 -20900 23000 -20830
rect 22680 -20930 23000 -20900
rect 22680 -21000 22700 -20930
rect 22770 -21000 22800 -20930
rect 22870 -21000 22900 -20930
rect 22970 -21000 23000 -20930
rect 22680 -21020 23000 -21000
rect 2210 -22660 3810 -22590
rect 2210 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3160 -22660
rect 3230 -22730 3270 -22660
rect 3340 -22730 3380 -22660
rect 3450 -22730 3490 -22660
rect 3560 -22730 3600 -22660
rect 3670 -22730 3710 -22660
rect 3780 -22730 3810 -22660
rect 2210 -22770 3810 -22730
rect 2210 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3160 -22770
rect 3230 -22840 3270 -22770
rect 3340 -22840 3380 -22770
rect 3450 -22840 3490 -22770
rect 3560 -22840 3600 -22770
rect 3670 -22840 3710 -22770
rect 3780 -22840 3810 -22770
rect 2210 -22860 3810 -22840
rect 11090 -22660 12690 -22590
rect 11090 -22730 11160 -22660
rect 11230 -22730 11270 -22660
rect 11340 -22730 11380 -22660
rect 11450 -22730 11490 -22660
rect 11560 -22730 11600 -22660
rect 11670 -22730 11710 -22660
rect 11780 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12690 -22660
rect 11090 -22770 12690 -22730
rect 11090 -22840 11160 -22770
rect 11230 -22840 11270 -22770
rect 11340 -22840 11380 -22770
rect 11450 -22840 11490 -22770
rect 11560 -22840 11600 -22770
rect 11670 -22840 11710 -22770
rect 11780 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12690 -22770
rect 11090 -22860 12690 -22840
<< via1 >>
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 25890 7140 25960 7210
rect 26000 7140 26070 7210
rect 26110 7140 26180 7210
rect 26220 7140 26290 7210
rect 25890 7030 25960 7100
rect 26000 7030 26070 7100
rect 26110 7030 26180 7100
rect 26220 7030 26290 7100
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 7380 6230 7440 6290
rect 7480 6230 7540 6290
rect 22780 6210 22850 6280
rect 22890 6210 22960 6280
rect 23000 6210 23070 6280
rect 23110 6210 23180 6280
rect 7380 6080 7440 6190
rect 7480 6080 7540 6190
rect 22780 6100 22850 6170
rect 22890 6100 22960 6170
rect 23000 6100 23070 6170
rect 23110 6100 23180 6170
rect 7380 5980 7440 6040
rect 7480 5980 7540 6040
rect 22780 5990 22850 6060
rect 22890 5990 22960 6060
rect 23000 5990 23070 6060
rect 23110 5990 23180 6060
rect 21820 5600 21890 5670
rect 21930 5600 22000 5670
rect 21820 5490 21890 5560
rect 21930 5490 22000 5560
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect 21820 5380 21890 5450
rect 21930 5380 22000 5450
rect 21820 5270 21890 5340
rect 21930 5270 22000 5340
rect 21820 5160 21890 5230
rect 21930 5160 22000 5230
rect 21820 5050 21890 5120
rect 21930 5050 22000 5120
rect 21820 4940 21890 5010
rect 21930 4940 22000 5010
rect 21820 4830 21890 4900
rect 21930 4830 22000 4900
rect 27710 4810 27770 4870
rect 27810 4810 27870 4870
rect 27910 4810 27970 4870
rect 21820 4720 21890 4790
rect 21930 4720 22000 4790
rect 27710 4710 27770 4770
rect 27810 4710 27870 4770
rect 27910 4710 27970 4770
rect 21820 4610 21890 4680
rect 21930 4610 22000 4680
rect 27710 4610 27770 4670
rect 27810 4610 27870 4670
rect 27910 4610 27970 4670
rect -1710 4550 -1700 4580
rect -1700 4550 -1640 4580
rect -1710 4510 -1640 4550
rect -1710 4430 -1640 4470
rect -1710 4400 -1700 4430
rect -1700 4400 -1640 4430
rect -1710 4350 -1640 4360
rect -1710 4310 -1700 4350
rect -1700 4310 -1640 4350
rect -1710 4290 -1640 4310
rect -1710 4230 -1700 4250
rect -1700 4230 -1640 4250
rect -1710 4190 -1640 4230
rect -1710 4180 -1700 4190
rect -1700 4180 -1640 4190
rect 16420 4550 16480 4580
rect 16480 4550 16490 4580
rect 16420 4510 16490 4550
rect 16420 4430 16490 4470
rect 16420 4400 16480 4430
rect 16480 4400 16490 4430
rect 16420 4350 16490 4360
rect 16420 4310 16480 4350
rect 16480 4310 16490 4350
rect 16420 4290 16490 4310
rect 16420 4230 16480 4250
rect 16480 4230 16490 4250
rect 16420 4190 16490 4230
rect 16420 4180 16480 4190
rect 16480 4180 16490 4190
rect 21820 4500 21890 4570
rect 21930 4500 22000 4570
rect 27710 4510 27770 4570
rect 27810 4510 27870 4570
rect 27910 4510 27970 4570
rect 27710 4410 27770 4470
rect 27810 4410 27870 4470
rect 27910 4410 27970 4470
rect 27710 4310 27770 4370
rect 27810 4310 27870 4370
rect 27910 4310 27970 4370
rect 27710 4210 27770 4270
rect 27810 4210 27870 4270
rect 27910 4210 27970 4270
rect 27710 4110 27770 4170
rect 27810 4110 27870 4170
rect 27910 4110 27970 4170
rect 27710 4010 27770 4070
rect 27810 4010 27870 4070
rect 27910 4010 27970 4070
rect 24720 3290 24790 3360
rect 24830 3290 24900 3360
rect 24940 3290 25010 3360
rect 7050 3180 7110 3240
rect 7150 3180 7210 3240
rect 7250 3180 7310 3240
rect 7590 3180 7650 3240
rect 7690 3180 7750 3240
rect 7790 3180 7850 3240
rect 24720 3180 24790 3250
rect 24830 3180 24900 3250
rect 24940 3180 25010 3250
rect 7050 3080 7110 3140
rect 7150 3080 7210 3140
rect 7250 3080 7310 3140
rect 7590 3080 7650 3140
rect 7690 3080 7750 3140
rect 7790 3080 7850 3140
rect 24720 3070 24790 3140
rect 24830 3070 24900 3140
rect 24940 3070 25010 3140
rect 7050 2980 7110 3040
rect 7150 2980 7210 3040
rect 7250 2980 7310 3040
rect 7590 2980 7650 3040
rect 7690 2980 7750 3040
rect 7790 2980 7850 3040
rect 4770 2830 4830 2890
rect 4870 2830 4930 2890
rect 4970 2830 5030 2890
rect 9870 2830 9930 2890
rect 9970 2830 10030 2890
rect 10070 2830 10130 2890
rect 4770 2730 4830 2790
rect 4870 2730 4930 2790
rect 4970 2730 5030 2790
rect 9870 2730 9930 2790
rect 9970 2730 10030 2790
rect 10070 2730 10130 2790
rect 4770 2630 4830 2690
rect 4870 2630 4930 2690
rect 4970 2630 5030 2690
rect 9870 2630 9930 2690
rect 9970 2630 10030 2690
rect 10070 2630 10130 2690
rect 22470 2530 22540 2600
rect 22580 2530 22650 2600
rect 22690 2530 22760 2600
rect 22800 2530 22870 2600
rect 22470 2420 22540 2490
rect 22580 2420 22650 2490
rect 22690 2420 22760 2490
rect 22800 2420 22870 2490
rect 26950 2530 27020 2600
rect 27060 2530 27130 2600
rect 27170 2530 27240 2600
rect 27280 2530 27350 2600
rect 26950 2420 27020 2490
rect 27060 2420 27130 2490
rect 27170 2420 27240 2490
rect 27280 2420 27350 2490
rect 14600 1090 14670 1160
rect 14700 1090 14770 1160
rect 14810 1090 14880 1160
rect 14600 980 14670 1050
rect 14700 980 14770 1050
rect 14810 980 14880 1050
rect 14600 870 14670 940
rect 14700 870 14770 940
rect 14810 870 14880 940
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect 25890 850 25960 920
rect 26000 850 26070 920
rect 26110 850 26180 920
rect 26220 850 26290 920
rect 25890 740 25960 810
rect 26000 740 26070 810
rect 26110 740 26180 810
rect 26220 740 26290 810
rect -300 -180 -270 -140
rect -270 -180 -230 -140
rect -190 -180 -150 -140
rect -150 -180 -120 -140
rect -80 -180 -70 -140
rect -70 -180 -30 -140
rect -30 -180 -10 -140
rect 30 -180 50 -140
rect 50 -180 90 -140
rect 90 -180 100 -140
rect -300 -210 -230 -180
rect -190 -210 -120 -180
rect -80 -210 -10 -180
rect 30 -210 100 -180
rect -300 -300 -230 -270
rect -190 -300 -120 -270
rect -80 -300 -10 -270
rect 30 -300 100 -270
rect -300 -340 -270 -300
rect -270 -340 -230 -300
rect -190 -340 -150 -300
rect -150 -340 -120 -300
rect -80 -340 -70 -300
rect -70 -340 -30 -300
rect -30 -340 -10 -300
rect 30 -340 50 -300
rect 50 -340 90 -300
rect 90 -340 100 -300
rect 7180 -140 7240 -120
rect 7280 -140 7340 -120
rect 7440 -140 7500 -120
rect 7540 -140 7600 -120
rect 7180 -180 7210 -140
rect 7210 -180 7240 -140
rect 7280 -180 7290 -140
rect 7290 -180 7330 -140
rect 7330 -180 7340 -140
rect 7440 -180 7450 -140
rect 7450 -180 7490 -140
rect 7490 -180 7500 -140
rect 7540 -180 7570 -140
rect 7570 -180 7600 -140
rect 7180 -220 7240 -210
rect 7280 -220 7340 -210
rect 7440 -220 7500 -210
rect 7540 -220 7600 -210
rect 7180 -260 7210 -220
rect 7210 -260 7240 -220
rect 7280 -260 7290 -220
rect 7290 -260 7330 -220
rect 7330 -260 7340 -220
rect 7440 -260 7450 -220
rect 7450 -260 7490 -220
rect 7490 -260 7500 -220
rect 7540 -260 7570 -220
rect 7570 -260 7600 -220
rect 7180 -270 7240 -260
rect 7280 -270 7340 -260
rect 7440 -270 7500 -260
rect 7540 -270 7600 -260
rect 7180 -340 7210 -300
rect 7210 -340 7240 -300
rect 7280 -340 7290 -300
rect 7290 -340 7330 -300
rect 7330 -340 7340 -300
rect 7440 -340 7450 -300
rect 7450 -340 7490 -300
rect 7490 -340 7500 -300
rect 7540 -340 7570 -300
rect 7570 -340 7600 -300
rect 7180 -360 7240 -340
rect 7280 -360 7340 -340
rect 7440 -360 7500 -340
rect 7540 -360 7600 -340
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 22780 -90 22850 -20
rect 22890 -90 22960 -20
rect 23000 -90 23070 -20
rect 23110 -90 23180 -20
rect 14660 -180 14690 -140
rect 14690 -180 14730 -140
rect 14770 -180 14810 -140
rect 14810 -180 14840 -140
rect 14880 -180 14890 -140
rect 14890 -180 14930 -140
rect 14930 -180 14950 -140
rect 14990 -180 15010 -140
rect 15010 -180 15050 -140
rect 15050 -180 15060 -140
rect 14660 -210 14730 -180
rect 14770 -210 14840 -180
rect 14880 -210 14950 -180
rect 14990 -210 15060 -180
rect 22780 -200 22850 -130
rect 22890 -200 22960 -130
rect 23000 -200 23070 -130
rect 23110 -200 23180 -130
rect 14660 -300 14730 -270
rect 14770 -300 14840 -270
rect 14880 -300 14950 -270
rect 14990 -300 15060 -270
rect 14660 -340 14690 -300
rect 14690 -340 14730 -300
rect 14770 -340 14810 -300
rect 14810 -340 14840 -300
rect 14880 -340 14890 -300
rect 14890 -340 14930 -300
rect 14930 -340 14950 -300
rect 14990 -340 15010 -300
rect 15010 -340 15050 -300
rect 15050 -340 15060 -300
rect 22780 -310 22850 -240
rect 22890 -310 22960 -240
rect 23000 -310 23070 -240
rect 23110 -310 23180 -240
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 21820 -920 21890 -850
rect 21930 -920 22000 -850
rect 21820 -1030 21890 -960
rect 21930 -1030 22000 -960
rect 21820 -1140 21890 -1070
rect 21930 -1140 22000 -1070
rect 21820 -1250 21890 -1180
rect 21930 -1250 22000 -1180
rect 21820 -1360 21890 -1290
rect 21930 -1360 22000 -1290
rect 21820 -1470 21890 -1400
rect 21930 -1470 22000 -1400
rect 27710 -1490 27770 -1430
rect 27810 -1490 27870 -1430
rect 27910 -1490 27970 -1430
rect 21820 -1580 21890 -1510
rect 21930 -1580 22000 -1510
rect 27710 -1590 27770 -1530
rect 27810 -1590 27870 -1530
rect 27910 -1590 27970 -1530
rect 21820 -1690 21890 -1620
rect 21930 -1690 22000 -1620
rect 27710 -1690 27770 -1630
rect 27810 -1690 27870 -1630
rect 27910 -1690 27970 -1630
rect 21820 -1800 21890 -1730
rect 21930 -1800 22000 -1730
rect 27710 -1790 27770 -1730
rect 27810 -1790 27870 -1730
rect 27910 -1790 27970 -1730
rect 21820 -1910 21890 -1840
rect 21930 -1910 22000 -1840
rect 27710 -1890 27770 -1830
rect 27810 -1890 27870 -1830
rect 27910 -1890 27970 -1830
rect 21820 -2020 21890 -1950
rect 21930 -2020 22000 -1950
rect 27710 -1990 27770 -1930
rect 27810 -1990 27870 -1930
rect 27910 -1990 27970 -1930
rect 27710 -2090 27770 -2030
rect 27810 -2090 27870 -2030
rect 27910 -2090 27970 -2030
rect 27710 -2190 27770 -2130
rect 27810 -2190 27870 -2130
rect 27910 -2190 27970 -2130
rect 27710 -2290 27770 -2230
rect 27810 -2290 27870 -2230
rect 27910 -2290 27970 -2230
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 24740 -3120 24810 -3050
rect 24850 -3120 24920 -3050
rect 24960 -3120 25030 -3050
rect 24740 -3230 24810 -3160
rect 24850 -3230 24920 -3160
rect 24960 -3230 25030 -3160
rect 24740 -3340 24810 -3270
rect 24850 -3340 24920 -3270
rect 24960 -3340 25030 -3270
rect 7380 -3400 7440 -3340
rect 7480 -3400 7540 -3340
rect 7380 -3550 7440 -3440
rect 7480 -3550 7540 -3440
rect 7380 -3650 7440 -3590
rect 7480 -3650 7540 -3590
rect 22470 -3760 22540 -3690
rect 22580 -3760 22650 -3690
rect 22690 -3760 22760 -3690
rect 22800 -3760 22870 -3690
rect 7310 -3950 7380 -3880
rect 7420 -3950 7490 -3880
rect 7530 -3950 7600 -3880
rect 22470 -3870 22540 -3800
rect 22580 -3870 22650 -3800
rect 22690 -3870 22760 -3800
rect 22800 -3870 22870 -3800
rect 26950 -3760 27020 -3690
rect 27060 -3760 27130 -3690
rect 27170 -3760 27240 -3690
rect 27280 -3760 27350 -3690
rect 26950 -3870 27020 -3800
rect 27060 -3870 27130 -3800
rect 27170 -3870 27240 -3800
rect 27280 -3870 27350 -3800
rect 7310 -4060 7380 -3990
rect 7420 -4060 7490 -3990
rect 7530 -4060 7600 -3990
rect 7310 -4170 7380 -4100
rect 7420 -4170 7490 -4100
rect 7530 -4170 7600 -4100
rect -1330 -4352 -1290 -4350
rect -1290 -4352 -1260 -4350
rect -1220 -4352 -1210 -4350
rect -1210 -4352 -1170 -4350
rect -1170 -4352 -1150 -4350
rect -1110 -4352 -1090 -4350
rect -1090 -4352 -1050 -4350
rect -1050 -4352 -1040 -4350
rect -1000 -4352 -970 -4350
rect -970 -4352 -930 -4350
rect -1330 -4392 -1260 -4352
rect -1220 -4392 -1150 -4352
rect -1110 -4392 -1040 -4352
rect -1000 -4392 -930 -4352
rect -1330 -4420 -1290 -4392
rect -1290 -4420 -1260 -4392
rect -1220 -4420 -1210 -4392
rect -1210 -4420 -1170 -4392
rect -1170 -4420 -1150 -4392
rect -1110 -4420 -1090 -4392
rect -1090 -4420 -1050 -4392
rect -1050 -4420 -1040 -4392
rect -1000 -4420 -970 -4392
rect -970 -4420 -930 -4392
rect -1330 -4472 -1260 -4460
rect -1220 -4472 -1150 -4460
rect -1110 -4472 -1040 -4460
rect -1000 -4472 -930 -4460
rect -1330 -4512 -1290 -4472
rect -1290 -4512 -1260 -4472
rect -1220 -4512 -1210 -4472
rect -1210 -4512 -1170 -4472
rect -1170 -4512 -1150 -4472
rect -1110 -4512 -1090 -4472
rect -1090 -4512 -1050 -4472
rect -1050 -4512 -1040 -4472
rect -1000 -4512 -970 -4472
rect -970 -4512 -930 -4472
rect -1330 -4530 -1260 -4512
rect -1220 -4530 -1150 -4512
rect -1110 -4530 -1040 -4512
rect -1000 -4530 -930 -4512
rect -560 -4312 -490 -4290
rect -450 -4312 -380 -4290
rect -340 -4312 -270 -4290
rect -230 -4312 -160 -4290
rect -560 -4352 -530 -4312
rect -530 -4352 -490 -4312
rect -450 -4352 -410 -4312
rect -410 -4352 -380 -4312
rect -340 -4352 -330 -4312
rect -330 -4352 -290 -4312
rect -290 -4352 -270 -4312
rect -230 -4352 -210 -4312
rect -210 -4352 -170 -4312
rect -170 -4352 -160 -4312
rect -560 -4360 -490 -4352
rect -450 -4360 -380 -4352
rect -340 -4360 -270 -4352
rect -230 -4360 -160 -4352
rect -560 -4432 -530 -4400
rect -530 -4432 -490 -4400
rect -450 -4432 -410 -4400
rect -410 -4432 -380 -4400
rect -340 -4432 -330 -4400
rect -330 -4432 -290 -4400
rect -290 -4432 -270 -4400
rect -230 -4432 -210 -4400
rect -210 -4432 -170 -4400
rect -170 -4432 -160 -4400
rect -560 -4470 -490 -4432
rect -450 -4470 -380 -4432
rect -340 -4470 -270 -4432
rect -230 -4470 -160 -4432
rect 14940 -4312 15010 -4290
rect 15050 -4312 15120 -4290
rect 15160 -4312 15230 -4290
rect 15270 -4312 15340 -4290
rect 14940 -4352 14950 -4312
rect 14950 -4352 14990 -4312
rect 14990 -4352 15010 -4312
rect 15050 -4352 15070 -4312
rect 15070 -4352 15110 -4312
rect 15110 -4352 15120 -4312
rect 15160 -4352 15190 -4312
rect 15190 -4352 15230 -4312
rect 15270 -4352 15310 -4312
rect 15310 -4352 15340 -4312
rect 14940 -4360 15010 -4352
rect 15050 -4360 15120 -4352
rect 15160 -4360 15230 -4352
rect 15270 -4360 15340 -4352
rect 14940 -4432 14950 -4400
rect 14950 -4432 14990 -4400
rect 14990 -4432 15010 -4400
rect 15050 -4432 15070 -4400
rect 15070 -4432 15110 -4400
rect 15110 -4432 15120 -4400
rect 15160 -4432 15190 -4400
rect 15190 -4432 15230 -4400
rect 15270 -4432 15310 -4400
rect 15310 -4432 15340 -4400
rect 14940 -4470 15010 -4432
rect 15050 -4470 15120 -4432
rect 15160 -4470 15230 -4432
rect 15270 -4470 15340 -4432
rect 15710 -4352 15750 -4350
rect 15750 -4352 15780 -4350
rect 15820 -4352 15830 -4350
rect 15830 -4352 15870 -4350
rect 15870 -4352 15890 -4350
rect 15930 -4352 15950 -4350
rect 15950 -4352 15990 -4350
rect 15990 -4352 16000 -4350
rect 16040 -4352 16070 -4350
rect 16070 -4352 16110 -4350
rect 15710 -4392 15780 -4352
rect 15820 -4392 15890 -4352
rect 15930 -4392 16000 -4352
rect 16040 -4392 16110 -4352
rect 15710 -4420 15750 -4392
rect 15750 -4420 15780 -4392
rect 15820 -4420 15830 -4392
rect 15830 -4420 15870 -4392
rect 15870 -4420 15890 -4392
rect 15930 -4420 15950 -4392
rect 15950 -4420 15990 -4392
rect 15990 -4420 16000 -4392
rect 16040 -4420 16070 -4392
rect 16070 -4420 16110 -4392
rect 15710 -4472 15780 -4460
rect 15820 -4472 15890 -4460
rect 15930 -4472 16000 -4460
rect 16040 -4472 16110 -4460
rect 15710 -4512 15750 -4472
rect 15750 -4512 15780 -4472
rect 15820 -4512 15830 -4472
rect 15830 -4512 15870 -4472
rect 15870 -4512 15890 -4472
rect 15930 -4512 15950 -4472
rect 15950 -4512 15990 -4472
rect 15990 -4512 16000 -4472
rect 16040 -4512 16070 -4472
rect 16070 -4512 16110 -4472
rect 15710 -4530 15780 -4512
rect 15820 -4530 15890 -4512
rect 15930 -4530 16000 -4512
rect 16040 -4530 16110 -4512
rect -1710 -6530 -1700 -6520
rect -1700 -6530 -1640 -6520
rect -1710 -6570 -1640 -6530
rect -1710 -6590 -1700 -6570
rect -1700 -6590 -1640 -6570
rect 7050 -6520 7110 -6460
rect 7150 -6520 7210 -6460
rect 7250 -6520 7310 -6460
rect 7590 -6520 7650 -6460
rect 7690 -6520 7750 -6460
rect 7790 -6520 7850 -6460
rect 7050 -6620 7110 -6560
rect 7150 -6620 7210 -6560
rect 7250 -6620 7310 -6560
rect 7590 -6620 7650 -6560
rect 7690 -6620 7750 -6560
rect 7790 -6620 7850 -6560
rect -1710 -6650 -1640 -6630
rect -1710 -6690 -1700 -6650
rect -1700 -6690 -1640 -6650
rect -1710 -6700 -1640 -6690
rect 4770 -6730 4830 -6670
rect 4870 -6730 4930 -6670
rect 4970 -6730 5030 -6670
rect 7050 -6720 7110 -6660
rect 7150 -6720 7210 -6660
rect 7250 -6720 7310 -6660
rect 7590 -6720 7650 -6660
rect 7690 -6720 7750 -6660
rect 7790 -6720 7850 -6660
rect 16420 -6530 16480 -6520
rect 16480 -6530 16490 -6520
rect 16420 -6570 16490 -6530
rect 16420 -6590 16480 -6570
rect 16480 -6590 16490 -6570
rect -1710 -6770 -1700 -6740
rect -1700 -6770 -1640 -6740
rect -1710 -6810 -1640 -6770
rect -1710 -6890 -1640 -6850
rect -1710 -6920 -1700 -6890
rect -1700 -6920 -1640 -6890
rect 9870 -6730 9930 -6670
rect 9970 -6730 10030 -6670
rect 10070 -6730 10130 -6670
rect 16420 -6650 16490 -6630
rect 16420 -6690 16480 -6650
rect 16480 -6690 16490 -6650
rect 16420 -6700 16490 -6690
rect 4770 -6830 4830 -6770
rect 4870 -6830 4930 -6770
rect 4970 -6830 5030 -6770
rect 7050 -6820 7110 -6760
rect 7150 -6820 7210 -6760
rect 7250 -6820 7310 -6760
rect 7590 -6820 7650 -6760
rect 7690 -6820 7750 -6760
rect 7790 -6820 7850 -6760
rect 9870 -6830 9930 -6770
rect 9970 -6830 10030 -6770
rect 10070 -6830 10130 -6770
rect 4770 -6930 4830 -6870
rect 4870 -6930 4930 -6870
rect 4970 -6930 5030 -6870
rect 9870 -6930 9930 -6870
rect 9970 -6930 10030 -6870
rect 10070 -6930 10130 -6870
rect 16420 -6770 16480 -6740
rect 16480 -6770 16490 -6740
rect 16420 -6810 16490 -6770
rect 16420 -6890 16490 -6850
rect 16420 -6920 16480 -6890
rect 16480 -6920 16490 -6890
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect 21630 -8430 21700 -8360
rect 21730 -8430 21800 -8360
rect 21830 -8430 21900 -8360
rect 21630 -8530 21700 -8460
rect 21730 -8530 21800 -8460
rect 21830 -8530 21900 -8460
rect 21630 -8630 21700 -8560
rect 21730 -8630 21800 -8560
rect 21830 -8630 21900 -8560
rect 22650 -9080 22720 -9010
rect 22750 -9080 22820 -9010
rect 22850 -9080 22920 -9010
rect 22650 -9180 22720 -9110
rect 22750 -9180 22820 -9110
rect 22850 -9180 22920 -9110
rect 22650 -9280 22720 -9210
rect 22750 -9280 22820 -9210
rect 22850 -9280 22920 -9210
rect -240 -9700 -210 -9660
rect -210 -9700 -170 -9660
rect -130 -9700 -90 -9660
rect -90 -9700 -60 -9660
rect -20 -9700 -10 -9660
rect -10 -9700 30 -9660
rect 30 -9700 50 -9660
rect 90 -9700 110 -9660
rect 110 -9700 150 -9660
rect 150 -9700 160 -9660
rect -240 -9730 -170 -9700
rect -130 -9730 -60 -9700
rect -20 -9730 50 -9700
rect 90 -9730 160 -9700
rect -240 -9820 -170 -9790
rect -130 -9820 -60 -9790
rect -20 -9820 50 -9790
rect 90 -9820 160 -9790
rect -240 -9860 -210 -9820
rect -210 -9860 -170 -9820
rect -130 -9860 -90 -9820
rect -90 -9860 -60 -9820
rect -20 -9860 -10 -9820
rect -10 -9860 30 -9820
rect 30 -9860 50 -9820
rect 90 -9860 110 -9820
rect 110 -9860 150 -9820
rect 150 -9860 160 -9820
rect 7240 -9660 7300 -9640
rect 7340 -9660 7400 -9640
rect 7500 -9660 7560 -9640
rect 7600 -9660 7660 -9640
rect 7240 -9700 7270 -9660
rect 7270 -9700 7300 -9660
rect 7340 -9700 7350 -9660
rect 7350 -9700 7390 -9660
rect 7390 -9700 7400 -9660
rect 7500 -9700 7510 -9660
rect 7510 -9700 7550 -9660
rect 7550 -9700 7560 -9660
rect 7600 -9700 7630 -9660
rect 7630 -9700 7660 -9660
rect 7240 -9740 7300 -9730
rect 7340 -9740 7400 -9730
rect 7500 -9740 7560 -9730
rect 7600 -9740 7660 -9730
rect 7240 -9780 7270 -9740
rect 7270 -9780 7300 -9740
rect 7340 -9780 7350 -9740
rect 7350 -9780 7390 -9740
rect 7390 -9780 7400 -9740
rect 7500 -9780 7510 -9740
rect 7510 -9780 7550 -9740
rect 7550 -9780 7560 -9740
rect 7600 -9780 7630 -9740
rect 7630 -9780 7660 -9740
rect 7240 -9790 7300 -9780
rect 7340 -9790 7400 -9780
rect 7500 -9790 7560 -9780
rect 7600 -9790 7660 -9780
rect 7240 -9860 7270 -9820
rect 7270 -9860 7300 -9820
rect 7340 -9860 7350 -9820
rect 7350 -9860 7390 -9820
rect 7390 -9860 7400 -9820
rect 7500 -9860 7510 -9820
rect 7510 -9860 7550 -9820
rect 7550 -9860 7560 -9820
rect 7600 -9860 7630 -9820
rect 7630 -9860 7660 -9820
rect 7240 -9880 7300 -9860
rect 7340 -9880 7400 -9860
rect 7500 -9880 7560 -9860
rect 7600 -9880 7660 -9860
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 14720 -9700 14750 -9660
rect 14750 -9700 14790 -9660
rect 14830 -9700 14870 -9660
rect 14870 -9700 14900 -9660
rect 14940 -9700 14950 -9660
rect 14950 -9700 14990 -9660
rect 14990 -9700 15010 -9660
rect 15050 -9700 15070 -9660
rect 15070 -9700 15110 -9660
rect 15110 -9700 15120 -9660
rect 14720 -9730 14790 -9700
rect 14830 -9730 14900 -9700
rect 14940 -9730 15010 -9700
rect 15050 -9730 15120 -9700
rect 14720 -9820 14790 -9790
rect 14830 -9820 14900 -9790
rect 14940 -9820 15010 -9790
rect 15050 -9820 15120 -9790
rect 14720 -9860 14750 -9820
rect 14750 -9860 14790 -9820
rect 14830 -9860 14870 -9820
rect 14870 -9860 14900 -9820
rect 14940 -9860 14950 -9820
rect 14950 -9860 14990 -9820
rect 14990 -9860 15010 -9820
rect 15050 -9860 15070 -9820
rect 15070 -9860 15110 -9820
rect 15110 -9860 15120 -9820
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 2240 -12370 2310 -12300
rect 2350 -12370 2420 -12300
rect 2460 -12370 2530 -12300
rect 2570 -12370 2640 -12300
rect 2680 -12370 2750 -12300
rect 2790 -12370 2860 -12300
rect 2900 -12370 2970 -12300
rect 3010 -12370 3080 -12300
rect 3120 -12370 3190 -12300
rect 3230 -12370 3300 -12300
rect 3340 -12370 3410 -12300
rect 3450 -12370 3520 -12300
rect 3560 -12370 3630 -12300
rect 3670 -12370 3740 -12300
rect 2240 -12480 2310 -12410
rect 2350 -12480 2420 -12410
rect 2460 -12480 2530 -12410
rect 2570 -12480 2640 -12410
rect 2680 -12480 2750 -12410
rect 2790 -12480 2860 -12410
rect 2900 -12480 2970 -12410
rect 3010 -12480 3080 -12410
rect 3120 -12480 3190 -12410
rect 3230 -12480 3300 -12410
rect 3340 -12480 3410 -12410
rect 3450 -12480 3520 -12410
rect 3560 -12480 3630 -12410
rect 3670 -12480 3740 -12410
rect 11120 -12370 11190 -12300
rect 11230 -12370 11300 -12300
rect 11340 -12370 11410 -12300
rect 11450 -12370 11520 -12300
rect 11560 -12370 11630 -12300
rect 11670 -12370 11740 -12300
rect 11780 -12370 11850 -12300
rect 11890 -12370 11960 -12300
rect 12000 -12370 12070 -12300
rect 12110 -12370 12180 -12300
rect 12220 -12370 12290 -12300
rect 12330 -12370 12400 -12300
rect 12440 -12370 12510 -12300
rect 12550 -12370 12620 -12300
rect 11120 -12480 11190 -12410
rect 11230 -12480 11300 -12410
rect 11340 -12480 11410 -12410
rect 11450 -12480 11520 -12410
rect 11560 -12480 11630 -12410
rect 11670 -12480 11740 -12410
rect 11780 -12480 11850 -12410
rect 11890 -12480 11960 -12410
rect 12000 -12480 12070 -12410
rect 12110 -12480 12180 -12410
rect 12220 -12480 12290 -12410
rect 12330 -12480 12400 -12410
rect 12440 -12480 12510 -12410
rect 12550 -12480 12620 -12410
rect 7010 -13310 7070 -13250
rect 7110 -13310 7170 -13250
rect 7210 -13310 7270 -13250
rect 7630 -13310 7690 -13250
rect 7730 -13310 7790 -13250
rect 7830 -13310 7890 -13250
rect 7010 -13400 7070 -13340
rect 7110 -13400 7170 -13340
rect 7210 -13400 7270 -13340
rect 7630 -13400 7690 -13340
rect 7730 -13400 7790 -13340
rect 7830 -13400 7890 -13340
rect 7010 -13490 7070 -13430
rect 7110 -13490 7170 -13430
rect 7210 -13490 7270 -13430
rect 7630 -13490 7690 -13430
rect 7730 -13490 7790 -13430
rect 7830 -13490 7890 -13430
rect 7010 -13590 7070 -13530
rect 7110 -13590 7170 -13530
rect 7210 -13590 7270 -13530
rect 7630 -13590 7690 -13530
rect 7730 -13590 7790 -13530
rect 7830 -13590 7890 -13530
rect 7010 -13680 7070 -13620
rect 7110 -13680 7170 -13620
rect 7210 -13680 7270 -13620
rect 7630 -13680 7690 -13620
rect 7730 -13680 7790 -13620
rect 7830 -13680 7890 -13620
rect 7010 -13770 7070 -13710
rect 7110 -13770 7170 -13710
rect 7210 -13770 7270 -13710
rect 7630 -13770 7690 -13710
rect 7730 -13770 7790 -13710
rect 7830 -13770 7890 -13710
rect 21630 -14090 21700 -14020
rect 21730 -14090 21800 -14020
rect 21830 -14090 21900 -14020
rect 21630 -14190 21700 -14120
rect 21730 -14190 21800 -14120
rect 21830 -14190 21900 -14120
rect 21630 -14290 21700 -14220
rect 21730 -14290 21800 -14220
rect 21830 -14290 21900 -14220
rect 22920 -14940 22990 -14870
rect 23020 -14940 23090 -14870
rect 23120 -14940 23190 -14870
rect 22920 -15040 22990 -14970
rect 23020 -15040 23090 -14970
rect 23120 -15040 23190 -14970
rect 22920 -15140 22990 -15070
rect 23020 -15140 23090 -15070
rect 23120 -15140 23190 -15070
rect 5040 -17160 5100 -17100
rect 5140 -17160 5200 -17100
rect 5240 -17160 5300 -17100
rect 9600 -17160 9660 -17100
rect 9700 -17160 9760 -17100
rect 9800 -17160 9860 -17100
rect 5040 -17260 5100 -17200
rect 5140 -17260 5200 -17200
rect 5240 -17260 5300 -17200
rect 9600 -17260 9660 -17200
rect 9700 -17260 9760 -17200
rect 9800 -17260 9860 -17200
rect 5040 -17360 5100 -17300
rect 5140 -17360 5200 -17300
rect 5240 -17360 5300 -17300
rect 9600 -17360 9660 -17300
rect 9700 -17360 9760 -17300
rect 9800 -17360 9860 -17300
rect 7230 -17670 7300 -17600
rect 7340 -17670 7410 -17600
rect 7450 -17670 7520 -17600
rect 7560 -17670 7630 -17600
rect 7230 -17780 7300 -17710
rect 7340 -17780 7410 -17710
rect 7450 -17780 7520 -17710
rect 7560 -17780 7630 -17710
rect 7230 -17890 7300 -17820
rect 7340 -17890 7410 -17820
rect 7450 -17890 7520 -17820
rect 7560 -17890 7630 -17820
rect 7230 -18000 7300 -17930
rect 7340 -18000 7410 -17930
rect 7450 -18000 7520 -17930
rect 7560 -18000 7630 -17930
rect 21630 -20170 21700 -20100
rect 21730 -20170 21800 -20100
rect 21830 -20170 21900 -20100
rect 21630 -20270 21700 -20200
rect 21730 -20270 21800 -20200
rect 21830 -20270 21900 -20200
rect 21630 -20370 21700 -20300
rect 21730 -20370 21800 -20300
rect 21830 -20370 21900 -20300
rect 22700 -20800 22770 -20730
rect 22800 -20800 22870 -20730
rect 22900 -20800 22970 -20730
rect 22700 -20900 22770 -20830
rect 22800 -20900 22870 -20830
rect 22900 -20900 22970 -20830
rect 22700 -21000 22770 -20930
rect 22800 -21000 22870 -20930
rect 22900 -21000 22970 -20930
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 3160 -22730 3230 -22660
rect 3270 -22730 3340 -22660
rect 3380 -22730 3450 -22660
rect 3490 -22730 3560 -22660
rect 3600 -22730 3670 -22660
rect 3710 -22730 3780 -22660
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 3160 -22840 3230 -22770
rect 3270 -22840 3340 -22770
rect 3380 -22840 3450 -22770
rect 3490 -22840 3560 -22770
rect 3600 -22840 3670 -22770
rect 3710 -22840 3780 -22770
rect 11160 -22730 11230 -22660
rect 11270 -22730 11340 -22660
rect 11380 -22730 11450 -22660
rect 11490 -22730 11560 -22660
rect 11600 -22730 11670 -22660
rect 11710 -22730 11780 -22660
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 11160 -22840 11230 -22770
rect 11270 -22840 11340 -22770
rect 11380 -22840 11450 -22770
rect 11490 -22840 11560 -22770
rect 11600 -22840 11670 -22770
rect 11710 -22840 11780 -22770
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
<< metal2 >>
rect 23460 7210 23940 7260
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 25860 7210 26340 7260
rect 25860 7140 25890 7210
rect 25960 7140 26000 7210
rect 26070 7140 26110 7210
rect 26180 7140 26220 7210
rect 26290 7140 26340 7210
rect 25860 7100 26340 7140
rect 25860 7030 25890 7100
rect 25960 7030 26000 7100
rect 26070 7030 26110 7100
rect 26180 7030 26220 7100
rect 26290 7030 26340 7100
rect 25860 7000 26340 7030
rect 1540 6850 3140 6900
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 11760 6880 13360 6930
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 1540 6640 3140 6670
rect 7350 6300 30940 6320
rect 7350 6290 30740 6300
rect 7350 6230 7380 6290
rect 7440 6230 7480 6290
rect 7540 6280 30740 6290
rect 7540 6230 22780 6280
rect 7350 6210 22780 6230
rect 22850 6210 22890 6280
rect 22960 6210 23000 6280
rect 23070 6210 23110 6280
rect 23180 6230 30740 6280
rect 30810 6230 30850 6300
rect 30920 6230 30940 6300
rect 23180 6210 30940 6230
rect 7350 6190 30940 6210
rect 7350 6080 7380 6190
rect 7440 6080 7480 6190
rect 7540 6170 30940 6190
rect 7540 6100 22780 6170
rect 22850 6100 22890 6170
rect 22960 6100 23000 6170
rect 23070 6100 23110 6170
rect 23180 6100 30740 6170
rect 30810 6100 30850 6170
rect 30920 6100 30940 6170
rect 7540 6080 30940 6100
rect 7350 6060 30940 6080
rect 7350 6040 22780 6060
rect 7350 5980 7380 6040
rect 7440 5980 7480 6040
rect 7540 5990 22780 6040
rect 22850 5990 22890 6060
rect 22960 5990 23000 6060
rect 23070 5990 23110 6060
rect 23180 6040 30940 6060
rect 23180 5990 30740 6040
rect 7540 5980 30740 5990
rect 7350 5970 30740 5980
rect 30810 5970 30850 6040
rect 30920 5970 30940 6040
rect 7350 5950 30940 5970
rect 21800 5670 22020 5690
rect 21800 5600 21820 5670
rect 21890 5600 21930 5670
rect 22000 5600 22020 5670
rect 21800 5560 22020 5600
rect 21800 5490 21820 5560
rect 21890 5490 21930 5560
rect 22000 5490 22020 5560
rect 21800 5450 22020 5490
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 21800 5380 21820 5450
rect 21890 5380 21930 5450
rect 22000 5380 22020 5450
rect 21800 5340 22020 5380
rect 21800 5270 21820 5340
rect 21890 5270 21930 5340
rect 22000 5270 22020 5340
rect 21800 5230 22020 5270
rect 21800 5160 21820 5230
rect 21890 5160 21930 5230
rect 22000 5160 22020 5230
rect 21800 5120 22020 5160
rect 21800 5050 21820 5120
rect 21890 5050 21930 5120
rect 22000 5050 22020 5120
rect 21800 5010 22020 5050
rect 21800 4940 21820 5010
rect 21890 4940 21930 5010
rect 22000 4940 22020 5010
rect 21800 4900 22020 4940
rect 21800 4830 21820 4900
rect 21890 4830 21930 4900
rect 22000 4830 22020 4900
rect 21800 4790 22020 4830
rect 7560 4760 7880 4790
rect 7560 4700 7590 4760
rect 7650 4700 7690 4760
rect 7750 4700 7790 4760
rect 7850 4700 7880 4760
rect 7560 4610 7880 4700
rect 21800 4720 21820 4790
rect 21890 4720 21930 4790
rect 22000 4720 22020 4790
rect 21800 4680 22020 4720
rect 21800 4610 21820 4680
rect 21890 4610 21930 4680
rect 22000 4610 22020 4680
rect -1740 4580 -1600 4610
rect -1740 4510 -1710 4580
rect -1640 4510 -1600 4580
rect -1740 4470 -1600 4510
rect -1740 4400 -1710 4470
rect -1640 4400 -1600 4470
rect -1740 4360 -1600 4400
rect -1740 4290 -1710 4360
rect -1640 4290 -1600 4360
rect -1740 4250 -1600 4290
rect -1740 4180 -1710 4250
rect -1640 4180 -1600 4250
rect -1740 4130 -1600 4180
rect 6670 4580 7880 4610
rect 6670 4520 6700 4580
rect 6760 4520 7880 4580
rect 6670 4460 7880 4520
rect 6670 4400 6700 4460
rect 6760 4400 7880 4460
rect 6670 4340 7880 4400
rect 6670 4280 6700 4340
rect 6760 4280 7880 4340
rect 6670 4220 7880 4280
rect 6670 4160 6700 4220
rect 6760 4160 7880 4220
rect 6670 4130 7880 4160
rect 16380 4580 16520 4610
rect 16380 4510 16420 4580
rect 16490 4510 16520 4580
rect 16380 4470 16520 4510
rect 21800 4570 22020 4610
rect 21800 4500 21820 4570
rect 21890 4500 21930 4570
rect 22000 4500 22020 4570
rect 21800 4480 22020 4500
rect 27680 4870 28280 4900
rect 27680 4810 27710 4870
rect 27770 4810 27810 4870
rect 27870 4810 27910 4870
rect 27970 4810 28280 4870
rect 27680 4770 28280 4810
rect 27680 4710 27710 4770
rect 27770 4710 27810 4770
rect 27870 4710 27910 4770
rect 27970 4710 28280 4770
rect 27680 4670 28280 4710
rect 27680 4610 27710 4670
rect 27770 4610 27810 4670
rect 27870 4610 27910 4670
rect 27970 4610 28280 4670
rect 27680 4570 28280 4610
rect 27680 4510 27710 4570
rect 27770 4510 27810 4570
rect 27870 4510 27910 4570
rect 27970 4510 28280 4570
rect 16380 4400 16420 4470
rect 16490 4400 16520 4470
rect 16380 4360 16520 4400
rect 16380 4290 16420 4360
rect 16490 4290 16520 4360
rect 16380 4250 16520 4290
rect 16380 4180 16420 4250
rect 16490 4180 16520 4250
rect 16380 4130 16520 4180
rect 27680 4470 28280 4510
rect 27680 4410 27710 4470
rect 27770 4410 27810 4470
rect 27870 4410 27910 4470
rect 27970 4410 28280 4470
rect 27680 4370 28280 4410
rect 27680 4310 27710 4370
rect 27770 4310 27810 4370
rect 27870 4310 27910 4370
rect 27970 4310 28280 4370
rect 27680 4270 28280 4310
rect 27680 4210 27710 4270
rect 27770 4210 27810 4270
rect 27870 4210 27910 4270
rect 27970 4210 28280 4270
rect 27680 4170 28280 4210
rect 7020 3240 7340 3270
rect 7020 3180 7050 3240
rect 7110 3180 7150 3240
rect 7210 3180 7250 3240
rect 7310 3180 7340 3240
rect 7020 3140 7340 3180
rect 7020 3080 7050 3140
rect 7110 3080 7150 3140
rect 7210 3080 7250 3140
rect 7310 3080 7340 3140
rect 7020 3040 7340 3080
rect 7020 2980 7050 3040
rect 7110 2980 7150 3040
rect 7210 2980 7250 3040
rect 7310 2980 7340 3040
rect 7020 2960 7340 2980
rect 7560 3240 7880 4130
rect 27680 4110 27710 4170
rect 27770 4110 27810 4170
rect 27870 4110 27910 4170
rect 27970 4110 28280 4170
rect 27680 4070 28280 4110
rect 27680 4010 27710 4070
rect 27770 4010 27810 4070
rect 27870 4010 27910 4070
rect 27970 4010 28280 4070
rect 27680 3980 28280 4010
rect 7560 3180 7590 3240
rect 7650 3180 7690 3240
rect 7750 3180 7790 3240
rect 7850 3180 7880 3240
rect 7560 3140 7880 3180
rect 7560 3080 7590 3140
rect 7650 3080 7690 3140
rect 7750 3080 7790 3140
rect 7850 3080 7880 3140
rect 7560 3040 7880 3080
rect 24700 3360 25030 3380
rect 24700 3290 24720 3360
rect 24790 3290 24830 3360
rect 24900 3290 24940 3360
rect 25010 3290 25030 3360
rect 24700 3250 25030 3290
rect 24700 3180 24720 3250
rect 24790 3180 24830 3250
rect 24900 3180 24940 3250
rect 25010 3180 25030 3250
rect 24700 3140 25030 3180
rect 24700 3070 24720 3140
rect 24790 3070 24830 3140
rect 24900 3070 24940 3140
rect 25010 3070 25030 3140
rect 24700 3050 25030 3070
rect 7560 2980 7590 3040
rect 7650 2980 7690 3040
rect 7750 2980 7790 3040
rect 7850 2980 7880 3040
rect 7560 2960 7880 2980
rect 4740 2890 5060 2920
rect 4740 2830 4770 2890
rect 4830 2830 4870 2890
rect 4930 2830 4970 2890
rect 5030 2830 5060 2890
rect 4740 2790 5060 2830
rect 4740 2730 4770 2790
rect 4830 2730 4870 2790
rect 4930 2730 4970 2790
rect 5030 2730 5060 2790
rect 4740 2690 5060 2730
rect 4740 2630 4770 2690
rect 4830 2630 4870 2690
rect 4930 2630 4970 2690
rect 5030 2630 5060 2690
rect 4740 2610 5060 2630
rect 9840 2890 10160 2920
rect 9840 2830 9870 2890
rect 9930 2830 9970 2890
rect 10030 2830 10070 2890
rect 10130 2830 10160 2890
rect 9840 2790 10160 2830
rect 9840 2730 9870 2790
rect 9930 2730 9970 2790
rect 10030 2730 10070 2790
rect 10130 2730 10160 2790
rect 9840 2690 10160 2730
rect 9840 2630 9870 2690
rect 9930 2630 9970 2690
rect 10030 2630 10070 2690
rect 10130 2630 10160 2690
rect 9840 2610 10160 2630
rect 22420 2600 22900 2630
rect 22420 2530 22470 2600
rect 22540 2530 22580 2600
rect 22650 2530 22690 2600
rect 22760 2530 22800 2600
rect 22870 2530 22900 2600
rect 22420 2490 22900 2530
rect 22420 2420 22470 2490
rect 22540 2420 22580 2490
rect 22650 2420 22690 2490
rect 22760 2420 22800 2490
rect 22870 2420 22900 2490
rect 22420 2370 22900 2420
rect 26900 2600 27380 2630
rect 26900 2530 26950 2600
rect 27020 2530 27060 2600
rect 27130 2530 27170 2600
rect 27240 2530 27280 2600
rect 27350 2530 27380 2600
rect 26900 2490 27380 2530
rect 26900 2420 26950 2490
rect 27020 2420 27060 2490
rect 27130 2420 27170 2490
rect 27240 2420 27280 2490
rect 27350 2420 27380 2490
rect 26900 2370 27380 2420
rect 28040 1980 28280 3980
rect 7150 1740 28280 1980
rect -330 -140 150 -100
rect -330 -210 -300 -140
rect -230 -210 -190 -140
rect -120 -210 -80 -140
rect -10 -210 30 -140
rect 100 -210 150 -140
rect -330 -270 150 -210
rect -330 -340 -300 -270
rect -230 -340 -190 -270
rect -120 -340 -80 -270
rect -10 -340 30 -270
rect 100 -340 150 -270
rect -330 -380 150 -340
rect 7150 -120 7630 1740
rect 14590 1160 14900 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 14900 1160
rect 14590 1050 14900 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 14900 1050
rect 14590 940 14900 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 14900 940
rect 14590 850 14900 870
rect 23460 920 23940 970
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 25860 920 26340 970
rect 25860 850 25890 920
rect 25960 850 26000 920
rect 26070 850 26110 920
rect 26180 850 26220 920
rect 26290 850 26340 920
rect 25860 810 26340 850
rect 25860 740 25890 810
rect 25960 740 26000 810
rect 26070 740 26110 810
rect 26180 740 26220 810
rect 26290 740 26340 810
rect 25860 710 26340 740
rect 19440 0 30940 20
rect 19440 -20 30740 0
rect 19440 -90 22780 -20
rect 22850 -90 22890 -20
rect 22960 -90 23000 -20
rect 23070 -90 23110 -20
rect 23180 -70 30740 -20
rect 30810 -70 30850 0
rect 30920 -70 30940 0
rect 23180 -90 30940 -70
rect 7150 -180 7180 -120
rect 7240 -180 7280 -120
rect 7340 -180 7440 -120
rect 7500 -180 7540 -120
rect 7600 -180 7630 -120
rect 7150 -210 7630 -180
rect 7150 -270 7180 -210
rect 7240 -270 7280 -210
rect 7340 -270 7440 -210
rect 7500 -270 7540 -210
rect 7600 -270 7630 -210
rect 7150 -300 7630 -270
rect 7150 -360 7180 -300
rect 7240 -360 7280 -300
rect 7340 -360 7440 -300
rect 7500 -360 7540 -300
rect 7600 -360 7630 -300
rect 7150 -380 7630 -360
rect 14630 -140 15110 -100
rect 14630 -210 14660 -140
rect 14730 -210 14770 -140
rect 14840 -210 14880 -140
rect 14950 -210 14990 -140
rect 15060 -210 15110 -140
rect 14630 -270 15110 -210
rect 14630 -340 14660 -270
rect 14730 -340 14770 -270
rect 14840 -340 14880 -270
rect 14950 -340 14990 -270
rect 15060 -340 15110 -270
rect 14630 -380 15110 -340
rect 19440 -130 30940 -90
rect 19440 -200 22780 -130
rect 22850 -200 22890 -130
rect 22960 -200 23000 -130
rect 23070 -200 23110 -130
rect 23180 -200 30740 -130
rect 30810 -200 30850 -130
rect 30920 -200 30940 -130
rect 19440 -240 30940 -200
rect 19440 -310 22780 -240
rect 22850 -310 22890 -240
rect 22960 -310 23000 -240
rect 23070 -310 23110 -240
rect 23180 -260 30940 -240
rect 23180 -310 30740 -260
rect 19440 -330 30740 -310
rect 30810 -330 30850 -260
rect 30920 -330 30940 -260
rect 19440 -350 30940 -330
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1020 2680 -970
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1020 13820 -970
rect 1540 -2780 3140 -2730
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 11760 -2780 13360 -2730
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect 19440 -3310 19680 -350
rect 21800 -850 22020 -830
rect 21800 -920 21820 -850
rect 21890 -920 21930 -850
rect 22000 -920 22020 -850
rect 21800 -960 22020 -920
rect 21800 -1030 21820 -960
rect 21890 -1030 21930 -960
rect 22000 -1030 22020 -960
rect 21800 -1070 22020 -1030
rect 21800 -1140 21820 -1070
rect 21890 -1140 21930 -1070
rect 22000 -1140 22020 -1070
rect 21800 -1180 22020 -1140
rect 21800 -1250 21820 -1180
rect 21890 -1250 21930 -1180
rect 22000 -1250 22020 -1180
rect 21800 -1290 22020 -1250
rect 21800 -1360 21820 -1290
rect 21890 -1360 21930 -1290
rect 22000 -1360 22020 -1290
rect 21800 -1400 22020 -1360
rect 21800 -1470 21820 -1400
rect 21890 -1470 21930 -1400
rect 22000 -1470 22020 -1400
rect 21800 -1510 22020 -1470
rect 21800 -1580 21820 -1510
rect 21890 -1580 21930 -1510
rect 22000 -1580 22020 -1510
rect 21800 -1620 22020 -1580
rect 21800 -1690 21820 -1620
rect 21890 -1690 21930 -1620
rect 22000 -1690 22020 -1620
rect 21800 -1730 22020 -1690
rect 21800 -1800 21820 -1730
rect 21890 -1800 21930 -1730
rect 22000 -1800 22020 -1730
rect 21800 -1840 22020 -1800
rect 21800 -1910 21820 -1840
rect 21890 -1910 21930 -1840
rect 22000 -1910 22020 -1840
rect 21800 -1950 22020 -1910
rect 21800 -2020 21820 -1950
rect 21890 -2020 21930 -1950
rect 22000 -2020 22020 -1950
rect 21800 -2040 22020 -2020
rect 27680 -1430 28280 -1400
rect 27680 -1490 27710 -1430
rect 27770 -1490 27810 -1430
rect 27870 -1490 27910 -1430
rect 27970 -1490 28280 -1430
rect 27680 -1530 28280 -1490
rect 27680 -1590 27710 -1530
rect 27770 -1590 27810 -1530
rect 27870 -1590 27910 -1530
rect 27970 -1590 28280 -1530
rect 27680 -1630 28280 -1590
rect 27680 -1690 27710 -1630
rect 27770 -1690 27810 -1630
rect 27870 -1690 27910 -1630
rect 27970 -1690 28280 -1630
rect 27680 -1730 28280 -1690
rect 27680 -1790 27710 -1730
rect 27770 -1790 27810 -1730
rect 27870 -1790 27910 -1730
rect 27970 -1790 28280 -1730
rect 27680 -1830 28280 -1790
rect 27680 -1890 27710 -1830
rect 27770 -1890 27810 -1830
rect 27870 -1890 27910 -1830
rect 27970 -1890 28280 -1830
rect 27680 -1930 28280 -1890
rect 27680 -1990 27710 -1930
rect 27770 -1990 27810 -1930
rect 27870 -1990 27910 -1930
rect 27970 -1990 28280 -1930
rect 27680 -2030 28280 -1990
rect 27680 -2090 27710 -2030
rect 27770 -2090 27810 -2030
rect 27870 -2090 27910 -2030
rect 27970 -2090 28280 -2030
rect 27680 -2130 28280 -2090
rect 27680 -2190 27710 -2130
rect 27770 -2190 27810 -2130
rect 27870 -2190 27910 -2130
rect 27970 -2190 28280 -2130
rect 27680 -2230 28280 -2190
rect 27680 -2290 27710 -2230
rect 27770 -2290 27810 -2230
rect 27870 -2290 27910 -2230
rect 27970 -2290 28280 -2230
rect 27680 -2320 28280 -2290
rect 7350 -3340 19680 -3310
rect 7350 -3400 7380 -3340
rect 7440 -3400 7480 -3340
rect 7540 -3400 19680 -3340
rect 24720 -3050 25050 -3030
rect 24720 -3120 24740 -3050
rect 24810 -3120 24850 -3050
rect 24920 -3120 24960 -3050
rect 25030 -3120 25050 -3050
rect 24720 -3160 25050 -3120
rect 24720 -3230 24740 -3160
rect 24810 -3230 24850 -3160
rect 24920 -3230 24960 -3160
rect 25030 -3230 25050 -3160
rect 24720 -3270 25050 -3230
rect 24720 -3340 24740 -3270
rect 24810 -3340 24850 -3270
rect 24920 -3340 24960 -3270
rect 25030 -3340 25050 -3270
rect 24720 -3360 25050 -3340
rect 7350 -3440 19680 -3400
rect 7350 -3550 7380 -3440
rect 7440 -3550 7480 -3440
rect 7540 -3550 19680 -3440
rect 7350 -3590 19680 -3550
rect 7350 -3650 7380 -3590
rect 7440 -3650 7480 -3590
rect 7540 -3650 19680 -3590
rect 7350 -3680 19680 -3650
rect 22420 -3690 22900 -3660
rect 22420 -3760 22470 -3690
rect 22540 -3760 22580 -3690
rect 22650 -3760 22690 -3690
rect 22760 -3760 22800 -3690
rect 22870 -3760 22900 -3690
rect 22420 -3800 22900 -3760
rect 7290 -3880 7620 -3860
rect 7290 -3950 7310 -3880
rect 7380 -3950 7420 -3880
rect 7490 -3950 7530 -3880
rect 7600 -3950 7620 -3880
rect 22420 -3870 22470 -3800
rect 22540 -3870 22580 -3800
rect 22650 -3870 22690 -3800
rect 22760 -3870 22800 -3800
rect 22870 -3870 22900 -3800
rect 22420 -3920 22900 -3870
rect 26900 -3690 27380 -3660
rect 26900 -3760 26950 -3690
rect 27020 -3760 27060 -3690
rect 27130 -3760 27170 -3690
rect 27240 -3760 27280 -3690
rect 27350 -3760 27380 -3690
rect 26900 -3800 27380 -3760
rect 26900 -3870 26950 -3800
rect 27020 -3870 27060 -3800
rect 27130 -3870 27170 -3800
rect 27240 -3870 27280 -3800
rect 27350 -3870 27380 -3800
rect 26900 -3920 27380 -3870
rect 7290 -3990 7620 -3950
rect 7290 -4060 7310 -3990
rect 7380 -4060 7420 -3990
rect 7490 -4060 7530 -3990
rect 7600 -4060 7620 -3990
rect 7290 -4100 7620 -4060
rect 7290 -4170 7310 -4100
rect 7380 -4170 7420 -4100
rect 7490 -4170 7530 -4100
rect 7600 -4170 7620 -4100
rect 7290 -4190 7620 -4170
rect -580 -4290 -140 -4270
rect -1350 -4350 -910 -4330
rect -1350 -4420 -1330 -4350
rect -1260 -4420 -1220 -4350
rect -1150 -4420 -1110 -4350
rect -1040 -4420 -1000 -4350
rect -930 -4420 -910 -4350
rect -1350 -4460 -910 -4420
rect -1350 -4530 -1330 -4460
rect -1260 -4530 -1220 -4460
rect -1150 -4530 -1110 -4460
rect -1040 -4530 -1000 -4460
rect -930 -4530 -910 -4460
rect -580 -4360 -560 -4290
rect -490 -4360 -450 -4290
rect -380 -4360 -340 -4290
rect -270 -4360 -230 -4290
rect -160 -4360 -140 -4290
rect -580 -4400 -140 -4360
rect -580 -4470 -560 -4400
rect -490 -4470 -450 -4400
rect -380 -4470 -340 -4400
rect -270 -4470 -230 -4400
rect -160 -4470 -140 -4400
rect -580 -4490 -140 -4470
rect 14920 -4290 15360 -4270
rect 14920 -4360 14940 -4290
rect 15010 -4360 15050 -4290
rect 15120 -4360 15160 -4290
rect 15230 -4360 15270 -4290
rect 15340 -4360 15360 -4290
rect 14920 -4400 15360 -4360
rect 14920 -4470 14940 -4400
rect 15010 -4470 15050 -4400
rect 15120 -4470 15160 -4400
rect 15230 -4470 15270 -4400
rect 15340 -4470 15360 -4400
rect 14920 -4490 15360 -4470
rect 15690 -4350 16130 -4330
rect 15690 -4420 15710 -4350
rect 15780 -4420 15820 -4350
rect 15890 -4420 15930 -4350
rect 16000 -4420 16040 -4350
rect 16110 -4420 16130 -4350
rect 28080 -4370 28280 -2320
rect 15690 -4460 16130 -4420
rect -1350 -4550 -910 -4530
rect 15690 -4530 15710 -4460
rect 15780 -4530 15820 -4460
rect 15890 -4530 15930 -4460
rect 16000 -4530 16040 -4460
rect 16110 -4530 16130 -4460
rect 15690 -4550 16130 -4530
rect 20180 -4600 28280 -4370
rect 7030 -6460 7340 -6420
rect -1740 -6520 -1600 -6470
rect -1740 -6590 -1710 -6520
rect -1640 -6590 -1600 -6520
rect -1740 -6630 -1600 -6590
rect -1740 -6700 -1710 -6630
rect -1640 -6700 -1600 -6630
rect 7030 -6520 7050 -6460
rect 7110 -6520 7150 -6460
rect 7210 -6520 7250 -6460
rect 7310 -6520 7340 -6460
rect 7030 -6560 7340 -6520
rect 7030 -6620 7050 -6560
rect 7110 -6620 7150 -6560
rect 7210 -6620 7250 -6560
rect 7310 -6620 7340 -6560
rect -1740 -6740 -1600 -6700
rect -1740 -6810 -1710 -6740
rect -1640 -6810 -1600 -6740
rect -1740 -6850 -1600 -6810
rect -1740 -6920 -1710 -6850
rect -1640 -6920 -1600 -6850
rect -1740 -6950 -1600 -6920
rect 4740 -6670 5060 -6640
rect 4740 -6730 4770 -6670
rect 4830 -6730 4870 -6670
rect 4930 -6730 4970 -6670
rect 5030 -6730 5060 -6670
rect 4740 -6770 5060 -6730
rect 4740 -6830 4770 -6770
rect 4830 -6830 4870 -6770
rect 4930 -6830 4970 -6770
rect 5030 -6830 5060 -6770
rect 4740 -6870 5060 -6830
rect 7030 -6660 7340 -6620
rect 7030 -6720 7050 -6660
rect 7110 -6720 7150 -6660
rect 7210 -6720 7250 -6660
rect 7310 -6720 7340 -6660
rect 7030 -6760 7340 -6720
rect 7030 -6820 7050 -6760
rect 7110 -6820 7150 -6760
rect 7210 -6820 7250 -6760
rect 7310 -6820 7340 -6760
rect 7030 -6850 7340 -6820
rect 7570 -6460 7870 -6420
rect 7570 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 7870 -6460
rect 7570 -6560 7870 -6520
rect 7570 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 7870 -6560
rect 7570 -6660 7870 -6620
rect 16380 -6520 16520 -6470
rect 16380 -6590 16420 -6520
rect 16490 -6590 16520 -6520
rect 16380 -6630 16520 -6590
rect 7570 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 7870 -6660
rect 7570 -6760 7870 -6720
rect 7570 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 7870 -6760
rect 7570 -6850 7870 -6820
rect 9840 -6670 10160 -6640
rect 9840 -6730 9870 -6670
rect 9930 -6730 9970 -6670
rect 10030 -6730 10070 -6670
rect 10130 -6730 10160 -6670
rect 9840 -6770 10160 -6730
rect 9840 -6830 9870 -6770
rect 9930 -6830 9970 -6770
rect 10030 -6830 10070 -6770
rect 10130 -6830 10160 -6770
rect 4740 -6930 4770 -6870
rect 4830 -6930 4870 -6870
rect 4930 -6930 4970 -6870
rect 5030 -6930 5060 -6870
rect 4740 -6950 5060 -6930
rect 9840 -6870 10160 -6830
rect 9840 -6930 9870 -6870
rect 9930 -6930 9970 -6870
rect 10030 -6930 10070 -6870
rect 10130 -6930 10160 -6870
rect 9840 -6950 10160 -6930
rect 16380 -6700 16420 -6630
rect 16490 -6700 16520 -6630
rect 16380 -6740 16520 -6700
rect 16380 -6810 16420 -6740
rect 16490 -6810 16520 -6740
rect 16380 -6850 16520 -6810
rect 16380 -6920 16420 -6850
rect 16490 -6920 16520 -6850
rect 16380 -6950 16520 -6920
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 20180 -9160 20490 -4600
rect 21610 -8360 21930 -8330
rect 21610 -8430 21630 -8360
rect 21700 -8430 21730 -8360
rect 21800 -8430 21830 -8360
rect 21900 -8430 21930 -8360
rect 21610 -8460 21930 -8430
rect 21610 -8530 21630 -8460
rect 21700 -8530 21730 -8460
rect 21800 -8530 21830 -8460
rect 21900 -8530 21930 -8460
rect 21610 -8560 21930 -8530
rect 21610 -8630 21630 -8560
rect 21700 -8630 21730 -8560
rect 21800 -8630 21830 -8560
rect 21900 -8630 21930 -8560
rect 21610 -8650 21930 -8630
rect 7210 -9440 20490 -9160
rect 22630 -9010 22950 -8980
rect 22630 -9080 22650 -9010
rect 22720 -9080 22750 -9010
rect 22820 -9080 22850 -9010
rect 22920 -9080 22950 -9010
rect 22630 -9110 22950 -9080
rect 22630 -9180 22650 -9110
rect 22720 -9180 22750 -9110
rect 22820 -9180 22850 -9110
rect 22920 -9180 22950 -9110
rect 22630 -9210 22950 -9180
rect 22630 -9280 22650 -9210
rect 22720 -9280 22750 -9210
rect 22820 -9280 22850 -9210
rect 22920 -9280 22950 -9210
rect 22630 -9300 22950 -9280
rect -270 -9660 210 -9620
rect -270 -9730 -240 -9660
rect -170 -9730 -130 -9660
rect -60 -9730 -20 -9660
rect 50 -9730 90 -9660
rect 160 -9730 210 -9660
rect -270 -9790 210 -9730
rect -270 -9860 -240 -9790
rect -170 -9860 -130 -9790
rect -60 -9860 -20 -9790
rect 50 -9860 90 -9790
rect 160 -9860 210 -9790
rect -270 -9900 210 -9860
rect 7210 -9640 7690 -9440
rect 7210 -9700 7240 -9640
rect 7300 -9700 7340 -9640
rect 7400 -9700 7500 -9640
rect 7560 -9700 7600 -9640
rect 7660 -9700 7690 -9640
rect 7210 -9730 7690 -9700
rect 7210 -9790 7240 -9730
rect 7300 -9790 7340 -9730
rect 7400 -9790 7500 -9730
rect 7560 -9790 7600 -9730
rect 7660 -9790 7690 -9730
rect 7210 -9820 7690 -9790
rect 7210 -9880 7240 -9820
rect 7300 -9880 7340 -9820
rect 7400 -9880 7500 -9820
rect 7560 -9880 7600 -9820
rect 7660 -9880 7690 -9820
rect 7210 -9900 7690 -9880
rect 14690 -9660 15170 -9620
rect 14690 -9730 14720 -9660
rect 14790 -9730 14830 -9660
rect 14900 -9730 14940 -9660
rect 15010 -9730 15050 -9660
rect 15120 -9730 15170 -9660
rect 14690 -9790 15170 -9730
rect 14690 -9860 14720 -9790
rect 14790 -9860 14830 -9790
rect 14900 -9860 14940 -9790
rect 15010 -9860 15050 -9790
rect 15120 -9860 15170 -9790
rect 14690 -9900 15170 -9860
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10570 2680 -10520
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10600 13820 -10550
rect 2210 -12300 3810 -12250
rect 2210 -12370 2240 -12300
rect 2310 -12370 2350 -12300
rect 2420 -12370 2460 -12300
rect 2530 -12370 2570 -12300
rect 2640 -12370 2680 -12300
rect 2750 -12370 2790 -12300
rect 2860 -12370 2900 -12300
rect 2970 -12370 3010 -12300
rect 3080 -12370 3120 -12300
rect 3190 -12370 3230 -12300
rect 3300 -12370 3340 -12300
rect 3410 -12370 3450 -12300
rect 3520 -12370 3560 -12300
rect 3630 -12370 3670 -12300
rect 3740 -12370 3810 -12300
rect 2210 -12410 3810 -12370
rect 2210 -12480 2240 -12410
rect 2310 -12480 2350 -12410
rect 2420 -12480 2460 -12410
rect 2530 -12480 2570 -12410
rect 2640 -12480 2680 -12410
rect 2750 -12480 2790 -12410
rect 2860 -12480 2900 -12410
rect 2970 -12480 3010 -12410
rect 3080 -12480 3120 -12410
rect 3190 -12480 3230 -12410
rect 3300 -12480 3340 -12410
rect 3410 -12480 3450 -12410
rect 3520 -12480 3560 -12410
rect 3630 -12480 3670 -12410
rect 3740 -12480 3810 -12410
rect 2210 -12510 3810 -12480
rect 11090 -12300 12690 -12250
rect 11090 -12370 11120 -12300
rect 11190 -12370 11230 -12300
rect 11300 -12370 11340 -12300
rect 11410 -12370 11450 -12300
rect 11520 -12370 11560 -12300
rect 11630 -12370 11670 -12300
rect 11740 -12370 11780 -12300
rect 11850 -12370 11890 -12300
rect 11960 -12370 12000 -12300
rect 12070 -12370 12110 -12300
rect 12180 -12370 12220 -12300
rect 12290 -12370 12330 -12300
rect 12400 -12370 12440 -12300
rect 12510 -12370 12550 -12300
rect 12620 -12370 12690 -12300
rect 11090 -12410 12690 -12370
rect 11090 -12480 11120 -12410
rect 11190 -12480 11230 -12410
rect 11300 -12480 11340 -12410
rect 11410 -12480 11450 -12410
rect 11520 -12480 11560 -12410
rect 11630 -12480 11670 -12410
rect 11740 -12480 11780 -12410
rect 11850 -12480 11890 -12410
rect 11960 -12480 12000 -12410
rect 12070 -12480 12110 -12410
rect 12180 -12480 12220 -12410
rect 12290 -12480 12330 -12410
rect 12400 -12480 12440 -12410
rect 12510 -12480 12550 -12410
rect 12620 -12480 12690 -12410
rect 11090 -12510 12690 -12480
rect 6980 -13250 7310 -13220
rect 6980 -13310 7010 -13250
rect 7070 -13310 7110 -13250
rect 7170 -13310 7210 -13250
rect 7270 -13310 7310 -13250
rect 6980 -13340 7310 -13310
rect 6980 -13400 7010 -13340
rect 7070 -13400 7110 -13340
rect 7170 -13400 7210 -13340
rect 7270 -13400 7310 -13340
rect 6980 -13430 7310 -13400
rect 6980 -13490 7010 -13430
rect 7070 -13490 7110 -13430
rect 7170 -13490 7210 -13430
rect 7270 -13490 7310 -13430
rect 6980 -13530 7310 -13490
rect 6980 -13590 7010 -13530
rect 7070 -13590 7110 -13530
rect 7170 -13590 7210 -13530
rect 7270 -13590 7310 -13530
rect 6980 -13620 7310 -13590
rect 6980 -13680 7010 -13620
rect 7070 -13680 7110 -13620
rect 7170 -13680 7210 -13620
rect 7270 -13680 7310 -13620
rect 6980 -13710 7310 -13680
rect 6980 -13770 7010 -13710
rect 7070 -13770 7110 -13710
rect 7170 -13770 7210 -13710
rect 7270 -13770 7310 -13710
rect 6980 -13800 7310 -13770
rect 7590 -13250 7920 -13220
rect 7590 -13310 7630 -13250
rect 7690 -13310 7730 -13250
rect 7790 -13310 7830 -13250
rect 7890 -13310 7920 -13250
rect 7590 -13340 7920 -13310
rect 7590 -13400 7630 -13340
rect 7690 -13400 7730 -13340
rect 7790 -13400 7830 -13340
rect 7890 -13400 7920 -13340
rect 7590 -13430 7920 -13400
rect 7590 -13490 7630 -13430
rect 7690 -13490 7730 -13430
rect 7790 -13490 7830 -13430
rect 7890 -13490 7920 -13430
rect 7590 -13530 7920 -13490
rect 7590 -13590 7630 -13530
rect 7690 -13590 7730 -13530
rect 7790 -13590 7830 -13530
rect 7890 -13590 7920 -13530
rect 7590 -13620 7920 -13590
rect 7590 -13680 7630 -13620
rect 7690 -13680 7730 -13620
rect 7790 -13680 7830 -13620
rect 7890 -13680 7920 -13620
rect 7590 -13710 7920 -13680
rect 7590 -13770 7630 -13710
rect 7690 -13770 7730 -13710
rect 7790 -13770 7830 -13710
rect 7890 -13770 7920 -13710
rect 7590 -13800 7920 -13770
rect 21610 -14020 21930 -13990
rect 21610 -14090 21630 -14020
rect 21700 -14090 21730 -14020
rect 21800 -14090 21830 -14020
rect 21900 -14090 21930 -14020
rect 21610 -14120 21930 -14090
rect 21610 -14190 21630 -14120
rect 21700 -14190 21730 -14120
rect 21800 -14190 21830 -14120
rect 21900 -14190 21930 -14120
rect 21610 -14220 21930 -14190
rect 21610 -14290 21630 -14220
rect 21700 -14290 21730 -14220
rect 21800 -14290 21830 -14220
rect 21900 -14290 21930 -14220
rect 21610 -14310 21930 -14290
rect 22900 -14870 23220 -14840
rect 22900 -14940 22920 -14870
rect 22990 -14940 23020 -14870
rect 23090 -14940 23120 -14870
rect 23190 -14940 23220 -14870
rect 22900 -14970 23220 -14940
rect 22900 -15040 22920 -14970
rect 22990 -15040 23020 -14970
rect 23090 -15040 23120 -14970
rect 23190 -15040 23220 -14970
rect 22900 -15070 23220 -15040
rect 22900 -15140 22920 -15070
rect 22990 -15140 23020 -15070
rect 23090 -15140 23120 -15070
rect 23190 -15140 23220 -15070
rect 22900 -15160 23220 -15140
rect 5010 -17100 5330 -17070
rect 5010 -17160 5040 -17100
rect 5100 -17160 5140 -17100
rect 5200 -17160 5240 -17100
rect 5300 -17160 5330 -17100
rect 5010 -17200 5330 -17160
rect 5010 -17260 5040 -17200
rect 5100 -17260 5140 -17200
rect 5200 -17260 5240 -17200
rect 5300 -17260 5330 -17200
rect 5010 -17300 5330 -17260
rect 5010 -17360 5040 -17300
rect 5100 -17360 5140 -17300
rect 5200 -17360 5240 -17300
rect 5300 -17360 5330 -17300
rect 5010 -17380 5330 -17360
rect 9570 -17100 9890 -17070
rect 9570 -17160 9600 -17100
rect 9660 -17160 9700 -17100
rect 9760 -17160 9800 -17100
rect 9860 -17160 9890 -17100
rect 9570 -17200 9890 -17160
rect 9570 -17260 9600 -17200
rect 9660 -17260 9700 -17200
rect 9760 -17260 9800 -17200
rect 9860 -17260 9890 -17200
rect 9570 -17300 9890 -17260
rect 9570 -17360 9600 -17300
rect 9660 -17360 9700 -17300
rect 9760 -17360 9800 -17300
rect 9860 -17360 9890 -17300
rect 9570 -17380 9890 -17360
rect 7210 -17600 7650 -17580
rect 7210 -17670 7230 -17600
rect 7300 -17670 7340 -17600
rect 7410 -17670 7450 -17600
rect 7520 -17670 7560 -17600
rect 7630 -17670 7650 -17600
rect 7210 -17710 7650 -17670
rect 7210 -17780 7230 -17710
rect 7300 -17780 7340 -17710
rect 7410 -17780 7450 -17710
rect 7520 -17780 7560 -17710
rect 7630 -17780 7650 -17710
rect 7210 -17820 7650 -17780
rect 7210 -17890 7230 -17820
rect 7300 -17890 7340 -17820
rect 7410 -17890 7450 -17820
rect 7520 -17890 7560 -17820
rect 7630 -17890 7650 -17820
rect 7210 -17930 7650 -17890
rect 7210 -18000 7230 -17930
rect 7300 -18000 7340 -17930
rect 7410 -18000 7450 -17930
rect 7520 -18000 7560 -17930
rect 7630 -18000 7650 -17930
rect 7210 -18020 7650 -18000
rect 21610 -20100 21930 -20070
rect 21610 -20170 21630 -20100
rect 21700 -20170 21730 -20100
rect 21800 -20170 21830 -20100
rect 21900 -20170 21930 -20100
rect 21610 -20200 21930 -20170
rect 21610 -20270 21630 -20200
rect 21700 -20270 21730 -20200
rect 21800 -20270 21830 -20200
rect 21900 -20270 21930 -20200
rect 21610 -20300 21930 -20270
rect 21610 -20370 21630 -20300
rect 21700 -20370 21730 -20300
rect 21800 -20370 21830 -20300
rect 21900 -20370 21930 -20300
rect 21610 -20390 21930 -20370
rect 22680 -20730 23000 -20700
rect 22680 -20800 22700 -20730
rect 22770 -20800 22800 -20730
rect 22870 -20800 22900 -20730
rect 22970 -20800 23000 -20730
rect 22680 -20830 23000 -20800
rect 22680 -20900 22700 -20830
rect 22770 -20900 22800 -20830
rect 22870 -20900 22900 -20830
rect 22970 -20900 23000 -20830
rect 22680 -20930 23000 -20900
rect 22680 -21000 22700 -20930
rect 22770 -21000 22800 -20930
rect 22870 -21000 22900 -20930
rect 22970 -21000 23000 -20930
rect 22680 -21020 23000 -21000
rect 2210 -22660 3810 -22630
rect 2210 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3160 -22660
rect 3230 -22730 3270 -22660
rect 3340 -22730 3380 -22660
rect 3450 -22730 3490 -22660
rect 3560 -22730 3600 -22660
rect 3670 -22730 3710 -22660
rect 3780 -22730 3810 -22660
rect 2210 -22770 3810 -22730
rect 2210 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3160 -22770
rect 3230 -22840 3270 -22770
rect 3340 -22840 3380 -22770
rect 3450 -22840 3490 -22770
rect 3560 -22840 3600 -22770
rect 3670 -22840 3710 -22770
rect 3780 -22840 3810 -22770
rect 2210 -22890 3810 -22840
rect 11090 -22660 12690 -22630
rect 11090 -22730 11160 -22660
rect 11230 -22730 11270 -22660
rect 11340 -22730 11380 -22660
rect 11450 -22730 11490 -22660
rect 11560 -22730 11600 -22660
rect 11670 -22730 11710 -22660
rect 11780 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12690 -22660
rect 11090 -22770 12690 -22730
rect 11090 -22840 11160 -22770
rect 11230 -22840 11270 -22770
rect 11340 -22840 11380 -22770
rect 11450 -22840 11490 -22770
rect 11560 -22840 11600 -22770
rect 11670 -22840 11710 -22770
rect 11780 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12690 -22770
rect 11090 -22890 12690 -22840
<< via2 >>
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 25890 7140 25960 7210
rect 26000 7140 26070 7210
rect 26110 7140 26180 7210
rect 26220 7140 26290 7210
rect 25890 7030 25960 7100
rect 26000 7030 26070 7100
rect 26110 7030 26180 7100
rect 26220 7030 26290 7100
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 30740 6230 30810 6300
rect 30850 6230 30920 6300
rect 30740 6100 30810 6170
rect 30850 6100 30920 6170
rect 30740 5970 30810 6040
rect 30850 5970 30920 6040
rect 21820 5600 21890 5670
rect 21930 5600 22000 5670
rect 21820 5490 21890 5560
rect 21930 5490 22000 5560
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect 21820 5380 21890 5450
rect 21930 5380 22000 5450
rect 21820 5270 21890 5340
rect 21930 5270 22000 5340
rect 21820 5160 21890 5230
rect 21930 5160 22000 5230
rect 21820 5050 21890 5120
rect 21930 5050 22000 5120
rect 21820 4940 21890 5010
rect 21930 4940 22000 5010
rect 21820 4830 21890 4900
rect 21930 4830 22000 4900
rect 7590 4700 7650 4760
rect 7690 4700 7750 4760
rect 7790 4700 7850 4760
rect 21820 4720 21890 4790
rect 21930 4720 22000 4790
rect 21820 4610 21890 4680
rect 21930 4610 22000 4680
rect -1710 4510 -1640 4580
rect -1710 4400 -1640 4470
rect -1710 4290 -1640 4360
rect -1710 4180 -1640 4250
rect 6700 4520 6760 4580
rect 6700 4400 6760 4460
rect 6700 4280 6760 4340
rect 6700 4160 6760 4220
rect 16420 4510 16490 4580
rect 21820 4500 21890 4570
rect 21930 4500 22000 4570
rect 16420 4400 16490 4470
rect 16420 4290 16490 4360
rect 16420 4180 16490 4250
rect 7050 3180 7110 3240
rect 7150 3180 7210 3240
rect 7250 3180 7310 3240
rect 7050 3080 7110 3140
rect 7150 3080 7210 3140
rect 7250 3080 7310 3140
rect 7050 2980 7110 3040
rect 7150 2980 7210 3040
rect 7250 2980 7310 3040
rect 24720 3290 24790 3360
rect 24830 3290 24900 3360
rect 24940 3290 25010 3360
rect 24720 3180 24790 3250
rect 24830 3180 24900 3250
rect 24940 3180 25010 3250
rect 24720 3070 24790 3140
rect 24830 3070 24900 3140
rect 24940 3070 25010 3140
rect 4770 2830 4830 2890
rect 4870 2830 4930 2890
rect 4970 2830 5030 2890
rect 4770 2730 4830 2790
rect 4870 2730 4930 2790
rect 4970 2730 5030 2790
rect 4770 2630 4830 2690
rect 4870 2630 4930 2690
rect 4970 2630 5030 2690
rect 9870 2830 9930 2890
rect 9970 2830 10030 2890
rect 10070 2830 10130 2890
rect 9870 2730 9930 2790
rect 9970 2730 10030 2790
rect 10070 2730 10130 2790
rect 9870 2630 9930 2690
rect 9970 2630 10030 2690
rect 10070 2630 10130 2690
rect 22470 2530 22540 2600
rect 22580 2530 22650 2600
rect 22690 2530 22760 2600
rect 22800 2530 22870 2600
rect 22470 2420 22540 2490
rect 22580 2420 22650 2490
rect 22690 2420 22760 2490
rect 22800 2420 22870 2490
rect 26950 2530 27020 2600
rect 27060 2530 27130 2600
rect 27170 2530 27240 2600
rect 27280 2530 27350 2600
rect 26950 2420 27020 2490
rect 27060 2420 27130 2490
rect 27170 2420 27240 2490
rect 27280 2420 27350 2490
rect -300 -210 -230 -140
rect -190 -210 -120 -140
rect -80 -210 -10 -140
rect 30 -210 100 -140
rect -300 -340 -230 -270
rect -190 -340 -120 -270
rect -80 -340 -10 -270
rect 30 -340 100 -270
rect 14600 1090 14670 1160
rect 14700 1090 14770 1160
rect 14810 1090 14880 1160
rect 14600 980 14670 1050
rect 14700 980 14770 1050
rect 14810 980 14880 1050
rect 14600 870 14670 940
rect 14700 870 14770 940
rect 14810 870 14880 940
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect 25890 850 25960 920
rect 26000 850 26070 920
rect 26110 850 26180 920
rect 26220 850 26290 920
rect 25890 740 25960 810
rect 26000 740 26070 810
rect 26110 740 26180 810
rect 26220 740 26290 810
rect 30740 -70 30810 0
rect 30850 -70 30920 0
rect 14660 -210 14730 -140
rect 14770 -210 14840 -140
rect 14880 -210 14950 -140
rect 14990 -210 15060 -140
rect 14660 -340 14730 -270
rect 14770 -340 14840 -270
rect 14880 -340 14950 -270
rect 14990 -340 15060 -270
rect 30740 -200 30810 -130
rect 30850 -200 30920 -130
rect 30740 -330 30810 -260
rect 30850 -330 30920 -260
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 21820 -920 21890 -850
rect 21930 -920 22000 -850
rect 21820 -1030 21890 -960
rect 21930 -1030 22000 -960
rect 21820 -1140 21890 -1070
rect 21930 -1140 22000 -1070
rect 21820 -1250 21890 -1180
rect 21930 -1250 22000 -1180
rect 21820 -1360 21890 -1290
rect 21930 -1360 22000 -1290
rect 21820 -1470 21890 -1400
rect 21930 -1470 22000 -1400
rect 21820 -1580 21890 -1510
rect 21930 -1580 22000 -1510
rect 21820 -1690 21890 -1620
rect 21930 -1690 22000 -1620
rect 21820 -1800 21890 -1730
rect 21930 -1800 22000 -1730
rect 21820 -1910 21890 -1840
rect 21930 -1910 22000 -1840
rect 21820 -2020 21890 -1950
rect 21930 -2020 22000 -1950
rect 24740 -3120 24810 -3050
rect 24850 -3120 24920 -3050
rect 24960 -3120 25030 -3050
rect 24740 -3230 24810 -3160
rect 24850 -3230 24920 -3160
rect 24960 -3230 25030 -3160
rect 24740 -3340 24810 -3270
rect 24850 -3340 24920 -3270
rect 24960 -3340 25030 -3270
rect 22470 -3760 22540 -3690
rect 22580 -3760 22650 -3690
rect 22690 -3760 22760 -3690
rect 22800 -3760 22870 -3690
rect 7310 -3950 7380 -3880
rect 7420 -3950 7490 -3880
rect 7530 -3950 7600 -3880
rect 22470 -3870 22540 -3800
rect 22580 -3870 22650 -3800
rect 22690 -3870 22760 -3800
rect 22800 -3870 22870 -3800
rect 26950 -3760 27020 -3690
rect 27060 -3760 27130 -3690
rect 27170 -3760 27240 -3690
rect 27280 -3760 27350 -3690
rect 26950 -3870 27020 -3800
rect 27060 -3870 27130 -3800
rect 27170 -3870 27240 -3800
rect 27280 -3870 27350 -3800
rect 7310 -4060 7380 -3990
rect 7420 -4060 7490 -3990
rect 7530 -4060 7600 -3990
rect 7310 -4170 7380 -4100
rect 7420 -4170 7490 -4100
rect 7530 -4170 7600 -4100
rect -1330 -4420 -1260 -4350
rect -1220 -4420 -1150 -4350
rect -1110 -4420 -1040 -4350
rect -1000 -4420 -930 -4350
rect -1330 -4530 -1260 -4460
rect -1220 -4530 -1150 -4460
rect -1110 -4530 -1040 -4460
rect -1000 -4530 -930 -4460
rect -560 -4360 -490 -4290
rect -450 -4360 -380 -4290
rect -340 -4360 -270 -4290
rect -230 -4360 -160 -4290
rect -560 -4470 -490 -4400
rect -450 -4470 -380 -4400
rect -340 -4470 -270 -4400
rect -230 -4470 -160 -4400
rect 14940 -4360 15010 -4290
rect 15050 -4360 15120 -4290
rect 15160 -4360 15230 -4290
rect 15270 -4360 15340 -4290
rect 14940 -4470 15010 -4400
rect 15050 -4470 15120 -4400
rect 15160 -4470 15230 -4400
rect 15270 -4470 15340 -4400
rect 15710 -4420 15780 -4350
rect 15820 -4420 15890 -4350
rect 15930 -4420 16000 -4350
rect 16040 -4420 16110 -4350
rect 15710 -4530 15780 -4460
rect 15820 -4530 15890 -4460
rect 15930 -4530 16000 -4460
rect 16040 -4530 16110 -4460
rect -1710 -6590 -1640 -6520
rect -1710 -6700 -1640 -6630
rect 7050 -6520 7110 -6460
rect 7150 -6520 7210 -6460
rect 7250 -6520 7310 -6460
rect 7050 -6620 7110 -6560
rect 7150 -6620 7210 -6560
rect 7250 -6620 7310 -6560
rect -1710 -6810 -1640 -6740
rect -1710 -6920 -1640 -6850
rect 4770 -6730 4830 -6670
rect 4870 -6730 4930 -6670
rect 4970 -6730 5030 -6670
rect 4770 -6830 4830 -6770
rect 4870 -6830 4930 -6770
rect 4970 -6830 5030 -6770
rect 7050 -6720 7110 -6660
rect 7150 -6720 7210 -6660
rect 7250 -6720 7310 -6660
rect 7050 -6820 7110 -6760
rect 7150 -6820 7210 -6760
rect 7250 -6820 7310 -6760
rect 7590 -6520 7650 -6460
rect 7690 -6520 7750 -6460
rect 7790 -6520 7850 -6460
rect 7590 -6620 7650 -6560
rect 7690 -6620 7750 -6560
rect 7790 -6620 7850 -6560
rect 16420 -6590 16490 -6520
rect 7590 -6720 7650 -6660
rect 7690 -6720 7750 -6660
rect 7790 -6720 7850 -6660
rect 7590 -6820 7650 -6760
rect 7690 -6820 7750 -6760
rect 7790 -6820 7850 -6760
rect 9870 -6730 9930 -6670
rect 9970 -6730 10030 -6670
rect 10070 -6730 10130 -6670
rect 9870 -6830 9930 -6770
rect 9970 -6830 10030 -6770
rect 10070 -6830 10130 -6770
rect 4770 -6930 4830 -6870
rect 4870 -6930 4930 -6870
rect 4970 -6930 5030 -6870
rect 9870 -6930 9930 -6870
rect 9970 -6930 10030 -6870
rect 10070 -6930 10130 -6870
rect 16420 -6700 16490 -6630
rect 16420 -6810 16490 -6740
rect 16420 -6920 16490 -6850
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect 21630 -8430 21700 -8360
rect 21730 -8430 21800 -8360
rect 21830 -8430 21900 -8360
rect 21630 -8530 21700 -8460
rect 21730 -8530 21800 -8460
rect 21830 -8530 21900 -8460
rect 21630 -8630 21700 -8560
rect 21730 -8630 21800 -8560
rect 21830 -8630 21900 -8560
rect 22650 -9080 22720 -9010
rect 22750 -9080 22820 -9010
rect 22850 -9080 22920 -9010
rect 22650 -9180 22720 -9110
rect 22750 -9180 22820 -9110
rect 22850 -9180 22920 -9110
rect 22650 -9280 22720 -9210
rect 22750 -9280 22820 -9210
rect 22850 -9280 22920 -9210
rect -240 -9730 -170 -9660
rect -130 -9730 -60 -9660
rect -20 -9730 50 -9660
rect 90 -9730 160 -9660
rect -240 -9860 -170 -9790
rect -130 -9860 -60 -9790
rect -20 -9860 50 -9790
rect 90 -9860 160 -9790
rect 14720 -9730 14790 -9660
rect 14830 -9730 14900 -9660
rect 14940 -9730 15010 -9660
rect 15050 -9730 15120 -9660
rect 14720 -9860 14790 -9790
rect 14830 -9860 14900 -9790
rect 14940 -9860 15010 -9790
rect 15050 -9860 15120 -9790
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 2240 -12370 2310 -12300
rect 2350 -12370 2420 -12300
rect 2460 -12370 2530 -12300
rect 2570 -12370 2640 -12300
rect 2680 -12370 2750 -12300
rect 2790 -12370 2860 -12300
rect 2900 -12370 2970 -12300
rect 3010 -12370 3080 -12300
rect 3120 -12370 3190 -12300
rect 3230 -12370 3300 -12300
rect 3340 -12370 3410 -12300
rect 3450 -12370 3520 -12300
rect 3560 -12370 3630 -12300
rect 3670 -12370 3740 -12300
rect 2240 -12480 2310 -12410
rect 2350 -12480 2420 -12410
rect 2460 -12480 2530 -12410
rect 2570 -12480 2640 -12410
rect 2680 -12480 2750 -12410
rect 2790 -12480 2860 -12410
rect 2900 -12480 2970 -12410
rect 3010 -12480 3080 -12410
rect 3120 -12480 3190 -12410
rect 3230 -12480 3300 -12410
rect 3340 -12480 3410 -12410
rect 3450 -12480 3520 -12410
rect 3560 -12480 3630 -12410
rect 3670 -12480 3740 -12410
rect 11120 -12370 11190 -12300
rect 11230 -12370 11300 -12300
rect 11340 -12370 11410 -12300
rect 11450 -12370 11520 -12300
rect 11560 -12370 11630 -12300
rect 11670 -12370 11740 -12300
rect 11780 -12370 11850 -12300
rect 11890 -12370 11960 -12300
rect 12000 -12370 12070 -12300
rect 12110 -12370 12180 -12300
rect 12220 -12370 12290 -12300
rect 12330 -12370 12400 -12300
rect 12440 -12370 12510 -12300
rect 12550 -12370 12620 -12300
rect 11120 -12480 11190 -12410
rect 11230 -12480 11300 -12410
rect 11340 -12480 11410 -12410
rect 11450 -12480 11520 -12410
rect 11560 -12480 11630 -12410
rect 11670 -12480 11740 -12410
rect 11780 -12480 11850 -12410
rect 11890 -12480 11960 -12410
rect 12000 -12480 12070 -12410
rect 12110 -12480 12180 -12410
rect 12220 -12480 12290 -12410
rect 12330 -12480 12400 -12410
rect 12440 -12480 12510 -12410
rect 12550 -12480 12620 -12410
rect 7010 -13310 7070 -13250
rect 7110 -13310 7170 -13250
rect 7210 -13310 7270 -13250
rect 7010 -13400 7070 -13340
rect 7110 -13400 7170 -13340
rect 7210 -13400 7270 -13340
rect 7010 -13490 7070 -13430
rect 7110 -13490 7170 -13430
rect 7210 -13490 7270 -13430
rect 7010 -13590 7070 -13530
rect 7110 -13590 7170 -13530
rect 7210 -13590 7270 -13530
rect 7010 -13680 7070 -13620
rect 7110 -13680 7170 -13620
rect 7210 -13680 7270 -13620
rect 7010 -13770 7070 -13710
rect 7110 -13770 7170 -13710
rect 7210 -13770 7270 -13710
rect 7630 -13310 7690 -13250
rect 7730 -13310 7790 -13250
rect 7830 -13310 7890 -13250
rect 7630 -13400 7690 -13340
rect 7730 -13400 7790 -13340
rect 7830 -13400 7890 -13340
rect 7630 -13490 7690 -13430
rect 7730 -13490 7790 -13430
rect 7830 -13490 7890 -13430
rect 7630 -13590 7690 -13530
rect 7730 -13590 7790 -13530
rect 7830 -13590 7890 -13530
rect 7630 -13680 7690 -13620
rect 7730 -13680 7790 -13620
rect 7830 -13680 7890 -13620
rect 7630 -13770 7690 -13710
rect 7730 -13770 7790 -13710
rect 7830 -13770 7890 -13710
rect 21630 -14090 21700 -14020
rect 21730 -14090 21800 -14020
rect 21830 -14090 21900 -14020
rect 21630 -14190 21700 -14120
rect 21730 -14190 21800 -14120
rect 21830 -14190 21900 -14120
rect 21630 -14290 21700 -14220
rect 21730 -14290 21800 -14220
rect 21830 -14290 21900 -14220
rect 22920 -14940 22990 -14870
rect 23020 -14940 23090 -14870
rect 23120 -14940 23190 -14870
rect 22920 -15040 22990 -14970
rect 23020 -15040 23090 -14970
rect 23120 -15040 23190 -14970
rect 22920 -15140 22990 -15070
rect 23020 -15140 23090 -15070
rect 23120 -15140 23190 -15070
rect 5040 -17160 5100 -17100
rect 5140 -17160 5200 -17100
rect 5240 -17160 5300 -17100
rect 5040 -17260 5100 -17200
rect 5140 -17260 5200 -17200
rect 5240 -17260 5300 -17200
rect 5040 -17360 5100 -17300
rect 5140 -17360 5200 -17300
rect 5240 -17360 5300 -17300
rect 9600 -17160 9660 -17100
rect 9700 -17160 9760 -17100
rect 9800 -17160 9860 -17100
rect 9600 -17260 9660 -17200
rect 9700 -17260 9760 -17200
rect 9800 -17260 9860 -17200
rect 9600 -17360 9660 -17300
rect 9700 -17360 9760 -17300
rect 9800 -17360 9860 -17300
rect 7230 -17670 7300 -17600
rect 7340 -17670 7410 -17600
rect 7450 -17670 7520 -17600
rect 7560 -17670 7630 -17600
rect 7230 -17780 7300 -17710
rect 7340 -17780 7410 -17710
rect 7450 -17780 7520 -17710
rect 7560 -17780 7630 -17710
rect 7230 -17890 7300 -17820
rect 7340 -17890 7410 -17820
rect 7450 -17890 7520 -17820
rect 7560 -17890 7630 -17820
rect 7230 -18000 7300 -17930
rect 7340 -18000 7410 -17930
rect 7450 -18000 7520 -17930
rect 7560 -18000 7630 -17930
rect 21630 -20170 21700 -20100
rect 21730 -20170 21800 -20100
rect 21830 -20170 21900 -20100
rect 21630 -20270 21700 -20200
rect 21730 -20270 21800 -20200
rect 21830 -20270 21900 -20200
rect 21630 -20370 21700 -20300
rect 21730 -20370 21800 -20300
rect 21830 -20370 21900 -20300
rect 22700 -20800 22770 -20730
rect 22800 -20800 22870 -20730
rect 22900 -20800 22970 -20730
rect 22700 -20900 22770 -20830
rect 22800 -20900 22870 -20830
rect 22900 -20900 22970 -20830
rect 22700 -21000 22770 -20930
rect 22800 -21000 22870 -20930
rect 22900 -21000 22970 -20930
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 3160 -22730 3230 -22660
rect 3270 -22730 3340 -22660
rect 3380 -22730 3450 -22660
rect 3490 -22730 3560 -22660
rect 3600 -22730 3670 -22660
rect 3710 -22730 3780 -22660
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 3160 -22840 3230 -22770
rect 3270 -22840 3340 -22770
rect 3380 -22840 3450 -22770
rect 3490 -22840 3560 -22770
rect 3600 -22840 3670 -22770
rect 3710 -22840 3780 -22770
rect 11160 -22730 11230 -22660
rect 11270 -22730 11340 -22660
rect 11380 -22730 11450 -22660
rect 11490 -22730 11560 -22660
rect 11600 -22730 11670 -22660
rect 11710 -22730 11780 -22660
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 11160 -22840 11230 -22770
rect 11270 -22840 11340 -22770
rect 11380 -22840 11450 -22770
rect 11490 -22840 11560 -22770
rect 11600 -22840 11670 -22770
rect 11710 -22840 11780 -22770
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
<< metal3 >>
rect -5020 21580 7290 21640
rect -5020 21510 -4730 21580
rect -4660 21510 -4640 21580
rect -4570 21510 -4550 21580
rect -4480 21510 -4460 21580
rect -4390 21510 -4370 21580
rect -4300 21510 -4280 21580
rect -4210 21510 -4190 21580
rect -4120 21510 -4100 21580
rect -4030 21510 -4010 21580
rect -3940 21510 -3920 21580
rect -3850 21510 -3830 21580
rect -3760 21510 -3740 21580
rect -3670 21510 -3650 21580
rect -3580 21510 -3560 21580
rect -3490 21510 -3470 21580
rect -3400 21510 -3380 21580
rect -3310 21510 -3290 21580
rect -3220 21510 -3200 21580
rect -3130 21510 -3110 21580
rect -3040 21510 -3020 21580
rect -2950 21510 -2930 21580
rect -2860 21510 -2840 21580
rect -2770 21510 -2750 21580
rect -2680 21510 -2660 21580
rect -2590 21510 -2570 21580
rect -2500 21510 -2480 21580
rect -2410 21510 -2390 21580
rect -2320 21510 -2300 21580
rect -2230 21510 -2210 21580
rect -2140 21510 -2120 21580
rect -2050 21510 -2030 21580
rect -1960 21510 -1940 21580
rect -1870 21510 -1850 21580
rect -1780 21510 -1720 21580
rect -1650 21510 -1630 21580
rect -1560 21510 -1540 21580
rect -1470 21510 -1450 21580
rect -1380 21510 -1360 21580
rect -1290 21510 -1270 21580
rect -1200 21510 -1180 21580
rect -1110 21510 -1090 21580
rect -1020 21510 -1000 21580
rect -930 21510 -910 21580
rect -840 21510 -820 21580
rect -750 21510 -730 21580
rect -660 21510 -640 21580
rect -570 21510 -550 21580
rect -480 21510 -460 21580
rect -390 21510 -370 21580
rect -300 21510 -280 21580
rect -210 21510 -190 21580
rect -120 21510 -100 21580
rect -30 21510 -10 21580
rect 60 21510 80 21580
rect 150 21510 170 21580
rect 240 21510 260 21580
rect 330 21510 350 21580
rect 420 21510 440 21580
rect 510 21510 530 21580
rect 600 21510 620 21580
rect 690 21510 710 21580
rect 780 21510 800 21580
rect 870 21510 890 21580
rect 960 21510 980 21580
rect 1050 21510 1070 21580
rect 1140 21510 1160 21580
rect 1230 21510 1290 21580
rect 1360 21510 1380 21580
rect 1450 21510 1470 21580
rect 1540 21510 1560 21580
rect 1630 21510 1650 21580
rect 1720 21510 1740 21580
rect 1810 21510 1830 21580
rect 1900 21510 1920 21580
rect 1990 21510 2010 21580
rect 2080 21510 2100 21580
rect 2170 21510 2190 21580
rect 2260 21510 2280 21580
rect 2350 21510 2370 21580
rect 2440 21510 2460 21580
rect 2530 21510 2550 21580
rect 2620 21510 2640 21580
rect 2710 21510 2730 21580
rect 2800 21510 2820 21580
rect 2890 21510 2910 21580
rect 2980 21510 3000 21580
rect 3070 21510 3090 21580
rect 3160 21510 3180 21580
rect 3250 21510 3270 21580
rect 3340 21510 3360 21580
rect 3430 21510 3450 21580
rect 3520 21510 3540 21580
rect 3610 21510 3630 21580
rect 3700 21510 3720 21580
rect 3790 21510 3810 21580
rect 3880 21510 3900 21580
rect 3970 21510 3990 21580
rect 4060 21510 4080 21580
rect 4150 21510 4170 21580
rect 4240 21510 4300 21580
rect 4370 21510 4390 21580
rect 4460 21510 4480 21580
rect 4550 21510 4570 21580
rect 4640 21510 4660 21580
rect 4730 21510 4750 21580
rect 4820 21510 4840 21580
rect 4910 21510 4930 21580
rect 5000 21510 5020 21580
rect 5090 21510 5110 21580
rect 5180 21510 5200 21580
rect 5270 21510 5290 21580
rect 5360 21510 5380 21580
rect 5450 21510 5470 21580
rect 5540 21510 5560 21580
rect 5630 21510 5650 21580
rect 5720 21510 5740 21580
rect 5810 21510 5830 21580
rect 5900 21510 5920 21580
rect 5990 21510 6010 21580
rect 6080 21510 6100 21580
rect 6170 21510 6190 21580
rect 6260 21510 6280 21580
rect 6350 21510 6370 21580
rect 6440 21510 6460 21580
rect 6530 21510 6550 21580
rect 6620 21510 6640 21580
rect 6710 21510 6730 21580
rect 6800 21510 6820 21580
rect 6890 21510 6910 21580
rect 6980 21510 7000 21580
rect 7070 21510 7090 21580
rect 7160 21510 7180 21580
rect 7250 21510 7290 21580
rect -5020 21490 7290 21510
rect -5020 21420 -4730 21490
rect -4660 21420 -4640 21490
rect -4570 21420 -4550 21490
rect -4480 21420 -4460 21490
rect -4390 21420 -4370 21490
rect -4300 21420 -4280 21490
rect -4210 21420 -4190 21490
rect -4120 21420 -4100 21490
rect -4030 21420 -4010 21490
rect -3940 21420 -3920 21490
rect -3850 21420 -3830 21490
rect -3760 21420 -3740 21490
rect -3670 21420 -3650 21490
rect -3580 21420 -3560 21490
rect -3490 21420 -3470 21490
rect -3400 21420 -3380 21490
rect -3310 21420 -3290 21490
rect -3220 21420 -3200 21490
rect -3130 21420 -3110 21490
rect -3040 21420 -3020 21490
rect -2950 21420 -2930 21490
rect -2860 21420 -2840 21490
rect -2770 21420 -2750 21490
rect -2680 21420 -2660 21490
rect -2590 21420 -2570 21490
rect -2500 21420 -2480 21490
rect -2410 21420 -2390 21490
rect -2320 21420 -2300 21490
rect -2230 21420 -2210 21490
rect -2140 21420 -2120 21490
rect -2050 21420 -2030 21490
rect -1960 21420 -1940 21490
rect -1870 21420 -1850 21490
rect -1780 21420 -1720 21490
rect -1650 21420 -1630 21490
rect -1560 21420 -1540 21490
rect -1470 21420 -1450 21490
rect -1380 21420 -1360 21490
rect -1290 21420 -1270 21490
rect -1200 21420 -1180 21490
rect -1110 21420 -1090 21490
rect -1020 21420 -1000 21490
rect -930 21420 -910 21490
rect -840 21420 -820 21490
rect -750 21420 -730 21490
rect -660 21420 -640 21490
rect -570 21420 -550 21490
rect -480 21420 -460 21490
rect -390 21420 -370 21490
rect -300 21420 -280 21490
rect -210 21420 -190 21490
rect -120 21420 -100 21490
rect -30 21420 -10 21490
rect 60 21420 80 21490
rect 150 21420 170 21490
rect 240 21420 260 21490
rect 330 21420 350 21490
rect 420 21420 440 21490
rect 510 21420 530 21490
rect 600 21420 620 21490
rect 690 21420 710 21490
rect 780 21420 800 21490
rect 870 21420 890 21490
rect 960 21420 980 21490
rect 1050 21420 1070 21490
rect 1140 21420 1160 21490
rect 1230 21420 1290 21490
rect 1360 21420 1380 21490
rect 1450 21420 1470 21490
rect 1540 21420 1560 21490
rect 1630 21420 1650 21490
rect 1720 21420 1740 21490
rect 1810 21420 1830 21490
rect 1900 21420 1920 21490
rect 1990 21420 2010 21490
rect 2080 21420 2100 21490
rect 2170 21420 2190 21490
rect 2260 21420 2280 21490
rect 2350 21420 2370 21490
rect 2440 21420 2460 21490
rect 2530 21420 2550 21490
rect 2620 21420 2640 21490
rect 2710 21420 2730 21490
rect 2800 21420 2820 21490
rect 2890 21420 2910 21490
rect 2980 21420 3000 21490
rect 3070 21420 3090 21490
rect 3160 21420 3180 21490
rect 3250 21420 3270 21490
rect 3340 21420 3360 21490
rect 3430 21420 3450 21490
rect 3520 21420 3540 21490
rect 3610 21420 3630 21490
rect 3700 21420 3720 21490
rect 3790 21420 3810 21490
rect 3880 21420 3900 21490
rect 3970 21420 3990 21490
rect 4060 21420 4080 21490
rect 4150 21420 4170 21490
rect 4240 21420 4300 21490
rect 4370 21420 4390 21490
rect 4460 21420 4480 21490
rect 4550 21420 4570 21490
rect 4640 21420 4660 21490
rect 4730 21420 4750 21490
rect 4820 21420 4840 21490
rect 4910 21420 4930 21490
rect 5000 21420 5020 21490
rect 5090 21420 5110 21490
rect 5180 21420 5200 21490
rect 5270 21420 5290 21490
rect 5360 21420 5380 21490
rect 5450 21420 5470 21490
rect 5540 21420 5560 21490
rect 5630 21420 5650 21490
rect 5720 21420 5740 21490
rect 5810 21420 5830 21490
rect 5900 21420 5920 21490
rect 5990 21420 6010 21490
rect 6080 21420 6100 21490
rect 6170 21420 6190 21490
rect 6260 21420 6280 21490
rect 6350 21420 6370 21490
rect 6440 21420 6460 21490
rect 6530 21420 6550 21490
rect 6620 21420 6640 21490
rect 6710 21420 6730 21490
rect 6800 21420 6820 21490
rect 6890 21420 6910 21490
rect 6980 21420 7000 21490
rect 7070 21420 7090 21490
rect 7160 21420 7180 21490
rect 7250 21420 7290 21490
rect -5020 21400 7290 21420
rect -5020 21330 -4730 21400
rect -4660 21330 -4640 21400
rect -4570 21330 -4550 21400
rect -4480 21330 -4460 21400
rect -4390 21330 -4370 21400
rect -4300 21330 -4280 21400
rect -4210 21330 -4190 21400
rect -4120 21330 -4100 21400
rect -4030 21330 -4010 21400
rect -3940 21330 -3920 21400
rect -3850 21330 -3830 21400
rect -3760 21330 -3740 21400
rect -3670 21330 -3650 21400
rect -3580 21330 -3560 21400
rect -3490 21330 -3470 21400
rect -3400 21330 -3380 21400
rect -3310 21330 -3290 21400
rect -3220 21330 -3200 21400
rect -3130 21330 -3110 21400
rect -3040 21330 -3020 21400
rect -2950 21330 -2930 21400
rect -2860 21330 -2840 21400
rect -2770 21330 -2750 21400
rect -2680 21330 -2660 21400
rect -2590 21330 -2570 21400
rect -2500 21330 -2480 21400
rect -2410 21330 -2390 21400
rect -2320 21330 -2300 21400
rect -2230 21330 -2210 21400
rect -2140 21330 -2120 21400
rect -2050 21330 -2030 21400
rect -1960 21330 -1940 21400
rect -1870 21330 -1850 21400
rect -1780 21330 -1720 21400
rect -1650 21330 -1630 21400
rect -1560 21330 -1540 21400
rect -1470 21330 -1450 21400
rect -1380 21330 -1360 21400
rect -1290 21330 -1270 21400
rect -1200 21330 -1180 21400
rect -1110 21330 -1090 21400
rect -1020 21330 -1000 21400
rect -930 21330 -910 21400
rect -840 21330 -820 21400
rect -750 21330 -730 21400
rect -660 21330 -640 21400
rect -570 21330 -550 21400
rect -480 21330 -460 21400
rect -390 21330 -370 21400
rect -300 21330 -280 21400
rect -210 21330 -190 21400
rect -120 21330 -100 21400
rect -30 21330 -10 21400
rect 60 21330 80 21400
rect 150 21330 170 21400
rect 240 21330 260 21400
rect 330 21330 350 21400
rect 420 21330 440 21400
rect 510 21330 530 21400
rect 600 21330 620 21400
rect 690 21330 710 21400
rect 780 21330 800 21400
rect 870 21330 890 21400
rect 960 21330 980 21400
rect 1050 21330 1070 21400
rect 1140 21330 1160 21400
rect 1230 21330 1290 21400
rect 1360 21330 1380 21400
rect 1450 21330 1470 21400
rect 1540 21330 1560 21400
rect 1630 21330 1650 21400
rect 1720 21330 1740 21400
rect 1810 21330 1830 21400
rect 1900 21330 1920 21400
rect 1990 21330 2010 21400
rect 2080 21330 2100 21400
rect 2170 21330 2190 21400
rect 2260 21330 2280 21400
rect 2350 21330 2370 21400
rect 2440 21330 2460 21400
rect 2530 21330 2550 21400
rect 2620 21330 2640 21400
rect 2710 21330 2730 21400
rect 2800 21330 2820 21400
rect 2890 21330 2910 21400
rect 2980 21330 3000 21400
rect 3070 21330 3090 21400
rect 3160 21330 3180 21400
rect 3250 21330 3270 21400
rect 3340 21330 3360 21400
rect 3430 21330 3450 21400
rect 3520 21330 3540 21400
rect 3610 21330 3630 21400
rect 3700 21330 3720 21400
rect 3790 21330 3810 21400
rect 3880 21330 3900 21400
rect 3970 21330 3990 21400
rect 4060 21330 4080 21400
rect 4150 21330 4170 21400
rect 4240 21330 4300 21400
rect 4370 21330 4390 21400
rect 4460 21330 4480 21400
rect 4550 21330 4570 21400
rect 4640 21330 4660 21400
rect 4730 21330 4750 21400
rect 4820 21330 4840 21400
rect 4910 21330 4930 21400
rect 5000 21330 5020 21400
rect 5090 21330 5110 21400
rect 5180 21330 5200 21400
rect 5270 21330 5290 21400
rect 5360 21330 5380 21400
rect 5450 21330 5470 21400
rect 5540 21330 5560 21400
rect 5630 21330 5650 21400
rect 5720 21330 5740 21400
rect 5810 21330 5830 21400
rect 5900 21330 5920 21400
rect 5990 21330 6010 21400
rect 6080 21330 6100 21400
rect 6170 21330 6190 21400
rect 6260 21330 6280 21400
rect 6350 21330 6370 21400
rect 6440 21330 6460 21400
rect 6530 21330 6550 21400
rect 6620 21330 6640 21400
rect 6710 21330 6730 21400
rect 6800 21330 6820 21400
rect 6890 21330 6910 21400
rect 6980 21330 7000 21400
rect 7070 21330 7090 21400
rect 7160 21330 7180 21400
rect 7250 21330 7290 21400
rect -5020 8690 7290 21330
rect 7610 21580 19920 21640
rect 7610 21510 7650 21580
rect 7720 21510 7740 21580
rect 7810 21510 7830 21580
rect 7900 21510 7920 21580
rect 7990 21510 8010 21580
rect 8080 21510 8100 21580
rect 8170 21510 8190 21580
rect 8260 21510 8280 21580
rect 8350 21510 8370 21580
rect 8440 21510 8460 21580
rect 8530 21510 8550 21580
rect 8620 21510 8640 21580
rect 8710 21510 8730 21580
rect 8800 21510 8820 21580
rect 8890 21510 8910 21580
rect 8980 21510 9000 21580
rect 9070 21510 9090 21580
rect 9160 21510 9180 21580
rect 9250 21510 9270 21580
rect 9340 21510 9360 21580
rect 9430 21510 9450 21580
rect 9520 21510 9540 21580
rect 9610 21510 9630 21580
rect 9700 21510 9720 21580
rect 9790 21510 9810 21580
rect 9880 21510 9900 21580
rect 9970 21510 9990 21580
rect 10060 21510 10080 21580
rect 10150 21510 10170 21580
rect 10240 21510 10260 21580
rect 10330 21510 10350 21580
rect 10420 21510 10440 21580
rect 10510 21510 10530 21580
rect 10600 21510 10660 21580
rect 10730 21510 10750 21580
rect 10820 21510 10840 21580
rect 10910 21510 10930 21580
rect 11000 21510 11020 21580
rect 11090 21510 11110 21580
rect 11180 21510 11200 21580
rect 11270 21510 11290 21580
rect 11360 21510 11380 21580
rect 11450 21510 11470 21580
rect 11540 21510 11560 21580
rect 11630 21510 11650 21580
rect 11720 21510 11740 21580
rect 11810 21510 11830 21580
rect 11900 21510 11920 21580
rect 11990 21510 12010 21580
rect 12080 21510 12100 21580
rect 12170 21510 12190 21580
rect 12260 21510 12280 21580
rect 12350 21510 12370 21580
rect 12440 21510 12460 21580
rect 12530 21510 12550 21580
rect 12620 21510 12640 21580
rect 12710 21510 12730 21580
rect 12800 21510 12820 21580
rect 12890 21510 12910 21580
rect 12980 21510 13000 21580
rect 13070 21510 13090 21580
rect 13160 21510 13180 21580
rect 13250 21510 13270 21580
rect 13340 21510 13360 21580
rect 13430 21510 13450 21580
rect 13520 21510 13540 21580
rect 13610 21510 13670 21580
rect 13740 21510 13760 21580
rect 13830 21510 13850 21580
rect 13920 21510 13940 21580
rect 14010 21510 14030 21580
rect 14100 21510 14120 21580
rect 14190 21510 14210 21580
rect 14280 21510 14300 21580
rect 14370 21510 14390 21580
rect 14460 21510 14480 21580
rect 14550 21510 14570 21580
rect 14640 21510 14660 21580
rect 14730 21510 14750 21580
rect 14820 21510 14840 21580
rect 14910 21510 14930 21580
rect 15000 21510 15020 21580
rect 15090 21510 15110 21580
rect 15180 21510 15200 21580
rect 15270 21510 15290 21580
rect 15360 21510 15380 21580
rect 15450 21510 15470 21580
rect 15540 21510 15560 21580
rect 15630 21510 15650 21580
rect 15720 21510 15740 21580
rect 15810 21510 15830 21580
rect 15900 21510 15920 21580
rect 15990 21510 16010 21580
rect 16080 21510 16100 21580
rect 16170 21510 16190 21580
rect 16260 21510 16280 21580
rect 16350 21510 16370 21580
rect 16440 21510 16460 21580
rect 16530 21510 16550 21580
rect 16620 21510 16680 21580
rect 16750 21510 16770 21580
rect 16840 21510 16860 21580
rect 16930 21510 16950 21580
rect 17020 21510 17040 21580
rect 17110 21510 17130 21580
rect 17200 21510 17220 21580
rect 17290 21510 17310 21580
rect 17380 21510 17400 21580
rect 17470 21510 17490 21580
rect 17560 21510 17580 21580
rect 17650 21510 17670 21580
rect 17740 21510 17760 21580
rect 17830 21510 17850 21580
rect 17920 21510 17940 21580
rect 18010 21510 18030 21580
rect 18100 21510 18120 21580
rect 18190 21510 18210 21580
rect 18280 21510 18300 21580
rect 18370 21510 18390 21580
rect 18460 21510 18480 21580
rect 18550 21510 18570 21580
rect 18640 21510 18660 21580
rect 18730 21510 18750 21580
rect 18820 21510 18840 21580
rect 18910 21510 18930 21580
rect 19000 21510 19020 21580
rect 19090 21510 19110 21580
rect 19180 21510 19200 21580
rect 19270 21510 19290 21580
rect 19360 21510 19380 21580
rect 19450 21510 19470 21580
rect 19540 21510 19560 21580
rect 19630 21510 19920 21580
rect 7610 21490 19920 21510
rect 7610 21420 7650 21490
rect 7720 21420 7740 21490
rect 7810 21420 7830 21490
rect 7900 21420 7920 21490
rect 7990 21420 8010 21490
rect 8080 21420 8100 21490
rect 8170 21420 8190 21490
rect 8260 21420 8280 21490
rect 8350 21420 8370 21490
rect 8440 21420 8460 21490
rect 8530 21420 8550 21490
rect 8620 21420 8640 21490
rect 8710 21420 8730 21490
rect 8800 21420 8820 21490
rect 8890 21420 8910 21490
rect 8980 21420 9000 21490
rect 9070 21420 9090 21490
rect 9160 21420 9180 21490
rect 9250 21420 9270 21490
rect 9340 21420 9360 21490
rect 9430 21420 9450 21490
rect 9520 21420 9540 21490
rect 9610 21420 9630 21490
rect 9700 21420 9720 21490
rect 9790 21420 9810 21490
rect 9880 21420 9900 21490
rect 9970 21420 9990 21490
rect 10060 21420 10080 21490
rect 10150 21420 10170 21490
rect 10240 21420 10260 21490
rect 10330 21420 10350 21490
rect 10420 21420 10440 21490
rect 10510 21420 10530 21490
rect 10600 21420 10660 21490
rect 10730 21420 10750 21490
rect 10820 21420 10840 21490
rect 10910 21420 10930 21490
rect 11000 21420 11020 21490
rect 11090 21420 11110 21490
rect 11180 21420 11200 21490
rect 11270 21420 11290 21490
rect 11360 21420 11380 21490
rect 11450 21420 11470 21490
rect 11540 21420 11560 21490
rect 11630 21420 11650 21490
rect 11720 21420 11740 21490
rect 11810 21420 11830 21490
rect 11900 21420 11920 21490
rect 11990 21420 12010 21490
rect 12080 21420 12100 21490
rect 12170 21420 12190 21490
rect 12260 21420 12280 21490
rect 12350 21420 12370 21490
rect 12440 21420 12460 21490
rect 12530 21420 12550 21490
rect 12620 21420 12640 21490
rect 12710 21420 12730 21490
rect 12800 21420 12820 21490
rect 12890 21420 12910 21490
rect 12980 21420 13000 21490
rect 13070 21420 13090 21490
rect 13160 21420 13180 21490
rect 13250 21420 13270 21490
rect 13340 21420 13360 21490
rect 13430 21420 13450 21490
rect 13520 21420 13540 21490
rect 13610 21420 13670 21490
rect 13740 21420 13760 21490
rect 13830 21420 13850 21490
rect 13920 21420 13940 21490
rect 14010 21420 14030 21490
rect 14100 21420 14120 21490
rect 14190 21420 14210 21490
rect 14280 21420 14300 21490
rect 14370 21420 14390 21490
rect 14460 21420 14480 21490
rect 14550 21420 14570 21490
rect 14640 21420 14660 21490
rect 14730 21420 14750 21490
rect 14820 21420 14840 21490
rect 14910 21420 14930 21490
rect 15000 21420 15020 21490
rect 15090 21420 15110 21490
rect 15180 21420 15200 21490
rect 15270 21420 15290 21490
rect 15360 21420 15380 21490
rect 15450 21420 15470 21490
rect 15540 21420 15560 21490
rect 15630 21420 15650 21490
rect 15720 21420 15740 21490
rect 15810 21420 15830 21490
rect 15900 21420 15920 21490
rect 15990 21420 16010 21490
rect 16080 21420 16100 21490
rect 16170 21420 16190 21490
rect 16260 21420 16280 21490
rect 16350 21420 16370 21490
rect 16440 21420 16460 21490
rect 16530 21420 16550 21490
rect 16620 21420 16680 21490
rect 16750 21420 16770 21490
rect 16840 21420 16860 21490
rect 16930 21420 16950 21490
rect 17020 21420 17040 21490
rect 17110 21420 17130 21490
rect 17200 21420 17220 21490
rect 17290 21420 17310 21490
rect 17380 21420 17400 21490
rect 17470 21420 17490 21490
rect 17560 21420 17580 21490
rect 17650 21420 17670 21490
rect 17740 21420 17760 21490
rect 17830 21420 17850 21490
rect 17920 21420 17940 21490
rect 18010 21420 18030 21490
rect 18100 21420 18120 21490
rect 18190 21420 18210 21490
rect 18280 21420 18300 21490
rect 18370 21420 18390 21490
rect 18460 21420 18480 21490
rect 18550 21420 18570 21490
rect 18640 21420 18660 21490
rect 18730 21420 18750 21490
rect 18820 21420 18840 21490
rect 18910 21420 18930 21490
rect 19000 21420 19020 21490
rect 19090 21420 19110 21490
rect 19180 21420 19200 21490
rect 19270 21420 19290 21490
rect 19360 21420 19380 21490
rect 19450 21420 19470 21490
rect 19540 21420 19560 21490
rect 19630 21420 19920 21490
rect 7610 21400 19920 21420
rect 7610 21330 7650 21400
rect 7720 21330 7740 21400
rect 7810 21330 7830 21400
rect 7900 21330 7920 21400
rect 7990 21330 8010 21400
rect 8080 21330 8100 21400
rect 8170 21330 8190 21400
rect 8260 21330 8280 21400
rect 8350 21330 8370 21400
rect 8440 21330 8460 21400
rect 8530 21330 8550 21400
rect 8620 21330 8640 21400
rect 8710 21330 8730 21400
rect 8800 21330 8820 21400
rect 8890 21330 8910 21400
rect 8980 21330 9000 21400
rect 9070 21330 9090 21400
rect 9160 21330 9180 21400
rect 9250 21330 9270 21400
rect 9340 21330 9360 21400
rect 9430 21330 9450 21400
rect 9520 21330 9540 21400
rect 9610 21330 9630 21400
rect 9700 21330 9720 21400
rect 9790 21330 9810 21400
rect 9880 21330 9900 21400
rect 9970 21330 9990 21400
rect 10060 21330 10080 21400
rect 10150 21330 10170 21400
rect 10240 21330 10260 21400
rect 10330 21330 10350 21400
rect 10420 21330 10440 21400
rect 10510 21330 10530 21400
rect 10600 21330 10660 21400
rect 10730 21330 10750 21400
rect 10820 21330 10840 21400
rect 10910 21330 10930 21400
rect 11000 21330 11020 21400
rect 11090 21330 11110 21400
rect 11180 21330 11200 21400
rect 11270 21330 11290 21400
rect 11360 21330 11380 21400
rect 11450 21330 11470 21400
rect 11540 21330 11560 21400
rect 11630 21330 11650 21400
rect 11720 21330 11740 21400
rect 11810 21330 11830 21400
rect 11900 21330 11920 21400
rect 11990 21330 12010 21400
rect 12080 21330 12100 21400
rect 12170 21330 12190 21400
rect 12260 21330 12280 21400
rect 12350 21330 12370 21400
rect 12440 21330 12460 21400
rect 12530 21330 12550 21400
rect 12620 21330 12640 21400
rect 12710 21330 12730 21400
rect 12800 21330 12820 21400
rect 12890 21330 12910 21400
rect 12980 21330 13000 21400
rect 13070 21330 13090 21400
rect 13160 21330 13180 21400
rect 13250 21330 13270 21400
rect 13340 21330 13360 21400
rect 13430 21330 13450 21400
rect 13520 21330 13540 21400
rect 13610 21330 13670 21400
rect 13740 21330 13760 21400
rect 13830 21330 13850 21400
rect 13920 21330 13940 21400
rect 14010 21330 14030 21400
rect 14100 21330 14120 21400
rect 14190 21330 14210 21400
rect 14280 21330 14300 21400
rect 14370 21330 14390 21400
rect 14460 21330 14480 21400
rect 14550 21330 14570 21400
rect 14640 21330 14660 21400
rect 14730 21330 14750 21400
rect 14820 21330 14840 21400
rect 14910 21330 14930 21400
rect 15000 21330 15020 21400
rect 15090 21330 15110 21400
rect 15180 21330 15200 21400
rect 15270 21330 15290 21400
rect 15360 21330 15380 21400
rect 15450 21330 15470 21400
rect 15540 21330 15560 21400
rect 15630 21330 15650 21400
rect 15720 21330 15740 21400
rect 15810 21330 15830 21400
rect 15900 21330 15920 21400
rect 15990 21330 16010 21400
rect 16080 21330 16100 21400
rect 16170 21330 16190 21400
rect 16260 21330 16280 21400
rect 16350 21330 16370 21400
rect 16440 21330 16460 21400
rect 16530 21330 16550 21400
rect 16620 21330 16680 21400
rect 16750 21330 16770 21400
rect 16840 21330 16860 21400
rect 16930 21330 16950 21400
rect 17020 21330 17040 21400
rect 17110 21330 17130 21400
rect 17200 21330 17220 21400
rect 17290 21330 17310 21400
rect 17380 21330 17400 21400
rect 17470 21330 17490 21400
rect 17560 21330 17580 21400
rect 17650 21330 17670 21400
rect 17740 21330 17760 21400
rect 17830 21330 17850 21400
rect 17920 21330 17940 21400
rect 18010 21330 18030 21400
rect 18100 21330 18120 21400
rect 18190 21330 18210 21400
rect 18280 21330 18300 21400
rect 18370 21330 18390 21400
rect 18460 21330 18480 21400
rect 18550 21330 18570 21400
rect 18640 21330 18660 21400
rect 18730 21330 18750 21400
rect 18820 21330 18840 21400
rect 18910 21330 18930 21400
rect 19000 21330 19020 21400
rect 19090 21330 19110 21400
rect 19180 21330 19200 21400
rect 19270 21330 19290 21400
rect 19360 21330 19380 21400
rect 19450 21330 19470 21400
rect 19540 21330 19560 21400
rect 19630 21330 19920 21400
rect 7610 8690 19920 21330
rect 7020 8410 7340 8430
rect 7020 8340 7040 8410
rect 7140 8340 7170 8410
rect 7270 8340 7340 8410
rect 7020 8320 7340 8340
rect 7020 8250 7040 8320
rect 7140 8250 7170 8320
rect 7270 8250 7340 8320
rect 1540 6850 3140 6900
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1750 6780 1790 6850
rect 1860 6780 1900 6850
rect 1970 6780 2010 6850
rect 2080 6780 2120 6850
rect 2190 6780 2230 6850
rect 2300 6780 2340 6850
rect 2410 6780 2450 6850
rect 2520 6780 2560 6850
rect 2630 6780 2670 6850
rect 2740 6780 2780 6850
rect 2850 6780 2890 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1750 6670 1790 6740
rect 1860 6670 1900 6740
rect 1970 6670 2010 6740
rect 2080 6670 2120 6740
rect 2190 6670 2230 6740
rect 2300 6670 2340 6740
rect 2410 6670 2450 6740
rect 2520 6670 2560 6740
rect 2630 6670 2670 6740
rect 2740 6670 2780 6740
rect 2850 6670 2890 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 1540 6640 3140 6670
rect 7020 4610 7340 8250
rect 7560 8410 7880 8430
rect 7560 8340 7630 8410
rect 7730 8340 7760 8410
rect 7860 8340 7880 8410
rect 7560 8320 7880 8340
rect 7560 8250 7630 8320
rect 7730 8250 7760 8320
rect 7860 8250 7880 8320
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5210 7490 5280
rect 7400 5170 7490 5210
rect 7400 5100 7410 5170
rect 7480 5100 7490 5170
rect 7400 5060 7490 5100
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 7560 4760 7880 8250
rect 31100 7820 38500 7910
rect 31100 7750 38190 7820
rect 38260 7750 38280 7820
rect 38350 7750 38370 7820
rect 38440 7750 38500 7820
rect 31100 7730 38500 7750
rect 31100 7660 38190 7730
rect 38260 7660 38280 7730
rect 38350 7660 38370 7730
rect 38440 7660 38500 7730
rect 31100 7640 38500 7660
rect 31100 7570 38190 7640
rect 38260 7570 38280 7640
rect 38350 7570 38370 7640
rect 38440 7570 38500 7640
rect 31100 7550 38500 7570
rect 31100 7480 38190 7550
rect 38260 7480 38280 7550
rect 38350 7480 38370 7550
rect 38440 7480 38500 7550
rect 31100 7460 38500 7480
rect 31100 7390 38190 7460
rect 38260 7390 38280 7460
rect 38350 7390 38370 7460
rect 38440 7390 38500 7460
rect 31100 7370 38500 7390
rect 31100 7300 38190 7370
rect 38260 7300 38280 7370
rect 38350 7300 38370 7370
rect 38440 7300 38500 7370
rect 31100 7280 38500 7300
rect 23460 7210 23940 7260
rect 23460 7140 23490 7210
rect 23560 7140 23600 7210
rect 23670 7140 23710 7210
rect 23780 7140 23820 7210
rect 23890 7140 23940 7210
rect 23460 7100 23940 7140
rect 23460 7030 23490 7100
rect 23560 7030 23600 7100
rect 23670 7030 23710 7100
rect 23780 7030 23820 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 25860 7210 26340 7260
rect 25860 7140 25890 7210
rect 25960 7140 26000 7210
rect 26070 7140 26110 7210
rect 26180 7140 26220 7210
rect 26290 7140 26340 7210
rect 25860 7100 26340 7140
rect 25860 7030 25890 7100
rect 25960 7030 26000 7100
rect 26070 7030 26110 7100
rect 26180 7030 26220 7100
rect 26290 7030 26340 7100
rect 25860 7000 26340 7030
rect 31100 7210 38190 7280
rect 38260 7210 38280 7280
rect 38350 7210 38370 7280
rect 38440 7210 38500 7280
rect 31100 7150 38500 7210
rect 31100 7080 38190 7150
rect 38260 7080 38280 7150
rect 38350 7080 38370 7150
rect 38440 7080 38500 7150
rect 31100 7060 38500 7080
rect 31100 6990 38190 7060
rect 38260 6990 38280 7060
rect 38350 6990 38370 7060
rect 38440 6990 38500 7060
rect 31100 6970 38500 6990
rect 11760 6880 13360 6930
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 11970 6810 12010 6880
rect 12080 6810 12120 6880
rect 12190 6810 12230 6880
rect 12300 6810 12340 6880
rect 12410 6810 12450 6880
rect 12520 6810 12560 6880
rect 12630 6810 12670 6880
rect 12740 6810 12780 6880
rect 12850 6810 12890 6880
rect 12960 6810 13000 6880
rect 13070 6810 13110 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 11970 6700 12010 6770
rect 12080 6700 12120 6770
rect 12190 6700 12230 6770
rect 12300 6700 12340 6770
rect 12410 6700 12450 6770
rect 12520 6700 12560 6770
rect 12630 6700 12670 6770
rect 12740 6700 12780 6770
rect 12850 6700 12890 6770
rect 12960 6700 13000 6770
rect 13070 6700 13110 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 31100 6900 38190 6970
rect 38260 6900 38280 6970
rect 38350 6900 38370 6970
rect 38440 6900 38500 6970
rect 31100 6880 38500 6900
rect 31100 6810 38190 6880
rect 38260 6810 38280 6880
rect 38350 6810 38370 6880
rect 38440 6810 38500 6880
rect 31100 6790 38500 6810
rect 31100 6720 38190 6790
rect 38260 6720 38280 6790
rect 38350 6720 38370 6790
rect 38440 6720 38500 6790
rect 31100 6700 38500 6720
rect 31100 6630 38190 6700
rect 38260 6630 38280 6700
rect 38350 6630 38370 6700
rect 38440 6630 38500 6700
rect 31100 6610 38500 6630
rect 31100 6540 38190 6610
rect 38260 6540 38280 6610
rect 38350 6540 38370 6610
rect 38440 6540 38500 6610
rect 31100 6520 38500 6540
rect 31100 6450 38190 6520
rect 38260 6450 38280 6520
rect 38350 6450 38370 6520
rect 38440 6450 38500 6520
rect 31100 6430 38500 6450
rect 31100 6360 38190 6430
rect 38260 6360 38280 6430
rect 38350 6360 38370 6430
rect 38440 6360 38500 6430
rect 31100 6340 38500 6360
rect 30720 6300 30940 6320
rect 30720 6230 30740 6300
rect 30810 6230 30850 6300
rect 30920 6230 30940 6300
rect 30720 6170 30940 6230
rect 30720 6100 30740 6170
rect 30810 6100 30850 6170
rect 30920 6100 30940 6170
rect 30720 6040 30940 6100
rect 30720 5970 30740 6040
rect 30810 5970 30850 6040
rect 30920 5970 30940 6040
rect 30720 5950 30940 5970
rect 31100 6270 38190 6340
rect 38260 6270 38280 6340
rect 38350 6270 38370 6340
rect 38440 6270 38500 6340
rect 31100 6250 38500 6270
rect 31100 6180 38190 6250
rect 38260 6180 38280 6250
rect 38350 6180 38370 6250
rect 38440 6180 38500 6250
rect 31100 6160 38500 6180
rect 31100 6090 38190 6160
rect 38260 6090 38280 6160
rect 38350 6090 38370 6160
rect 38440 6090 38500 6160
rect 31100 6070 38500 6090
rect 31100 6000 38190 6070
rect 38260 6000 38280 6070
rect 38350 6000 38370 6070
rect 38440 6000 38500 6070
rect 31100 5980 38500 6000
rect 31100 5910 38190 5980
rect 38260 5910 38280 5980
rect 38350 5910 38370 5980
rect 38440 5910 38500 5980
rect 31100 5890 38500 5910
rect 31100 5820 38190 5890
rect 38260 5820 38280 5890
rect 38350 5820 38370 5890
rect 38440 5820 38500 5890
rect 31100 5800 38500 5820
rect 31100 5730 38190 5800
rect 38260 5730 38280 5800
rect 38350 5730 38370 5800
rect 38440 5730 38500 5800
rect 31100 5710 38500 5730
rect 7560 4700 7590 4760
rect 7650 4700 7690 4760
rect 7750 4700 7790 4760
rect 7850 4700 7880 4760
rect 7560 4670 7880 4700
rect 21800 5670 22020 5690
rect 21800 5600 21820 5670
rect 21890 5600 21930 5670
rect 22000 5600 22020 5670
rect 21800 5560 22020 5600
rect 21800 5490 21820 5560
rect 21890 5490 21930 5560
rect 22000 5490 22020 5560
rect 21800 5450 22020 5490
rect 21800 5380 21820 5450
rect 21890 5380 21930 5450
rect 22000 5380 22020 5450
rect 21800 5340 22020 5380
rect 21800 5270 21820 5340
rect 21890 5270 21930 5340
rect 22000 5270 22020 5340
rect 21800 5230 22020 5270
rect 21800 5160 21820 5230
rect 21890 5160 21930 5230
rect 22000 5160 22020 5230
rect 21800 5120 22020 5160
rect 21800 5050 21820 5120
rect 21890 5050 21930 5120
rect 22000 5050 22020 5120
rect 21800 5010 22020 5050
rect 21800 4940 21820 5010
rect 21890 4940 21930 5010
rect 22000 4940 22020 5010
rect 21800 4900 22020 4940
rect 21800 4830 21820 4900
rect 21890 4830 21930 4900
rect 22000 4830 22020 4900
rect 21800 4790 22020 4830
rect 21800 4720 21820 4790
rect 21890 4720 21930 4790
rect 22000 4720 22020 4790
rect 21800 4680 22020 4720
rect 21800 4610 21820 4680
rect 21890 4610 21930 4680
rect 22000 4610 22020 4680
rect -1740 4580 6790 4610
rect -1740 4510 -1710 4580
rect -1640 4520 6700 4580
rect 6760 4520 6790 4580
rect -1640 4510 6790 4520
rect -1740 4470 6790 4510
rect -1740 4400 -1710 4470
rect -1640 4460 6790 4470
rect -1640 4400 6700 4460
rect 6760 4400 6790 4460
rect -1740 4360 6790 4400
rect -1740 4290 -1710 4360
rect -1640 4340 6790 4360
rect -1640 4290 6700 4340
rect -1740 4280 6700 4290
rect 6760 4280 6790 4340
rect -1740 4250 6790 4280
rect -1740 4180 -1710 4250
rect -1640 4220 6790 4250
rect -1640 4180 6700 4220
rect -1740 4160 6700 4180
rect 6760 4160 6790 4220
rect -1740 4130 6790 4160
rect 7020 4580 16520 4610
rect 7020 4510 16420 4580
rect 16490 4510 16520 4580
rect 7020 4470 16520 4510
rect 21800 4570 22020 4610
rect 21800 4500 21820 4570
rect 21890 4500 21930 4570
rect 22000 4500 22020 4570
rect 21800 4480 22020 4500
rect 31100 5640 38190 5710
rect 38260 5640 38280 5710
rect 38350 5640 38370 5710
rect 38440 5640 38500 5710
rect 31100 5620 38500 5640
rect 31100 5550 38190 5620
rect 38260 5550 38280 5620
rect 38350 5550 38370 5620
rect 38440 5550 38500 5620
rect 31100 5530 38500 5550
rect 31100 5460 38190 5530
rect 38260 5460 38280 5530
rect 38350 5460 38370 5530
rect 38440 5460 38500 5530
rect 31100 5440 38500 5460
rect 31100 5370 38190 5440
rect 38260 5370 38280 5440
rect 38350 5370 38370 5440
rect 38440 5370 38500 5440
rect 31100 5350 38500 5370
rect 31100 5280 38190 5350
rect 38260 5280 38280 5350
rect 38350 5280 38370 5350
rect 38440 5280 38500 5350
rect 31100 5260 38500 5280
rect 31100 5190 38190 5260
rect 38260 5190 38280 5260
rect 38350 5190 38370 5260
rect 38440 5190 38500 5260
rect 31100 5170 38500 5190
rect 31100 5100 38190 5170
rect 38260 5100 38280 5170
rect 38350 5100 38370 5170
rect 38440 5100 38500 5170
rect 31100 5080 38500 5100
rect 31100 5010 38190 5080
rect 38260 5010 38280 5080
rect 38350 5010 38370 5080
rect 38440 5010 38500 5080
rect 31100 4990 38500 5010
rect 31100 4920 38190 4990
rect 38260 4920 38280 4990
rect 38350 4920 38370 4990
rect 38440 4920 38500 4990
rect 31100 4900 38500 4920
rect 31100 4830 38190 4900
rect 38260 4830 38280 4900
rect 38350 4830 38370 4900
rect 38440 4830 38500 4900
rect 31100 4810 38500 4830
rect 31100 4740 38190 4810
rect 38260 4740 38280 4810
rect 38350 4740 38370 4810
rect 38440 4740 38500 4810
rect 31100 4720 38500 4740
rect 31100 4650 38190 4720
rect 38260 4650 38280 4720
rect 38350 4650 38370 4720
rect 38440 4650 38500 4720
rect 31100 4630 38500 4650
rect 31100 4560 38190 4630
rect 38260 4560 38280 4630
rect 38350 4560 38370 4630
rect 38440 4560 38500 4630
rect 31100 4540 38500 4560
rect 7020 4400 16420 4470
rect 16490 4400 16520 4470
rect 7020 4360 16520 4400
rect 7020 4290 16420 4360
rect 16490 4290 16520 4360
rect 7020 4250 16520 4290
rect 7020 4180 16420 4250
rect 16490 4180 16520 4250
rect 7020 4130 16520 4180
rect 31100 4470 38190 4540
rect 38260 4470 38280 4540
rect 38350 4470 38370 4540
rect 38440 4470 38500 4540
rect 31100 4450 38500 4470
rect 31100 4380 38190 4450
rect 38260 4380 38280 4450
rect 38350 4380 38370 4450
rect 38440 4380 38500 4450
rect 31100 4360 38500 4380
rect 31100 4290 38190 4360
rect 38260 4290 38280 4360
rect 38350 4290 38370 4360
rect 38440 4290 38500 4360
rect 31100 4270 38500 4290
rect 31100 4200 38190 4270
rect 38260 4200 38280 4270
rect 38350 4200 38370 4270
rect 38440 4200 38500 4270
rect 31100 4140 38500 4200
rect 7020 3240 7340 4130
rect 31100 4070 38190 4140
rect 38260 4070 38280 4140
rect 38350 4070 38370 4140
rect 38440 4070 38500 4140
rect 31100 4050 38500 4070
rect 31100 3980 38190 4050
rect 38260 3980 38280 4050
rect 38350 3980 38370 4050
rect 38440 3980 38500 4050
rect 31100 3960 38500 3980
rect 31100 3890 38190 3960
rect 38260 3890 38280 3960
rect 38350 3890 38370 3960
rect 38440 3890 38500 3960
rect 31100 3870 38500 3890
rect 31100 3800 38190 3870
rect 38260 3800 38280 3870
rect 38350 3800 38370 3870
rect 38440 3800 38500 3870
rect 31100 3780 38500 3800
rect 31100 3710 38190 3780
rect 38260 3710 38280 3780
rect 38350 3710 38370 3780
rect 38440 3710 38500 3780
rect 31100 3690 38500 3710
rect 31100 3620 38190 3690
rect 38260 3620 38280 3690
rect 38350 3620 38370 3690
rect 38440 3620 38500 3690
rect 31100 3600 38500 3620
rect 31100 3530 38190 3600
rect 38260 3530 38280 3600
rect 38350 3530 38370 3600
rect 38440 3530 38500 3600
rect 31100 3510 38500 3530
rect 31100 3440 38190 3510
rect 38260 3440 38280 3510
rect 38350 3440 38370 3510
rect 38440 3440 38500 3510
rect 31100 3420 38500 3440
rect 7020 3180 7050 3240
rect 7110 3180 7150 3240
rect 7210 3180 7250 3240
rect 7310 3180 7340 3240
rect 7020 3140 7340 3180
rect 7020 3080 7050 3140
rect 7110 3080 7150 3140
rect 7210 3080 7250 3140
rect 7310 3080 7340 3140
rect 7020 3040 7340 3080
rect 24700 3360 25030 3380
rect 24700 3290 24720 3360
rect 24790 3290 24830 3360
rect 24900 3290 24940 3360
rect 25010 3290 25030 3360
rect 24700 3250 25030 3290
rect 24700 3180 24720 3250
rect 24790 3180 24830 3250
rect 24900 3180 24940 3250
rect 25010 3180 25030 3250
rect 24700 3140 25030 3180
rect 24700 3070 24720 3140
rect 24790 3070 24830 3140
rect 24900 3070 24940 3140
rect 25010 3070 25030 3140
rect 24700 3050 25030 3070
rect 31100 3350 38190 3420
rect 38260 3350 38280 3420
rect 38350 3350 38370 3420
rect 38440 3350 38500 3420
rect 31100 3330 38500 3350
rect 31100 3260 38190 3330
rect 38260 3260 38280 3330
rect 38350 3260 38370 3330
rect 38440 3260 38500 3330
rect 31100 3240 38500 3260
rect 31100 3170 38190 3240
rect 38260 3170 38280 3240
rect 38350 3170 38370 3240
rect 38440 3170 38500 3240
rect 31100 3150 38500 3170
rect 31100 3080 38190 3150
rect 38260 3080 38280 3150
rect 38350 3080 38370 3150
rect 38440 3080 38500 3150
rect 31100 3060 38500 3080
rect 7020 2980 7050 3040
rect 7110 2980 7150 3040
rect 7210 2980 7250 3040
rect 7310 2980 7340 3040
rect 7020 2960 7340 2980
rect 31100 2990 38190 3060
rect 38260 2990 38280 3060
rect 38350 2990 38370 3060
rect 38440 2990 38500 3060
rect 31100 2970 38500 2990
rect 4740 2890 6750 2920
rect 4740 2830 4770 2890
rect 4830 2830 4870 2890
rect 4930 2830 4970 2890
rect 5030 2830 6750 2890
rect 4740 2790 6750 2830
rect 4740 2730 4770 2790
rect 4830 2730 4870 2790
rect 4930 2730 4970 2790
rect 5030 2730 6750 2790
rect 4740 2690 6750 2730
rect 4740 2630 4770 2690
rect 4830 2630 4870 2690
rect 4930 2630 4970 2690
rect 5030 2630 6750 2690
rect 4740 2610 6750 2630
rect 6440 -100 6750 2610
rect -330 -140 6750 -100
rect -330 -210 -300 -140
rect -230 -210 -190 -140
rect -120 -210 -80 -140
rect -10 -210 30 -140
rect 100 -210 6750 -140
rect -330 -270 6750 -210
rect -330 -340 -300 -270
rect -230 -340 -190 -270
rect -120 -340 -80 -270
rect -10 -340 30 -270
rect 100 -340 6750 -270
rect -330 -380 6750 -340
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1330 -860 1370 -790
rect 1440 -860 1480 -790
rect 1550 -860 1590 -790
rect 1660 -860 1700 -790
rect 1770 -860 1810 -790
rect 1880 -860 1920 -790
rect 1990 -860 2030 -790
rect 2100 -860 2140 -790
rect 2210 -860 2250 -790
rect 2320 -860 2360 -790
rect 2430 -860 2470 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1330 -970 1370 -900
rect 1440 -970 1480 -900
rect 1550 -970 1590 -900
rect 1660 -970 1700 -900
rect 1770 -970 1810 -900
rect 1880 -970 1920 -900
rect 1990 -970 2030 -900
rect 2100 -970 2140 -900
rect 2210 -970 2250 -900
rect 2320 -970 2360 -900
rect 2430 -970 2470 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1020 2680 -970
rect 1540 -2780 3140 -2730
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1750 -2850 1790 -2780
rect 1860 -2850 1900 -2780
rect 1970 -2850 2010 -2780
rect 2080 -2850 2120 -2780
rect 2190 -2850 2230 -2780
rect 2300 -2850 2340 -2780
rect 2410 -2850 2450 -2780
rect 2520 -2850 2560 -2780
rect 2630 -2850 2670 -2780
rect 2740 -2850 2780 -2780
rect 2850 -2850 2890 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1750 -2960 1790 -2890
rect 1860 -2960 1900 -2890
rect 1970 -2960 2010 -2890
rect 2080 -2960 2120 -2890
rect 2190 -2960 2230 -2890
rect 2300 -2960 2340 -2890
rect 2410 -2960 2450 -2890
rect 2520 -2960 2560 -2890
rect 2630 -2960 2670 -2890
rect 2740 -2960 2780 -2890
rect 2850 -2960 2890 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 6440 -4270 6750 -380
rect 8180 2890 10160 2920
rect 8180 2830 9870 2890
rect 9930 2830 9970 2890
rect 10030 2830 10070 2890
rect 10130 2830 10160 2890
rect 8180 2790 10160 2830
rect 8180 2730 9870 2790
rect 9930 2730 9970 2790
rect 10030 2730 10070 2790
rect 10130 2730 10160 2790
rect 8180 2690 10160 2730
rect 8180 2630 9870 2690
rect 9930 2630 9970 2690
rect 10030 2630 10070 2690
rect 10130 2630 10160 2690
rect 31100 2900 38190 2970
rect 38260 2900 38280 2970
rect 38350 2900 38370 2970
rect 38440 2900 38500 2970
rect 31100 2880 38500 2900
rect 31100 2810 38190 2880
rect 38260 2810 38280 2880
rect 38350 2810 38370 2880
rect 38440 2810 38500 2880
rect 31100 2790 38500 2810
rect 31100 2720 38190 2790
rect 38260 2720 38280 2790
rect 38350 2720 38370 2790
rect 38440 2720 38500 2790
rect 31100 2700 38500 2720
rect 31100 2630 38190 2700
rect 38260 2630 38280 2700
rect 38350 2630 38370 2700
rect 38440 2630 38500 2700
rect 8180 2610 10160 2630
rect 8180 -100 8490 2610
rect 22420 2600 22900 2630
rect 22420 2530 22470 2600
rect 22540 2530 22580 2600
rect 22650 2530 22690 2600
rect 22760 2530 22800 2600
rect 22870 2530 22900 2600
rect 22420 2490 22900 2530
rect 22420 2420 22470 2490
rect 22540 2420 22580 2490
rect 22650 2420 22690 2490
rect 22760 2420 22800 2490
rect 22870 2420 22900 2490
rect 22420 2370 22900 2420
rect 26900 2600 27380 2630
rect 26900 2530 26950 2600
rect 27020 2530 27060 2600
rect 27130 2530 27170 2600
rect 27240 2530 27280 2600
rect 27350 2530 27380 2600
rect 26900 2490 27380 2530
rect 26900 2420 26950 2490
rect 27020 2420 27060 2490
rect 27130 2420 27170 2490
rect 27240 2420 27280 2490
rect 27350 2420 27380 2490
rect 26900 2370 27380 2420
rect 31100 2610 38500 2630
rect 31100 2540 38190 2610
rect 38260 2540 38280 2610
rect 38350 2540 38370 2610
rect 38440 2540 38500 2610
rect 31100 2520 38500 2540
rect 31100 2450 38190 2520
rect 38260 2450 38280 2520
rect 38350 2450 38370 2520
rect 38440 2450 38500 2520
rect 31100 2430 38500 2450
rect 31100 2360 38190 2430
rect 38260 2360 38280 2430
rect 38350 2360 38370 2430
rect 38440 2360 38500 2430
rect 31100 2340 38500 2360
rect 31100 2270 38190 2340
rect 38260 2270 38280 2340
rect 38350 2270 38370 2340
rect 38440 2270 38500 2340
rect 31100 2250 38500 2270
rect 31100 2180 38190 2250
rect 38260 2180 38280 2250
rect 38350 2180 38370 2250
rect 38440 2180 38500 2250
rect 31100 2160 38500 2180
rect 31100 2090 38190 2160
rect 38260 2090 38280 2160
rect 38350 2090 38370 2160
rect 38440 2090 38500 2160
rect 31100 2070 38500 2090
rect 31100 2000 38190 2070
rect 38260 2000 38280 2070
rect 38350 2000 38370 2070
rect 38440 2000 38500 2070
rect 31100 1980 38500 2000
rect 31100 1910 38190 1980
rect 38260 1910 38280 1980
rect 38350 1910 38370 1980
rect 38440 1910 38500 1980
rect 31100 1890 38500 1910
rect 31100 1820 38190 1890
rect 38260 1820 38280 1890
rect 38350 1820 38370 1890
rect 38440 1820 38500 1890
rect 31100 1800 38500 1820
rect 31100 1730 38190 1800
rect 38260 1730 38280 1800
rect 38350 1730 38370 1800
rect 38440 1730 38500 1800
rect 31100 1710 38500 1730
rect 31100 1640 38190 1710
rect 38260 1640 38280 1710
rect 38350 1640 38370 1710
rect 38440 1640 38500 1710
rect 31100 1620 38500 1640
rect 31100 1550 38190 1620
rect 38260 1550 38280 1620
rect 38350 1550 38370 1620
rect 38440 1550 38500 1620
rect 31100 1530 38500 1550
rect 31100 1460 38190 1530
rect 38260 1460 38280 1530
rect 38350 1460 38370 1530
rect 38440 1460 38500 1530
rect 31100 1440 38500 1460
rect 31100 1370 38190 1440
rect 38260 1370 38280 1440
rect 38350 1370 38370 1440
rect 38440 1370 38500 1440
rect 31100 1350 38500 1370
rect 31100 1280 38190 1350
rect 38260 1280 38280 1350
rect 38350 1280 38370 1350
rect 38440 1280 38500 1350
rect 31100 1260 38500 1280
rect 31100 1190 38190 1260
rect 38260 1190 38280 1260
rect 38350 1190 38370 1260
rect 38440 1190 38500 1260
rect 14590 1160 17580 1180
rect 14590 1090 14600 1160
rect 14670 1090 14700 1160
rect 14770 1090 14810 1160
rect 14880 1090 17480 1160
rect 17550 1090 17580 1160
rect 31100 1150 38500 1190
rect 14590 1050 17580 1090
rect 14590 980 14600 1050
rect 14670 980 14700 1050
rect 14770 980 14810 1050
rect 14880 980 17480 1050
rect 17550 980 17580 1050
rect 14590 940 17580 980
rect 14590 870 14600 940
rect 14670 870 14700 940
rect 14770 870 14810 940
rect 14880 870 17480 940
rect 17550 870 17580 940
rect 14590 850 17580 870
rect 23460 920 23940 970
rect 23460 850 23490 920
rect 23560 850 23600 920
rect 23670 850 23710 920
rect 23780 850 23820 920
rect 23890 850 23940 920
rect 23460 810 23940 850
rect 23460 740 23490 810
rect 23560 740 23600 810
rect 23670 740 23710 810
rect 23780 740 23820 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 25860 920 26340 970
rect 25860 850 25890 920
rect 25960 850 26000 920
rect 26070 850 26110 920
rect 26180 850 26220 920
rect 26290 850 26340 920
rect 25860 810 26340 850
rect 25860 740 25890 810
rect 25960 740 26000 810
rect 26070 740 26110 810
rect 26180 740 26220 810
rect 26290 740 26340 810
rect 25860 710 26340 740
rect 31100 220 38500 310
rect 31100 150 38190 220
rect 38260 150 38280 220
rect 38350 150 38370 220
rect 38440 150 38500 220
rect 31100 130 38500 150
rect 31100 60 38190 130
rect 38260 60 38280 130
rect 38350 60 38370 130
rect 38440 60 38500 130
rect 31100 40 38500 60
rect 30720 0 30940 20
rect 30720 -70 30740 0
rect 30810 -70 30850 0
rect 30920 -70 30940 0
rect 8180 -140 15110 -100
rect 8180 -210 14660 -140
rect 14730 -210 14770 -140
rect 14840 -210 14880 -140
rect 14950 -210 14990 -140
rect 15060 -210 15110 -140
rect 8180 -270 15110 -210
rect 8180 -340 14660 -270
rect 14730 -340 14770 -270
rect 14840 -340 14880 -270
rect 14950 -340 14990 -270
rect 15060 -340 15110 -270
rect 8180 -380 15110 -340
rect 30720 -130 30940 -70
rect 30720 -200 30740 -130
rect 30810 -200 30850 -130
rect 30920 -200 30940 -130
rect 30720 -260 30940 -200
rect 30720 -330 30740 -260
rect 30810 -330 30850 -260
rect 30920 -330 30940 -260
rect 30720 -350 30940 -330
rect 31100 -30 38190 40
rect 38260 -30 38280 40
rect 38350 -30 38370 40
rect 38440 -30 38500 40
rect 31100 -50 38500 -30
rect 31100 -120 38190 -50
rect 38260 -120 38280 -50
rect 38350 -120 38370 -50
rect 38440 -120 38500 -50
rect 31100 -140 38500 -120
rect 31100 -210 38190 -140
rect 38260 -210 38280 -140
rect 38350 -210 38370 -140
rect 38440 -210 38500 -140
rect 31100 -230 38500 -210
rect 31100 -300 38190 -230
rect 38260 -300 38280 -230
rect 38350 -300 38370 -230
rect 38440 -300 38500 -230
rect 31100 -320 38500 -300
rect 7290 -3880 7620 -3860
rect 7290 -3950 7310 -3880
rect 7380 -3950 7420 -3880
rect 7490 -3950 7530 -3880
rect 7600 -3950 7620 -3880
rect 7290 -3990 7620 -3950
rect 7290 -4060 7310 -3990
rect 7380 -4060 7420 -3990
rect 7490 -4060 7530 -3990
rect 7600 -4060 7620 -3990
rect 7290 -4100 7620 -4060
rect 7290 -4170 7310 -4100
rect 7380 -4170 7420 -4100
rect 7490 -4170 7530 -4100
rect 7600 -4170 7620 -4100
rect 7290 -4190 7620 -4170
rect -590 -4290 6750 -4270
rect -1350 -4350 -910 -4330
rect -1350 -4420 -1330 -4350
rect -1260 -4420 -1220 -4350
rect -1150 -4420 -1110 -4350
rect -1040 -4420 -1000 -4350
rect -930 -4420 -910 -4350
rect -1350 -4460 -910 -4420
rect -1350 -4530 -1330 -4460
rect -1260 -4530 -1220 -4460
rect -1150 -4530 -1110 -4460
rect -1040 -4530 -1000 -4460
rect -930 -4530 -910 -4460
rect -1350 -4550 -910 -4530
rect -590 -4360 -560 -4290
rect -490 -4360 -450 -4290
rect -380 -4360 -340 -4290
rect -270 -4360 -230 -4290
rect -160 -4360 6750 -4290
rect -590 -4400 6750 -4360
rect -590 -4470 -560 -4400
rect -490 -4470 -450 -4400
rect -380 -4470 -340 -4400
rect -270 -4470 -230 -4400
rect -160 -4470 6750 -4400
rect -590 -4550 6750 -4470
rect -1350 -6330 260 -4630
rect -1350 -6400 -1160 -6330
rect -1090 -6400 -1070 -6330
rect -1000 -6400 -980 -6330
rect -910 -6400 -890 -6330
rect -820 -6400 -800 -6330
rect -730 -6400 -710 -6330
rect -640 -6400 -620 -6330
rect -550 -6400 -530 -6330
rect -460 -6400 -440 -6330
rect -370 -6400 -350 -6330
rect -280 -6400 -260 -6330
rect -190 -6400 -170 -6330
rect -100 -6400 -80 -6330
rect -10 -6400 10 -6330
rect 80 -6400 260 -6330
rect -1350 -6420 260 -6400
rect -1740 -6520 -1600 -6470
rect -1740 -6590 -1710 -6520
rect -1640 -6590 -1600 -6520
rect -1740 -6630 -1600 -6590
rect -1740 -6700 -1710 -6630
rect -1640 -6640 -1600 -6630
rect -1350 -6490 -1160 -6420
rect -1090 -6490 -1070 -6420
rect -1000 -6490 -980 -6420
rect -910 -6490 -890 -6420
rect -820 -6490 -800 -6420
rect -730 -6490 -710 -6420
rect -640 -6490 -620 -6420
rect -550 -6490 -530 -6420
rect -460 -6490 -440 -6420
rect -370 -6490 -350 -6420
rect -280 -6490 -260 -6420
rect -190 -6490 -170 -6420
rect -100 -6490 -80 -6420
rect -10 -6490 10 -6420
rect 80 -6490 260 -6420
rect -1350 -6510 260 -6490
rect -1350 -6580 -1160 -6510
rect -1090 -6580 -1070 -6510
rect -1000 -6580 -980 -6510
rect -910 -6580 -890 -6510
rect -820 -6580 -800 -6510
rect -730 -6580 -710 -6510
rect -640 -6580 -620 -6510
rect -550 -6580 -530 -6510
rect -460 -6580 -440 -6510
rect -370 -6580 -350 -6510
rect -280 -6580 -260 -6510
rect -190 -6580 -170 -6510
rect -100 -6580 -80 -6510
rect -10 -6580 10 -6510
rect 80 -6580 260 -6510
rect -1350 -6640 260 -6580
rect 6440 -6420 6750 -4550
rect 8180 -4270 8490 -380
rect 31100 -390 38190 -320
rect 38260 -390 38280 -320
rect 38350 -390 38370 -320
rect 38440 -390 38500 -320
rect 31100 -450 38500 -390
rect 31100 -520 38190 -450
rect 38260 -520 38280 -450
rect 38350 -520 38370 -450
rect 38440 -520 38500 -450
rect 31100 -540 38500 -520
rect 31100 -610 38190 -540
rect 38260 -610 38280 -540
rect 38350 -610 38370 -540
rect 38440 -610 38500 -540
rect 31100 -630 38500 -610
rect 31100 -700 38190 -630
rect 38260 -700 38280 -630
rect 38350 -700 38370 -630
rect 38440 -700 38500 -630
rect 31100 -720 38500 -700
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12430 -860 12470 -790
rect 12540 -860 12580 -790
rect 12650 -860 12690 -790
rect 12760 -860 12800 -790
rect 12870 -860 12910 -790
rect 12980 -860 13020 -790
rect 13090 -860 13130 -790
rect 13200 -860 13240 -790
rect 13310 -860 13350 -790
rect 13420 -860 13460 -790
rect 13530 -860 13570 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 31100 -790 38190 -720
rect 38260 -790 38280 -720
rect 38350 -790 38370 -720
rect 38440 -790 38500 -720
rect 31100 -810 38500 -790
rect 12220 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12430 -970 12470 -900
rect 12540 -970 12580 -900
rect 12650 -970 12690 -900
rect 12760 -970 12800 -900
rect 12870 -970 12910 -900
rect 12980 -970 13020 -900
rect 13090 -970 13130 -900
rect 13200 -970 13240 -900
rect 13310 -970 13350 -900
rect 13420 -970 13460 -900
rect 13530 -970 13570 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1020 13820 -970
rect 21800 -850 22020 -830
rect 21800 -920 21820 -850
rect 21890 -920 21930 -850
rect 22000 -920 22020 -850
rect 21800 -960 22020 -920
rect 21800 -1030 21820 -960
rect 21890 -1030 21930 -960
rect 22000 -1030 22020 -960
rect 21800 -1070 22020 -1030
rect 21800 -1140 21820 -1070
rect 21890 -1140 21930 -1070
rect 22000 -1140 22020 -1070
rect 21800 -1180 22020 -1140
rect 21800 -1250 21820 -1180
rect 21890 -1250 21930 -1180
rect 22000 -1250 22020 -1180
rect 21800 -1290 22020 -1250
rect 21800 -1360 21820 -1290
rect 21890 -1360 21930 -1290
rect 22000 -1360 22020 -1290
rect 21800 -1400 22020 -1360
rect 21800 -1470 21820 -1400
rect 21890 -1470 21930 -1400
rect 22000 -1470 22020 -1400
rect 21800 -1510 22020 -1470
rect 21800 -1580 21820 -1510
rect 21890 -1580 21930 -1510
rect 22000 -1580 22020 -1510
rect 21800 -1620 22020 -1580
rect 21800 -1690 21820 -1620
rect 21890 -1690 21930 -1620
rect 22000 -1690 22020 -1620
rect 21800 -1730 22020 -1690
rect 21800 -1800 21820 -1730
rect 21890 -1800 21930 -1730
rect 22000 -1800 22020 -1730
rect 21800 -1840 22020 -1800
rect 21800 -1910 21820 -1840
rect 21890 -1910 21930 -1840
rect 22000 -1910 22020 -1840
rect 21800 -1950 22020 -1910
rect 21800 -2020 21820 -1950
rect 21890 -2020 21930 -1950
rect 22000 -2020 22020 -1950
rect 21800 -2040 22020 -2020
rect 31100 -880 38190 -810
rect 38260 -880 38280 -810
rect 38350 -880 38370 -810
rect 38440 -880 38500 -810
rect 31100 -900 38500 -880
rect 31100 -970 38190 -900
rect 38260 -970 38280 -900
rect 38350 -970 38370 -900
rect 38440 -970 38500 -900
rect 31100 -990 38500 -970
rect 31100 -1060 38190 -990
rect 38260 -1060 38280 -990
rect 38350 -1060 38370 -990
rect 38440 -1060 38500 -990
rect 31100 -1080 38500 -1060
rect 31100 -1150 38190 -1080
rect 38260 -1150 38280 -1080
rect 38350 -1150 38370 -1080
rect 38440 -1150 38500 -1080
rect 31100 -1170 38500 -1150
rect 31100 -1240 38190 -1170
rect 38260 -1240 38280 -1170
rect 38350 -1240 38370 -1170
rect 38440 -1240 38500 -1170
rect 31100 -1260 38500 -1240
rect 31100 -1330 38190 -1260
rect 38260 -1330 38280 -1260
rect 38350 -1330 38370 -1260
rect 38440 -1330 38500 -1260
rect 31100 -1350 38500 -1330
rect 31100 -1420 38190 -1350
rect 38260 -1420 38280 -1350
rect 38350 -1420 38370 -1350
rect 38440 -1420 38500 -1350
rect 31100 -1440 38500 -1420
rect 31100 -1510 38190 -1440
rect 38260 -1510 38280 -1440
rect 38350 -1510 38370 -1440
rect 38440 -1510 38500 -1440
rect 31100 -1530 38500 -1510
rect 31100 -1600 38190 -1530
rect 38260 -1600 38280 -1530
rect 38350 -1600 38370 -1530
rect 38440 -1600 38500 -1530
rect 31100 -1620 38500 -1600
rect 31100 -1690 38190 -1620
rect 38260 -1690 38280 -1620
rect 38350 -1690 38370 -1620
rect 38440 -1690 38500 -1620
rect 31100 -1710 38500 -1690
rect 31100 -1780 38190 -1710
rect 38260 -1780 38280 -1710
rect 38350 -1780 38370 -1710
rect 38440 -1780 38500 -1710
rect 31100 -1800 38500 -1780
rect 31100 -1870 38190 -1800
rect 38260 -1870 38280 -1800
rect 38350 -1870 38370 -1800
rect 38440 -1870 38500 -1800
rect 31100 -1890 38500 -1870
rect 31100 -1960 38190 -1890
rect 38260 -1960 38280 -1890
rect 38350 -1960 38370 -1890
rect 38440 -1960 38500 -1890
rect 31100 -1980 38500 -1960
rect 31100 -2050 38190 -1980
rect 38260 -2050 38280 -1980
rect 38350 -2050 38370 -1980
rect 38440 -2050 38500 -1980
rect 31100 -2070 38500 -2050
rect 31100 -2140 38190 -2070
rect 38260 -2140 38280 -2070
rect 38350 -2140 38370 -2070
rect 38440 -2140 38500 -2070
rect 31100 -2160 38500 -2140
rect 31100 -2230 38190 -2160
rect 38260 -2230 38280 -2160
rect 38350 -2230 38370 -2160
rect 38440 -2230 38500 -2160
rect 31100 -2250 38500 -2230
rect 31100 -2320 38190 -2250
rect 38260 -2320 38280 -2250
rect 38350 -2320 38370 -2250
rect 38440 -2320 38500 -2250
rect 31100 -2340 38500 -2320
rect 31100 -2410 38190 -2340
rect 38260 -2410 38280 -2340
rect 38350 -2410 38370 -2340
rect 38440 -2410 38500 -2340
rect 31100 -2430 38500 -2410
rect 31100 -2500 38190 -2430
rect 38260 -2500 38280 -2430
rect 38350 -2500 38370 -2430
rect 38440 -2500 38500 -2430
rect 31100 -2520 38500 -2500
rect 31100 -2590 38190 -2520
rect 38260 -2590 38280 -2520
rect 38350 -2590 38370 -2520
rect 38440 -2590 38500 -2520
rect 31100 -2610 38500 -2590
rect 31100 -2680 38190 -2610
rect 38260 -2680 38280 -2610
rect 38350 -2680 38370 -2610
rect 38440 -2680 38500 -2610
rect 31100 -2700 38500 -2680
rect 11760 -2780 13360 -2730
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 11970 -2850 12010 -2780
rect 12080 -2850 12120 -2780
rect 12190 -2850 12230 -2780
rect 12300 -2850 12340 -2780
rect 12410 -2850 12450 -2780
rect 12520 -2850 12560 -2780
rect 12630 -2850 12670 -2780
rect 12740 -2850 12780 -2780
rect 12850 -2850 12890 -2780
rect 12960 -2850 13000 -2780
rect 13070 -2850 13110 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 11970 -2960 12010 -2890
rect 12080 -2960 12120 -2890
rect 12190 -2960 12230 -2890
rect 12300 -2960 12340 -2890
rect 12410 -2960 12450 -2890
rect 12520 -2960 12560 -2890
rect 12630 -2960 12670 -2890
rect 12740 -2960 12780 -2890
rect 12850 -2960 12890 -2890
rect 12960 -2960 13000 -2890
rect 13070 -2960 13110 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect 31100 -2770 38190 -2700
rect 38260 -2770 38280 -2700
rect 38350 -2770 38370 -2700
rect 38440 -2770 38500 -2700
rect 31100 -2790 38500 -2770
rect 31100 -2860 38190 -2790
rect 38260 -2860 38280 -2790
rect 38350 -2860 38370 -2790
rect 38440 -2860 38500 -2790
rect 31100 -2880 38500 -2860
rect 31100 -2950 38190 -2880
rect 38260 -2950 38280 -2880
rect 38350 -2950 38370 -2880
rect 38440 -2950 38500 -2880
rect 31100 -2970 38500 -2950
rect 24720 -3050 25050 -3030
rect 24720 -3120 24740 -3050
rect 24810 -3120 24850 -3050
rect 24920 -3120 24960 -3050
rect 25030 -3120 25050 -3050
rect 24720 -3160 25050 -3120
rect 24720 -3230 24740 -3160
rect 24810 -3230 24850 -3160
rect 24920 -3230 24960 -3160
rect 25030 -3230 25050 -3160
rect 24720 -3270 25050 -3230
rect 24720 -3340 24740 -3270
rect 24810 -3340 24850 -3270
rect 24920 -3340 24960 -3270
rect 25030 -3340 25050 -3270
rect 24720 -3360 25050 -3340
rect 31100 -3040 38190 -2970
rect 38260 -3040 38280 -2970
rect 38350 -3040 38370 -2970
rect 38440 -3040 38500 -2970
rect 31100 -3060 38500 -3040
rect 31100 -3130 38190 -3060
rect 38260 -3130 38280 -3060
rect 38350 -3130 38370 -3060
rect 38440 -3130 38500 -3060
rect 31100 -3150 38500 -3130
rect 31100 -3220 38190 -3150
rect 38260 -3220 38280 -3150
rect 38350 -3220 38370 -3150
rect 38440 -3220 38500 -3150
rect 31100 -3240 38500 -3220
rect 31100 -3310 38190 -3240
rect 38260 -3310 38280 -3240
rect 38350 -3310 38370 -3240
rect 38440 -3310 38500 -3240
rect 31100 -3330 38500 -3310
rect 31100 -3400 38190 -3330
rect 38260 -3400 38280 -3330
rect 38350 -3400 38370 -3330
rect 38440 -3400 38500 -3330
rect 31100 -3460 38500 -3400
rect 31100 -3530 38190 -3460
rect 38260 -3530 38280 -3460
rect 38350 -3530 38370 -3460
rect 38440 -3530 38500 -3460
rect 31100 -3550 38500 -3530
rect 31100 -3620 38190 -3550
rect 38260 -3620 38280 -3550
rect 38350 -3620 38370 -3550
rect 38440 -3620 38500 -3550
rect 31100 -3640 38500 -3620
rect 22420 -3690 22900 -3660
rect 22420 -3760 22470 -3690
rect 22540 -3760 22580 -3690
rect 22650 -3760 22690 -3690
rect 22760 -3760 22800 -3690
rect 22870 -3760 22900 -3690
rect 22420 -3800 22900 -3760
rect 22420 -3870 22470 -3800
rect 22540 -3870 22580 -3800
rect 22650 -3870 22690 -3800
rect 22760 -3870 22800 -3800
rect 22870 -3870 22900 -3800
rect 22420 -3920 22900 -3870
rect 26900 -3690 27380 -3660
rect 26900 -3760 26950 -3690
rect 27020 -3760 27060 -3690
rect 27130 -3760 27170 -3690
rect 27240 -3760 27280 -3690
rect 27350 -3760 27380 -3690
rect 26900 -3800 27380 -3760
rect 26900 -3870 26950 -3800
rect 27020 -3870 27060 -3800
rect 27130 -3870 27170 -3800
rect 27240 -3870 27280 -3800
rect 27350 -3870 27380 -3800
rect 26900 -3920 27380 -3870
rect 31100 -3710 38190 -3640
rect 38260 -3710 38280 -3640
rect 38350 -3710 38370 -3640
rect 38440 -3710 38500 -3640
rect 31100 -3730 38500 -3710
rect 31100 -3800 38190 -3730
rect 38260 -3800 38280 -3730
rect 38350 -3800 38370 -3730
rect 38440 -3800 38500 -3730
rect 31100 -3820 38500 -3800
rect 31100 -3890 38190 -3820
rect 38260 -3890 38280 -3820
rect 38350 -3890 38370 -3820
rect 38440 -3890 38500 -3820
rect 31100 -3910 38500 -3890
rect 31100 -3980 38190 -3910
rect 38260 -3980 38280 -3910
rect 38350 -3980 38370 -3910
rect 38440 -3980 38500 -3910
rect 31100 -4000 38500 -3980
rect 31100 -4070 38190 -4000
rect 38260 -4070 38280 -4000
rect 38350 -4070 38370 -4000
rect 38440 -4070 38500 -4000
rect 31100 -4090 38500 -4070
rect 31100 -4160 38190 -4090
rect 38260 -4160 38280 -4090
rect 38350 -4160 38370 -4090
rect 38440 -4160 38500 -4090
rect 31100 -4180 38500 -4160
rect 31100 -4250 38190 -4180
rect 38260 -4250 38280 -4180
rect 38350 -4250 38370 -4180
rect 38440 -4250 38500 -4180
rect 31100 -4270 38500 -4250
rect 8180 -4290 15370 -4270
rect 8180 -4360 14940 -4290
rect 15010 -4360 15050 -4290
rect 15120 -4360 15160 -4290
rect 15230 -4360 15270 -4290
rect 15340 -4360 15370 -4290
rect 8180 -4400 15370 -4360
rect 8180 -4470 14940 -4400
rect 15010 -4470 15050 -4400
rect 15120 -4470 15160 -4400
rect 15230 -4470 15270 -4400
rect 15340 -4470 15370 -4400
rect 8180 -4550 15370 -4470
rect 15690 -4350 16130 -4330
rect 15690 -4420 15710 -4350
rect 15780 -4420 15820 -4350
rect 15890 -4420 15930 -4350
rect 16000 -4420 16040 -4350
rect 16110 -4420 16130 -4350
rect 15690 -4460 16130 -4420
rect 15690 -4530 15710 -4460
rect 15780 -4530 15820 -4460
rect 15890 -4530 15930 -4460
rect 16000 -4530 16040 -4460
rect 16110 -4530 16130 -4460
rect 15690 -4550 16130 -4530
rect 31100 -4340 38190 -4270
rect 38260 -4340 38280 -4270
rect 38350 -4340 38370 -4270
rect 38440 -4340 38500 -4270
rect 31100 -4360 38500 -4340
rect 31100 -4430 38190 -4360
rect 38260 -4430 38280 -4360
rect 38350 -4430 38370 -4360
rect 38440 -4430 38500 -4360
rect 31100 -4450 38500 -4430
rect 31100 -4520 38190 -4450
rect 38260 -4520 38280 -4450
rect 38350 -4520 38370 -4450
rect 38440 -4520 38500 -4450
rect 31100 -4540 38500 -4520
rect 8180 -6420 8490 -4550
rect 31100 -4610 38190 -4540
rect 38260 -4610 38280 -4540
rect 38350 -4610 38370 -4540
rect 38440 -4610 38500 -4540
rect 31100 -4630 38500 -4610
rect 6440 -6460 7340 -6420
rect 6440 -6520 7050 -6460
rect 7110 -6520 7150 -6460
rect 7210 -6520 7250 -6460
rect 7310 -6520 7340 -6460
rect 6440 -6560 7340 -6520
rect 6440 -6620 7050 -6560
rect 7110 -6620 7150 -6560
rect 7210 -6620 7250 -6560
rect 7310 -6620 7340 -6560
rect -1640 -6670 6190 -6640
rect -1640 -6700 4770 -6670
rect -1740 -6730 4770 -6700
rect 4830 -6730 4870 -6670
rect 4930 -6730 4970 -6670
rect 5030 -6730 6190 -6670
rect -1740 -6740 6190 -6730
rect -1740 -6810 -1710 -6740
rect -1640 -6770 6190 -6740
rect -1640 -6810 4770 -6770
rect -1740 -6830 4770 -6810
rect 4830 -6830 4870 -6770
rect 4930 -6830 4970 -6770
rect 5030 -6830 6190 -6770
rect -1740 -6850 6190 -6830
rect 6440 -6660 7340 -6620
rect 6440 -6720 7050 -6660
rect 7110 -6720 7150 -6660
rect 7210 -6720 7250 -6660
rect 7310 -6720 7340 -6660
rect 6440 -6760 7340 -6720
rect 6440 -6820 7050 -6760
rect 7110 -6820 7150 -6760
rect 7210 -6820 7250 -6760
rect 7310 -6820 7340 -6760
rect 6440 -6850 7340 -6820
rect 7560 -6460 8490 -6420
rect 7560 -6520 7590 -6460
rect 7650 -6520 7690 -6460
rect 7750 -6520 7790 -6460
rect 7850 -6520 8490 -6460
rect 7560 -6560 8490 -6520
rect 7560 -6620 7590 -6560
rect 7650 -6620 7690 -6560
rect 7750 -6620 7790 -6560
rect 7850 -6620 8490 -6560
rect 7560 -6660 8490 -6620
rect 14520 -6330 16130 -4630
rect 14520 -6400 14700 -6330
rect 14770 -6400 14790 -6330
rect 14860 -6400 14880 -6330
rect 14950 -6400 14970 -6330
rect 15040 -6400 15060 -6330
rect 15130 -6400 15150 -6330
rect 15220 -6400 15240 -6330
rect 15310 -6400 15330 -6330
rect 15400 -6400 15420 -6330
rect 15490 -6400 15510 -6330
rect 15580 -6400 15600 -6330
rect 15670 -6400 15690 -6330
rect 15760 -6400 15780 -6330
rect 15850 -6400 15870 -6330
rect 15940 -6400 16130 -6330
rect 14520 -6420 16130 -6400
rect 14520 -6490 14700 -6420
rect 14770 -6490 14790 -6420
rect 14860 -6490 14880 -6420
rect 14950 -6490 14970 -6420
rect 15040 -6490 15060 -6420
rect 15130 -6490 15150 -6420
rect 15220 -6490 15240 -6420
rect 15310 -6490 15330 -6420
rect 15400 -6490 15420 -6420
rect 15490 -6490 15510 -6420
rect 15580 -6490 15600 -6420
rect 15670 -6490 15690 -6420
rect 15760 -6490 15780 -6420
rect 15850 -6490 15870 -6420
rect 15940 -6490 16130 -6420
rect 31100 -4700 38190 -4630
rect 38260 -4700 38280 -4630
rect 38350 -4700 38370 -4630
rect 38440 -4700 38500 -4630
rect 31100 -4720 38500 -4700
rect 31100 -4790 38190 -4720
rect 38260 -4790 38280 -4720
rect 38350 -4790 38370 -4720
rect 38440 -4790 38500 -4720
rect 31100 -4810 38500 -4790
rect 31100 -4880 38190 -4810
rect 38260 -4880 38280 -4810
rect 38350 -4880 38370 -4810
rect 38440 -4880 38500 -4810
rect 31100 -4900 38500 -4880
rect 31100 -4970 38190 -4900
rect 38260 -4970 38280 -4900
rect 38350 -4970 38370 -4900
rect 38440 -4970 38500 -4900
rect 31100 -4990 38500 -4970
rect 31100 -5060 38190 -4990
rect 38260 -5060 38280 -4990
rect 38350 -5060 38370 -4990
rect 38440 -5060 38500 -4990
rect 31100 -5080 38500 -5060
rect 31100 -5150 38190 -5080
rect 38260 -5150 38280 -5080
rect 38350 -5150 38370 -5080
rect 38440 -5150 38500 -5080
rect 31100 -5170 38500 -5150
rect 31100 -5240 38190 -5170
rect 38260 -5240 38280 -5170
rect 38350 -5240 38370 -5170
rect 38440 -5240 38500 -5170
rect 31100 -5260 38500 -5240
rect 31100 -5330 38190 -5260
rect 38260 -5330 38280 -5260
rect 38350 -5330 38370 -5260
rect 38440 -5330 38500 -5260
rect 31100 -5350 38500 -5330
rect 31100 -5420 38190 -5350
rect 38260 -5420 38280 -5350
rect 38350 -5420 38370 -5350
rect 38440 -5420 38500 -5350
rect 31100 -5440 38500 -5420
rect 31100 -5510 38190 -5440
rect 38260 -5510 38280 -5440
rect 38350 -5510 38370 -5440
rect 38440 -5510 38500 -5440
rect 31100 -5530 38500 -5510
rect 31100 -5600 38190 -5530
rect 38260 -5600 38280 -5530
rect 38350 -5600 38370 -5530
rect 38440 -5600 38500 -5530
rect 31100 -5620 38500 -5600
rect 31100 -5690 38190 -5620
rect 38260 -5690 38280 -5620
rect 38350 -5690 38370 -5620
rect 38440 -5690 38500 -5620
rect 31100 -5710 38500 -5690
rect 31100 -5780 38190 -5710
rect 38260 -5780 38280 -5710
rect 38350 -5780 38370 -5710
rect 38440 -5780 38500 -5710
rect 31100 -5800 38500 -5780
rect 31100 -5870 38190 -5800
rect 38260 -5870 38280 -5800
rect 38350 -5870 38370 -5800
rect 38440 -5870 38500 -5800
rect 31100 -5890 38500 -5870
rect 31100 -5960 38190 -5890
rect 38260 -5960 38280 -5890
rect 38350 -5960 38370 -5890
rect 38440 -5960 38500 -5890
rect 31100 -5980 38500 -5960
rect 31100 -6050 38190 -5980
rect 38260 -6050 38280 -5980
rect 38350 -6050 38370 -5980
rect 38440 -6050 38500 -5980
rect 31100 -6070 38500 -6050
rect 31100 -6140 38190 -6070
rect 38260 -6140 38280 -6070
rect 38350 -6140 38370 -6070
rect 38440 -6140 38500 -6070
rect 31100 -6160 38500 -6140
rect 31100 -6230 38190 -6160
rect 38260 -6230 38280 -6160
rect 38350 -6230 38370 -6160
rect 38440 -6230 38500 -6160
rect 31100 -6250 38500 -6230
rect 31100 -6320 38190 -6250
rect 38260 -6320 38280 -6250
rect 38350 -6320 38370 -6250
rect 38440 -6320 38500 -6250
rect 31100 -6340 38500 -6320
rect 31100 -6410 38190 -6340
rect 38260 -6410 38280 -6340
rect 38350 -6410 38370 -6340
rect 38440 -6410 38500 -6340
rect 31100 -6450 38500 -6410
rect 14520 -6510 16130 -6490
rect 14520 -6580 14700 -6510
rect 14770 -6580 14790 -6510
rect 14860 -6580 14880 -6510
rect 14950 -6580 14970 -6510
rect 15040 -6580 15060 -6510
rect 15130 -6580 15150 -6510
rect 15220 -6580 15240 -6510
rect 15310 -6580 15330 -6510
rect 15400 -6580 15420 -6510
rect 15490 -6580 15510 -6510
rect 15580 -6580 15600 -6510
rect 15670 -6580 15690 -6510
rect 15760 -6580 15780 -6510
rect 15850 -6580 15870 -6510
rect 15940 -6580 16130 -6510
rect 14520 -6640 16130 -6580
rect 16380 -6520 16520 -6470
rect 16380 -6590 16420 -6520
rect 16490 -6590 16520 -6520
rect 16380 -6630 16520 -6590
rect 16380 -6640 16420 -6630
rect 7560 -6720 7590 -6660
rect 7650 -6720 7690 -6660
rect 7750 -6720 7790 -6660
rect 7850 -6720 8490 -6660
rect 7560 -6760 8490 -6720
rect 7560 -6820 7590 -6760
rect 7650 -6820 7690 -6760
rect 7750 -6820 7790 -6760
rect 7850 -6820 8490 -6760
rect 7560 -6850 8490 -6820
rect 8710 -6670 16420 -6640
rect 8710 -6730 9870 -6670
rect 9930 -6730 9970 -6670
rect 10030 -6730 10070 -6670
rect 10130 -6700 16420 -6670
rect 16490 -6700 16520 -6630
rect 10130 -6730 16520 -6700
rect 8710 -6740 16520 -6730
rect 8710 -6770 16420 -6740
rect 8710 -6830 9870 -6770
rect 9930 -6830 9970 -6770
rect 10030 -6830 10070 -6770
rect 10130 -6810 16420 -6770
rect 16490 -6810 16520 -6740
rect 10130 -6830 16520 -6810
rect 8710 -6850 16520 -6830
rect -1740 -6920 -1710 -6850
rect -1640 -6870 6190 -6850
rect -1640 -6920 4770 -6870
rect -1740 -6930 4770 -6920
rect 4830 -6930 4870 -6870
rect 4930 -6930 4970 -6870
rect 5030 -6930 6190 -6870
rect -1740 -6950 6190 -6930
rect 5880 -9620 6190 -6950
rect -270 -9660 6190 -9620
rect -270 -9730 -240 -9660
rect -170 -9730 -130 -9660
rect -60 -9730 -20 -9660
rect 50 -9730 90 -9660
rect 160 -9730 6190 -9660
rect -270 -9790 6190 -9730
rect -270 -9860 -240 -9790
rect -170 -9860 -130 -9790
rect -60 -9860 -20 -9790
rect 50 -9860 90 -9790
rect 160 -9860 6190 -9790
rect -270 -9900 6190 -9860
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1330 -10410 1370 -10340
rect 1440 -10410 1480 -10340
rect 1550 -10410 1590 -10340
rect 1660 -10410 1700 -10340
rect 1770 -10410 1810 -10340
rect 1880 -10410 1920 -10340
rect 1990 -10410 2030 -10340
rect 2100 -10410 2140 -10340
rect 2210 -10410 2250 -10340
rect 2320 -10410 2360 -10340
rect 2430 -10410 2470 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1330 -10520 1370 -10450
rect 1440 -10520 1480 -10450
rect 1550 -10520 1590 -10450
rect 1660 -10520 1700 -10450
rect 1770 -10520 1810 -10450
rect 1880 -10520 1920 -10450
rect 1990 -10520 2030 -10450
rect 2100 -10520 2140 -10450
rect 2210 -10520 2250 -10450
rect 2320 -10520 2360 -10450
rect 2430 -10520 2470 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10570 2680 -10520
rect 2210 -12300 3810 -12250
rect 2210 -12370 2240 -12300
rect 2310 -12370 2350 -12300
rect 2420 -12370 2460 -12300
rect 2530 -12370 2570 -12300
rect 2640 -12370 2680 -12300
rect 2750 -12370 2790 -12300
rect 2860 -12370 2900 -12300
rect 2970 -12370 3010 -12300
rect 3080 -12370 3120 -12300
rect 3190 -12370 3230 -12300
rect 3300 -12370 3340 -12300
rect 3410 -12370 3450 -12300
rect 3520 -12370 3560 -12300
rect 3630 -12370 3670 -12300
rect 3740 -12370 3810 -12300
rect 2210 -12410 3810 -12370
rect 2210 -12480 2240 -12410
rect 2310 -12480 2350 -12410
rect 2420 -12480 2460 -12410
rect 2530 -12480 2570 -12410
rect 2640 -12480 2680 -12410
rect 2750 -12480 2790 -12410
rect 2860 -12480 2900 -12410
rect 2970 -12480 3010 -12410
rect 3080 -12480 3120 -12410
rect 3190 -12480 3230 -12410
rect 3300 -12480 3340 -12410
rect 3410 -12480 3450 -12410
rect 3520 -12480 3560 -12410
rect 3630 -12480 3670 -12410
rect 3740 -12480 3810 -12410
rect 2210 -12510 3810 -12480
rect 5880 -13220 6190 -9900
rect 8710 -6870 16420 -6850
rect 8710 -6930 9870 -6870
rect 9930 -6930 9970 -6870
rect 10030 -6930 10070 -6870
rect 10130 -6920 16420 -6870
rect 16490 -6920 16520 -6850
rect 10130 -6930 16520 -6920
rect 8710 -6950 16520 -6930
rect 8710 -9620 9020 -6950
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8340 14900 -8300
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 14900 -8340
rect 14590 -8450 14900 -8410
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 21610 -8360 21930 -8330
rect 21610 -8430 21630 -8360
rect 21700 -8430 21730 -8360
rect 21800 -8430 21830 -8360
rect 21900 -8430 21930 -8360
rect 21610 -8460 21930 -8430
rect 21610 -8530 21630 -8460
rect 21700 -8530 21730 -8460
rect 21800 -8530 21830 -8460
rect 21900 -8530 21930 -8460
rect 21610 -8560 21930 -8530
rect 21610 -8630 21630 -8560
rect 21700 -8630 21730 -8560
rect 21800 -8630 21830 -8560
rect 21900 -8630 21930 -8560
rect 21610 -8650 21930 -8630
rect 22630 -9010 22950 -8980
rect 22630 -9080 22650 -9010
rect 22720 -9080 22750 -9010
rect 22820 -9080 22850 -9010
rect 22920 -9080 22950 -9010
rect 22630 -9110 22950 -9080
rect 22630 -9180 22650 -9110
rect 22720 -9180 22750 -9110
rect 22820 -9180 22850 -9110
rect 22920 -9180 22950 -9110
rect 22630 -9210 22950 -9180
rect 22630 -9280 22650 -9210
rect 22720 -9280 22750 -9210
rect 22820 -9280 22850 -9210
rect 22920 -9280 22950 -9210
rect 22630 -9300 22950 -9280
rect 8710 -9660 15170 -9620
rect 8710 -9730 14720 -9660
rect 14790 -9730 14830 -9660
rect 14900 -9730 14940 -9660
rect 15010 -9730 15050 -9660
rect 15120 -9730 15170 -9660
rect 8710 -9790 15170 -9730
rect 8710 -9860 14720 -9790
rect 14790 -9860 14830 -9790
rect 14900 -9860 14940 -9790
rect 15010 -9860 15050 -9790
rect 15120 -9860 15170 -9790
rect 8710 -9900 15170 -9860
rect 8710 -13220 9020 -9900
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12470 -10440 12510 -10370
rect 12580 -10440 12620 -10370
rect 12690 -10440 12730 -10370
rect 12800 -10440 12840 -10370
rect 12910 -10440 12950 -10370
rect 13020 -10440 13060 -10370
rect 13130 -10440 13170 -10370
rect 13240 -10440 13280 -10370
rect 13350 -10440 13390 -10370
rect 13460 -10440 13500 -10370
rect 13570 -10440 13610 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12470 -10550 12510 -10480
rect 12580 -10550 12620 -10480
rect 12690 -10550 12730 -10480
rect 12800 -10550 12840 -10480
rect 12910 -10550 12950 -10480
rect 13020 -10550 13060 -10480
rect 13130 -10550 13170 -10480
rect 13240 -10550 13280 -10480
rect 13350 -10550 13390 -10480
rect 13460 -10550 13500 -10480
rect 13570 -10550 13610 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10600 13820 -10550
rect 29960 -10520 30790 -10510
rect 29960 -10590 29990 -10520
rect 30060 -10590 30700 -10520
rect 30770 -10590 30790 -10520
rect 29960 -10630 30790 -10590
rect 29960 -10700 29990 -10630
rect 30060 -10700 30700 -10630
rect 30770 -10700 30790 -10630
rect 29960 -10740 30790 -10700
rect 29960 -10810 29990 -10740
rect 30060 -10810 30700 -10740
rect 30770 -10810 30790 -10740
rect 29960 -10830 30790 -10810
rect 11090 -12300 12690 -12250
rect 11090 -12370 11120 -12300
rect 11190 -12370 11230 -12300
rect 11300 -12370 11340 -12300
rect 11410 -12370 11450 -12300
rect 11520 -12370 11560 -12300
rect 11630 -12370 11670 -12300
rect 11740 -12370 11780 -12300
rect 11850 -12370 11890 -12300
rect 11960 -12370 12000 -12300
rect 12070 -12370 12110 -12300
rect 12180 -12370 12220 -12300
rect 12290 -12370 12330 -12300
rect 12400 -12370 12440 -12300
rect 12510 -12370 12550 -12300
rect 12620 -12370 12690 -12300
rect 11090 -12410 12690 -12370
rect 11090 -12480 11120 -12410
rect 11190 -12480 11230 -12410
rect 11300 -12480 11340 -12410
rect 11410 -12480 11450 -12410
rect 11520 -12480 11560 -12410
rect 11630 -12480 11670 -12410
rect 11740 -12480 11780 -12410
rect 11850 -12480 11890 -12410
rect 11960 -12480 12000 -12410
rect 12070 -12480 12110 -12410
rect 12180 -12480 12220 -12410
rect 12290 -12480 12330 -12410
rect 12400 -12480 12440 -12410
rect 12510 -12480 12550 -12410
rect 12620 -12480 12690 -12410
rect 11090 -12510 12690 -12480
rect 5880 -13250 7310 -13220
rect 5880 -13310 7010 -13250
rect 7070 -13310 7110 -13250
rect 7170 -13310 7210 -13250
rect 7270 -13310 7310 -13250
rect 5880 -13340 7310 -13310
rect 5880 -13400 7010 -13340
rect 7070 -13400 7110 -13340
rect 7170 -13400 7210 -13340
rect 7270 -13400 7310 -13340
rect 5880 -13430 7310 -13400
rect 5880 -13490 7010 -13430
rect 7070 -13490 7110 -13430
rect 7170 -13490 7210 -13430
rect 7270 -13490 7310 -13430
rect 5880 -13530 7310 -13490
rect 5880 -13590 7010 -13530
rect 7070 -13590 7110 -13530
rect 7170 -13590 7210 -13530
rect 7270 -13590 7310 -13530
rect 5880 -13620 7310 -13590
rect 5880 -13680 7010 -13620
rect 7070 -13680 7110 -13620
rect 7170 -13680 7210 -13620
rect 7270 -13680 7310 -13620
rect 5880 -13710 7310 -13680
rect 5880 -13770 7010 -13710
rect 7070 -13770 7110 -13710
rect 7170 -13770 7210 -13710
rect 7270 -13770 7310 -13710
rect 5880 -13800 7310 -13770
rect 7590 -13250 9020 -13220
rect 7590 -13310 7630 -13250
rect 7690 -13310 7730 -13250
rect 7790 -13310 7830 -13250
rect 7890 -13310 9020 -13250
rect 7590 -13340 9020 -13310
rect 7590 -13400 7630 -13340
rect 7690 -13400 7730 -13340
rect 7790 -13400 7830 -13340
rect 7890 -13400 9020 -13340
rect 7590 -13430 9020 -13400
rect 7590 -13490 7630 -13430
rect 7690 -13490 7730 -13430
rect 7790 -13490 7830 -13430
rect 7890 -13490 9020 -13430
rect 7590 -13530 9020 -13490
rect 7590 -13590 7630 -13530
rect 7690 -13590 7730 -13530
rect 7790 -13590 7830 -13530
rect 7890 -13590 9020 -13530
rect 7590 -13620 9020 -13590
rect 7590 -13680 7630 -13620
rect 7690 -13680 7730 -13620
rect 7790 -13680 7830 -13620
rect 7890 -13680 9020 -13620
rect 7590 -13710 9020 -13680
rect 7590 -13770 7630 -13710
rect 7690 -13770 7730 -13710
rect 7790 -13770 7830 -13710
rect 7890 -13770 9020 -13710
rect 7590 -13800 9020 -13770
rect 21610 -14020 21930 -13990
rect 21610 -14090 21630 -14020
rect 21700 -14090 21730 -14020
rect 21800 -14090 21830 -14020
rect 21900 -14090 21930 -14020
rect 21610 -14120 21930 -14090
rect 21610 -14190 21630 -14120
rect 21700 -14190 21730 -14120
rect 21800 -14190 21830 -14120
rect 21900 -14190 21930 -14120
rect 21610 -14220 21930 -14190
rect 21610 -14290 21630 -14220
rect 21700 -14290 21730 -14220
rect 21800 -14290 21830 -14220
rect 21900 -14290 21930 -14220
rect 21610 -14310 21930 -14290
rect 22900 -14870 23220 -14840
rect 22900 -14940 22920 -14870
rect 22990 -14940 23020 -14870
rect 23090 -14940 23120 -14870
rect 23190 -14940 23220 -14870
rect 22900 -14970 23220 -14940
rect 22900 -15040 22920 -14970
rect 22990 -15040 23020 -14970
rect 23090 -15040 23120 -14970
rect 23190 -15040 23220 -14970
rect 22900 -15070 23220 -15040
rect 22900 -15140 22920 -15070
rect 22990 -15140 23020 -15070
rect 23090 -15140 23120 -15070
rect 23190 -15140 23220 -15070
rect 22900 -15160 23220 -15140
rect 5010 -17100 5330 -17070
rect 5010 -17160 5040 -17100
rect 5100 -17160 5140 -17100
rect 5200 -17160 5240 -17100
rect 5300 -17160 5330 -17100
rect 5010 -17200 5330 -17160
rect 5010 -17260 5040 -17200
rect 5100 -17260 5140 -17200
rect 5200 -17260 5240 -17200
rect 5300 -17260 5330 -17200
rect 5010 -17300 5330 -17260
rect 5010 -17360 5040 -17300
rect 5100 -17360 5140 -17300
rect 5200 -17360 5240 -17300
rect 5300 -17360 5330 -17300
rect 2210 -22660 3810 -22630
rect 2210 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2460 -22730 2500 -22660
rect 2570 -22730 2610 -22660
rect 2680 -22730 2720 -22660
rect 2790 -22730 2830 -22660
rect 2900 -22730 2940 -22660
rect 3010 -22730 3050 -22660
rect 3120 -22730 3160 -22660
rect 3230 -22730 3270 -22660
rect 3340 -22730 3380 -22660
rect 3450 -22730 3490 -22660
rect 3560 -22730 3600 -22660
rect 3670 -22730 3710 -22660
rect 3780 -22730 3810 -22660
rect 2210 -22770 3810 -22730
rect 2210 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2460 -22840 2500 -22770
rect 2570 -22840 2610 -22770
rect 2680 -22840 2720 -22770
rect 2790 -22840 2830 -22770
rect 2900 -22840 2940 -22770
rect 3010 -22840 3050 -22770
rect 3120 -22840 3160 -22770
rect 3230 -22840 3270 -22770
rect 3340 -22840 3380 -22770
rect 3450 -22840 3490 -22770
rect 3560 -22840 3600 -22770
rect 3670 -22840 3710 -22770
rect 3780 -22840 3810 -22770
rect 2210 -22890 3810 -22840
rect 5010 -24030 5330 -17360
rect 9570 -17100 9890 -17070
rect 9570 -17160 9600 -17100
rect 9660 -17160 9700 -17100
rect 9760 -17160 9800 -17100
rect 9860 -17160 9890 -17100
rect 9570 -17200 9890 -17160
rect 9570 -17260 9600 -17200
rect 9660 -17260 9700 -17200
rect 9760 -17260 9800 -17200
rect 9860 -17260 9890 -17200
rect 9570 -17300 9890 -17260
rect 9570 -17360 9600 -17300
rect 9660 -17360 9700 -17300
rect 9760 -17360 9800 -17300
rect 9860 -17360 9890 -17300
rect 7210 -17600 7650 -17580
rect 7210 -17670 7230 -17600
rect 7300 -17670 7340 -17600
rect 7410 -17670 7450 -17600
rect 7520 -17670 7560 -17600
rect 7630 -17670 7650 -17600
rect 7210 -17710 7650 -17670
rect 7210 -17780 7230 -17710
rect 7300 -17780 7340 -17710
rect 7410 -17780 7450 -17710
rect 7520 -17780 7560 -17710
rect 7630 -17780 7650 -17710
rect 7210 -17820 7650 -17780
rect 7210 -17890 7230 -17820
rect 7300 -17890 7340 -17820
rect 7410 -17890 7450 -17820
rect 7520 -17890 7560 -17820
rect 7630 -17890 7650 -17820
rect 7210 -17930 7650 -17890
rect 7210 -18000 7230 -17930
rect 7300 -18000 7340 -17930
rect 7410 -18000 7450 -17930
rect 7520 -18000 7560 -17930
rect 7630 -18000 7650 -17930
rect 7210 -18020 7650 -18000
rect 9570 -24030 9890 -17360
rect 21610 -20100 21930 -20070
rect 21610 -20170 21630 -20100
rect 21700 -20170 21730 -20100
rect 21800 -20170 21830 -20100
rect 21900 -20170 21930 -20100
rect 21610 -20200 21930 -20170
rect 21610 -20270 21630 -20200
rect 21700 -20270 21730 -20200
rect 21800 -20270 21830 -20200
rect 21900 -20270 21930 -20200
rect 21610 -20300 21930 -20270
rect 21610 -20370 21630 -20300
rect 21700 -20370 21730 -20300
rect 21800 -20370 21830 -20300
rect 21900 -20370 21930 -20300
rect 21610 -20390 21930 -20370
rect 22680 -20730 23000 -20700
rect 22680 -20800 22700 -20730
rect 22770 -20800 22800 -20730
rect 22870 -20800 22900 -20730
rect 22970 -20800 23000 -20730
rect 22680 -20830 23000 -20800
rect 22680 -20900 22700 -20830
rect 22770 -20900 22800 -20830
rect 22870 -20900 22900 -20830
rect 22970 -20900 23000 -20830
rect 22680 -20930 23000 -20900
rect 22680 -21000 22700 -20930
rect 22770 -21000 22800 -20930
rect 22870 -21000 22900 -20930
rect 22970 -21000 23000 -20930
rect 22680 -21020 23000 -21000
rect 11090 -22660 12690 -22630
rect 11090 -22730 11160 -22660
rect 11230 -22730 11270 -22660
rect 11340 -22730 11380 -22660
rect 11450 -22730 11490 -22660
rect 11560 -22730 11600 -22660
rect 11670 -22730 11710 -22660
rect 11780 -22730 11820 -22660
rect 11890 -22730 11930 -22660
rect 12000 -22730 12040 -22660
rect 12110 -22730 12150 -22660
rect 12220 -22730 12260 -22660
rect 12330 -22730 12370 -22660
rect 12440 -22730 12480 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12690 -22660
rect 11090 -22770 12690 -22730
rect 11090 -22840 11160 -22770
rect 11230 -22840 11270 -22770
rect 11340 -22840 11380 -22770
rect 11450 -22840 11490 -22770
rect 11560 -22840 11600 -22770
rect 11670 -22840 11710 -22770
rect 11780 -22840 11820 -22770
rect 11890 -22840 11930 -22770
rect 12000 -22840 12040 -22770
rect 12110 -22840 12150 -22770
rect 12220 -22840 12260 -22770
rect 12330 -22840 12370 -22770
rect 12440 -22840 12480 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12690 -22770
rect 11090 -22890 12690 -22840
<< via3 >>
rect -4730 21510 -4660 21580
rect -4640 21510 -4570 21580
rect -4550 21510 -4480 21580
rect -4460 21510 -4390 21580
rect -4370 21510 -4300 21580
rect -4280 21510 -4210 21580
rect -4190 21510 -4120 21580
rect -4100 21510 -4030 21580
rect -4010 21510 -3940 21580
rect -3920 21510 -3850 21580
rect -3830 21510 -3760 21580
rect -3740 21510 -3670 21580
rect -3650 21510 -3580 21580
rect -3560 21510 -3490 21580
rect -3470 21510 -3400 21580
rect -3380 21510 -3310 21580
rect -3290 21510 -3220 21580
rect -3200 21510 -3130 21580
rect -3110 21510 -3040 21580
rect -3020 21510 -2950 21580
rect -2930 21510 -2860 21580
rect -2840 21510 -2770 21580
rect -2750 21510 -2680 21580
rect -2660 21510 -2590 21580
rect -2570 21510 -2500 21580
rect -2480 21510 -2410 21580
rect -2390 21510 -2320 21580
rect -2300 21510 -2230 21580
rect -2210 21510 -2140 21580
rect -2120 21510 -2050 21580
rect -2030 21510 -1960 21580
rect -1940 21510 -1870 21580
rect -1850 21510 -1780 21580
rect -1720 21510 -1650 21580
rect -1630 21510 -1560 21580
rect -1540 21510 -1470 21580
rect -1450 21510 -1380 21580
rect -1360 21510 -1290 21580
rect -1270 21510 -1200 21580
rect -1180 21510 -1110 21580
rect -1090 21510 -1020 21580
rect -1000 21510 -930 21580
rect -910 21510 -840 21580
rect -820 21510 -750 21580
rect -730 21510 -660 21580
rect -640 21510 -570 21580
rect -550 21510 -480 21580
rect -460 21510 -390 21580
rect -370 21510 -300 21580
rect -280 21510 -210 21580
rect -190 21510 -120 21580
rect -100 21510 -30 21580
rect -10 21510 60 21580
rect 80 21510 150 21580
rect 170 21510 240 21580
rect 260 21510 330 21580
rect 350 21510 420 21580
rect 440 21510 510 21580
rect 530 21510 600 21580
rect 620 21510 690 21580
rect 710 21510 780 21580
rect 800 21510 870 21580
rect 890 21510 960 21580
rect 980 21510 1050 21580
rect 1070 21510 1140 21580
rect 1160 21510 1230 21580
rect 1290 21510 1360 21580
rect 1380 21510 1450 21580
rect 1470 21510 1540 21580
rect 1560 21510 1630 21580
rect 1650 21510 1720 21580
rect 1740 21510 1810 21580
rect 1830 21510 1900 21580
rect 1920 21510 1990 21580
rect 2010 21510 2080 21580
rect 2100 21510 2170 21580
rect 2190 21510 2260 21580
rect 2280 21510 2350 21580
rect 2370 21510 2440 21580
rect 2460 21510 2530 21580
rect 2550 21510 2620 21580
rect 2640 21510 2710 21580
rect 2730 21510 2800 21580
rect 2820 21510 2890 21580
rect 2910 21510 2980 21580
rect 3000 21510 3070 21580
rect 3090 21510 3160 21580
rect 3180 21510 3250 21580
rect 3270 21510 3340 21580
rect 3360 21510 3430 21580
rect 3450 21510 3520 21580
rect 3540 21510 3610 21580
rect 3630 21510 3700 21580
rect 3720 21510 3790 21580
rect 3810 21510 3880 21580
rect 3900 21510 3970 21580
rect 3990 21510 4060 21580
rect 4080 21510 4150 21580
rect 4170 21510 4240 21580
rect 4300 21510 4370 21580
rect 4390 21510 4460 21580
rect 4480 21510 4550 21580
rect 4570 21510 4640 21580
rect 4660 21510 4730 21580
rect 4750 21510 4820 21580
rect 4840 21510 4910 21580
rect 4930 21510 5000 21580
rect 5020 21510 5090 21580
rect 5110 21510 5180 21580
rect 5200 21510 5270 21580
rect 5290 21510 5360 21580
rect 5380 21510 5450 21580
rect 5470 21510 5540 21580
rect 5560 21510 5630 21580
rect 5650 21510 5720 21580
rect 5740 21510 5810 21580
rect 5830 21510 5900 21580
rect 5920 21510 5990 21580
rect 6010 21510 6080 21580
rect 6100 21510 6170 21580
rect 6190 21510 6260 21580
rect 6280 21510 6350 21580
rect 6370 21510 6440 21580
rect 6460 21510 6530 21580
rect 6550 21510 6620 21580
rect 6640 21510 6710 21580
rect 6730 21510 6800 21580
rect 6820 21510 6890 21580
rect 6910 21510 6980 21580
rect 7000 21510 7070 21580
rect 7090 21510 7160 21580
rect 7180 21510 7250 21580
rect -4730 21420 -4660 21490
rect -4640 21420 -4570 21490
rect -4550 21420 -4480 21490
rect -4460 21420 -4390 21490
rect -4370 21420 -4300 21490
rect -4280 21420 -4210 21490
rect -4190 21420 -4120 21490
rect -4100 21420 -4030 21490
rect -4010 21420 -3940 21490
rect -3920 21420 -3850 21490
rect -3830 21420 -3760 21490
rect -3740 21420 -3670 21490
rect -3650 21420 -3580 21490
rect -3560 21420 -3490 21490
rect -3470 21420 -3400 21490
rect -3380 21420 -3310 21490
rect -3290 21420 -3220 21490
rect -3200 21420 -3130 21490
rect -3110 21420 -3040 21490
rect -3020 21420 -2950 21490
rect -2930 21420 -2860 21490
rect -2840 21420 -2770 21490
rect -2750 21420 -2680 21490
rect -2660 21420 -2590 21490
rect -2570 21420 -2500 21490
rect -2480 21420 -2410 21490
rect -2390 21420 -2320 21490
rect -2300 21420 -2230 21490
rect -2210 21420 -2140 21490
rect -2120 21420 -2050 21490
rect -2030 21420 -1960 21490
rect -1940 21420 -1870 21490
rect -1850 21420 -1780 21490
rect -1720 21420 -1650 21490
rect -1630 21420 -1560 21490
rect -1540 21420 -1470 21490
rect -1450 21420 -1380 21490
rect -1360 21420 -1290 21490
rect -1270 21420 -1200 21490
rect -1180 21420 -1110 21490
rect -1090 21420 -1020 21490
rect -1000 21420 -930 21490
rect -910 21420 -840 21490
rect -820 21420 -750 21490
rect -730 21420 -660 21490
rect -640 21420 -570 21490
rect -550 21420 -480 21490
rect -460 21420 -390 21490
rect -370 21420 -300 21490
rect -280 21420 -210 21490
rect -190 21420 -120 21490
rect -100 21420 -30 21490
rect -10 21420 60 21490
rect 80 21420 150 21490
rect 170 21420 240 21490
rect 260 21420 330 21490
rect 350 21420 420 21490
rect 440 21420 510 21490
rect 530 21420 600 21490
rect 620 21420 690 21490
rect 710 21420 780 21490
rect 800 21420 870 21490
rect 890 21420 960 21490
rect 980 21420 1050 21490
rect 1070 21420 1140 21490
rect 1160 21420 1230 21490
rect 1290 21420 1360 21490
rect 1380 21420 1450 21490
rect 1470 21420 1540 21490
rect 1560 21420 1630 21490
rect 1650 21420 1720 21490
rect 1740 21420 1810 21490
rect 1830 21420 1900 21490
rect 1920 21420 1990 21490
rect 2010 21420 2080 21490
rect 2100 21420 2170 21490
rect 2190 21420 2260 21490
rect 2280 21420 2350 21490
rect 2370 21420 2440 21490
rect 2460 21420 2530 21490
rect 2550 21420 2620 21490
rect 2640 21420 2710 21490
rect 2730 21420 2800 21490
rect 2820 21420 2890 21490
rect 2910 21420 2980 21490
rect 3000 21420 3070 21490
rect 3090 21420 3160 21490
rect 3180 21420 3250 21490
rect 3270 21420 3340 21490
rect 3360 21420 3430 21490
rect 3450 21420 3520 21490
rect 3540 21420 3610 21490
rect 3630 21420 3700 21490
rect 3720 21420 3790 21490
rect 3810 21420 3880 21490
rect 3900 21420 3970 21490
rect 3990 21420 4060 21490
rect 4080 21420 4150 21490
rect 4170 21420 4240 21490
rect 4300 21420 4370 21490
rect 4390 21420 4460 21490
rect 4480 21420 4550 21490
rect 4570 21420 4640 21490
rect 4660 21420 4730 21490
rect 4750 21420 4820 21490
rect 4840 21420 4910 21490
rect 4930 21420 5000 21490
rect 5020 21420 5090 21490
rect 5110 21420 5180 21490
rect 5200 21420 5270 21490
rect 5290 21420 5360 21490
rect 5380 21420 5450 21490
rect 5470 21420 5540 21490
rect 5560 21420 5630 21490
rect 5650 21420 5720 21490
rect 5740 21420 5810 21490
rect 5830 21420 5900 21490
rect 5920 21420 5990 21490
rect 6010 21420 6080 21490
rect 6100 21420 6170 21490
rect 6190 21420 6260 21490
rect 6280 21420 6350 21490
rect 6370 21420 6440 21490
rect 6460 21420 6530 21490
rect 6550 21420 6620 21490
rect 6640 21420 6710 21490
rect 6730 21420 6800 21490
rect 6820 21420 6890 21490
rect 6910 21420 6980 21490
rect 7000 21420 7070 21490
rect 7090 21420 7160 21490
rect 7180 21420 7250 21490
rect -4730 21330 -4660 21400
rect -4640 21330 -4570 21400
rect -4550 21330 -4480 21400
rect -4460 21330 -4390 21400
rect -4370 21330 -4300 21400
rect -4280 21330 -4210 21400
rect -4190 21330 -4120 21400
rect -4100 21330 -4030 21400
rect -4010 21330 -3940 21400
rect -3920 21330 -3850 21400
rect -3830 21330 -3760 21400
rect -3740 21330 -3670 21400
rect -3650 21330 -3580 21400
rect -3560 21330 -3490 21400
rect -3470 21330 -3400 21400
rect -3380 21330 -3310 21400
rect -3290 21330 -3220 21400
rect -3200 21330 -3130 21400
rect -3110 21330 -3040 21400
rect -3020 21330 -2950 21400
rect -2930 21330 -2860 21400
rect -2840 21330 -2770 21400
rect -2750 21330 -2680 21400
rect -2660 21330 -2590 21400
rect -2570 21330 -2500 21400
rect -2480 21330 -2410 21400
rect -2390 21330 -2320 21400
rect -2300 21330 -2230 21400
rect -2210 21330 -2140 21400
rect -2120 21330 -2050 21400
rect -2030 21330 -1960 21400
rect -1940 21330 -1870 21400
rect -1850 21330 -1780 21400
rect -1720 21330 -1650 21400
rect -1630 21330 -1560 21400
rect -1540 21330 -1470 21400
rect -1450 21330 -1380 21400
rect -1360 21330 -1290 21400
rect -1270 21330 -1200 21400
rect -1180 21330 -1110 21400
rect -1090 21330 -1020 21400
rect -1000 21330 -930 21400
rect -910 21330 -840 21400
rect -820 21330 -750 21400
rect -730 21330 -660 21400
rect -640 21330 -570 21400
rect -550 21330 -480 21400
rect -460 21330 -390 21400
rect -370 21330 -300 21400
rect -280 21330 -210 21400
rect -190 21330 -120 21400
rect -100 21330 -30 21400
rect -10 21330 60 21400
rect 80 21330 150 21400
rect 170 21330 240 21400
rect 260 21330 330 21400
rect 350 21330 420 21400
rect 440 21330 510 21400
rect 530 21330 600 21400
rect 620 21330 690 21400
rect 710 21330 780 21400
rect 800 21330 870 21400
rect 890 21330 960 21400
rect 980 21330 1050 21400
rect 1070 21330 1140 21400
rect 1160 21330 1230 21400
rect 1290 21330 1360 21400
rect 1380 21330 1450 21400
rect 1470 21330 1540 21400
rect 1560 21330 1630 21400
rect 1650 21330 1720 21400
rect 1740 21330 1810 21400
rect 1830 21330 1900 21400
rect 1920 21330 1990 21400
rect 2010 21330 2080 21400
rect 2100 21330 2170 21400
rect 2190 21330 2260 21400
rect 2280 21330 2350 21400
rect 2370 21330 2440 21400
rect 2460 21330 2530 21400
rect 2550 21330 2620 21400
rect 2640 21330 2710 21400
rect 2730 21330 2800 21400
rect 2820 21330 2890 21400
rect 2910 21330 2980 21400
rect 3000 21330 3070 21400
rect 3090 21330 3160 21400
rect 3180 21330 3250 21400
rect 3270 21330 3340 21400
rect 3360 21330 3430 21400
rect 3450 21330 3520 21400
rect 3540 21330 3610 21400
rect 3630 21330 3700 21400
rect 3720 21330 3790 21400
rect 3810 21330 3880 21400
rect 3900 21330 3970 21400
rect 3990 21330 4060 21400
rect 4080 21330 4150 21400
rect 4170 21330 4240 21400
rect 4300 21330 4370 21400
rect 4390 21330 4460 21400
rect 4480 21330 4550 21400
rect 4570 21330 4640 21400
rect 4660 21330 4730 21400
rect 4750 21330 4820 21400
rect 4840 21330 4910 21400
rect 4930 21330 5000 21400
rect 5020 21330 5090 21400
rect 5110 21330 5180 21400
rect 5200 21330 5270 21400
rect 5290 21330 5360 21400
rect 5380 21330 5450 21400
rect 5470 21330 5540 21400
rect 5560 21330 5630 21400
rect 5650 21330 5720 21400
rect 5740 21330 5810 21400
rect 5830 21330 5900 21400
rect 5920 21330 5990 21400
rect 6010 21330 6080 21400
rect 6100 21330 6170 21400
rect 6190 21330 6260 21400
rect 6280 21330 6350 21400
rect 6370 21330 6440 21400
rect 6460 21330 6530 21400
rect 6550 21330 6620 21400
rect 6640 21330 6710 21400
rect 6730 21330 6800 21400
rect 6820 21330 6890 21400
rect 6910 21330 6980 21400
rect 7000 21330 7070 21400
rect 7090 21330 7160 21400
rect 7180 21330 7250 21400
rect 7650 21510 7720 21580
rect 7740 21510 7810 21580
rect 7830 21510 7900 21580
rect 7920 21510 7990 21580
rect 8010 21510 8080 21580
rect 8100 21510 8170 21580
rect 8190 21510 8260 21580
rect 8280 21510 8350 21580
rect 8370 21510 8440 21580
rect 8460 21510 8530 21580
rect 8550 21510 8620 21580
rect 8640 21510 8710 21580
rect 8730 21510 8800 21580
rect 8820 21510 8890 21580
rect 8910 21510 8980 21580
rect 9000 21510 9070 21580
rect 9090 21510 9160 21580
rect 9180 21510 9250 21580
rect 9270 21510 9340 21580
rect 9360 21510 9430 21580
rect 9450 21510 9520 21580
rect 9540 21510 9610 21580
rect 9630 21510 9700 21580
rect 9720 21510 9790 21580
rect 9810 21510 9880 21580
rect 9900 21510 9970 21580
rect 9990 21510 10060 21580
rect 10080 21510 10150 21580
rect 10170 21510 10240 21580
rect 10260 21510 10330 21580
rect 10350 21510 10420 21580
rect 10440 21510 10510 21580
rect 10530 21510 10600 21580
rect 10660 21510 10730 21580
rect 10750 21510 10820 21580
rect 10840 21510 10910 21580
rect 10930 21510 11000 21580
rect 11020 21510 11090 21580
rect 11110 21510 11180 21580
rect 11200 21510 11270 21580
rect 11290 21510 11360 21580
rect 11380 21510 11450 21580
rect 11470 21510 11540 21580
rect 11560 21510 11630 21580
rect 11650 21510 11720 21580
rect 11740 21510 11810 21580
rect 11830 21510 11900 21580
rect 11920 21510 11990 21580
rect 12010 21510 12080 21580
rect 12100 21510 12170 21580
rect 12190 21510 12260 21580
rect 12280 21510 12350 21580
rect 12370 21510 12440 21580
rect 12460 21510 12530 21580
rect 12550 21510 12620 21580
rect 12640 21510 12710 21580
rect 12730 21510 12800 21580
rect 12820 21510 12890 21580
rect 12910 21510 12980 21580
rect 13000 21510 13070 21580
rect 13090 21510 13160 21580
rect 13180 21510 13250 21580
rect 13270 21510 13340 21580
rect 13360 21510 13430 21580
rect 13450 21510 13520 21580
rect 13540 21510 13610 21580
rect 13670 21510 13740 21580
rect 13760 21510 13830 21580
rect 13850 21510 13920 21580
rect 13940 21510 14010 21580
rect 14030 21510 14100 21580
rect 14120 21510 14190 21580
rect 14210 21510 14280 21580
rect 14300 21510 14370 21580
rect 14390 21510 14460 21580
rect 14480 21510 14550 21580
rect 14570 21510 14640 21580
rect 14660 21510 14730 21580
rect 14750 21510 14820 21580
rect 14840 21510 14910 21580
rect 14930 21510 15000 21580
rect 15020 21510 15090 21580
rect 15110 21510 15180 21580
rect 15200 21510 15270 21580
rect 15290 21510 15360 21580
rect 15380 21510 15450 21580
rect 15470 21510 15540 21580
rect 15560 21510 15630 21580
rect 15650 21510 15720 21580
rect 15740 21510 15810 21580
rect 15830 21510 15900 21580
rect 15920 21510 15990 21580
rect 16010 21510 16080 21580
rect 16100 21510 16170 21580
rect 16190 21510 16260 21580
rect 16280 21510 16350 21580
rect 16370 21510 16440 21580
rect 16460 21510 16530 21580
rect 16550 21510 16620 21580
rect 16680 21510 16750 21580
rect 16770 21510 16840 21580
rect 16860 21510 16930 21580
rect 16950 21510 17020 21580
rect 17040 21510 17110 21580
rect 17130 21510 17200 21580
rect 17220 21510 17290 21580
rect 17310 21510 17380 21580
rect 17400 21510 17470 21580
rect 17490 21510 17560 21580
rect 17580 21510 17650 21580
rect 17670 21510 17740 21580
rect 17760 21510 17830 21580
rect 17850 21510 17920 21580
rect 17940 21510 18010 21580
rect 18030 21510 18100 21580
rect 18120 21510 18190 21580
rect 18210 21510 18280 21580
rect 18300 21510 18370 21580
rect 18390 21510 18460 21580
rect 18480 21510 18550 21580
rect 18570 21510 18640 21580
rect 18660 21510 18730 21580
rect 18750 21510 18820 21580
rect 18840 21510 18910 21580
rect 18930 21510 19000 21580
rect 19020 21510 19090 21580
rect 19110 21510 19180 21580
rect 19200 21510 19270 21580
rect 19290 21510 19360 21580
rect 19380 21510 19450 21580
rect 19470 21510 19540 21580
rect 19560 21510 19630 21580
rect 7650 21420 7720 21490
rect 7740 21420 7810 21490
rect 7830 21420 7900 21490
rect 7920 21420 7990 21490
rect 8010 21420 8080 21490
rect 8100 21420 8170 21490
rect 8190 21420 8260 21490
rect 8280 21420 8350 21490
rect 8370 21420 8440 21490
rect 8460 21420 8530 21490
rect 8550 21420 8620 21490
rect 8640 21420 8710 21490
rect 8730 21420 8800 21490
rect 8820 21420 8890 21490
rect 8910 21420 8980 21490
rect 9000 21420 9070 21490
rect 9090 21420 9160 21490
rect 9180 21420 9250 21490
rect 9270 21420 9340 21490
rect 9360 21420 9430 21490
rect 9450 21420 9520 21490
rect 9540 21420 9610 21490
rect 9630 21420 9700 21490
rect 9720 21420 9790 21490
rect 9810 21420 9880 21490
rect 9900 21420 9970 21490
rect 9990 21420 10060 21490
rect 10080 21420 10150 21490
rect 10170 21420 10240 21490
rect 10260 21420 10330 21490
rect 10350 21420 10420 21490
rect 10440 21420 10510 21490
rect 10530 21420 10600 21490
rect 10660 21420 10730 21490
rect 10750 21420 10820 21490
rect 10840 21420 10910 21490
rect 10930 21420 11000 21490
rect 11020 21420 11090 21490
rect 11110 21420 11180 21490
rect 11200 21420 11270 21490
rect 11290 21420 11360 21490
rect 11380 21420 11450 21490
rect 11470 21420 11540 21490
rect 11560 21420 11630 21490
rect 11650 21420 11720 21490
rect 11740 21420 11810 21490
rect 11830 21420 11900 21490
rect 11920 21420 11990 21490
rect 12010 21420 12080 21490
rect 12100 21420 12170 21490
rect 12190 21420 12260 21490
rect 12280 21420 12350 21490
rect 12370 21420 12440 21490
rect 12460 21420 12530 21490
rect 12550 21420 12620 21490
rect 12640 21420 12710 21490
rect 12730 21420 12800 21490
rect 12820 21420 12890 21490
rect 12910 21420 12980 21490
rect 13000 21420 13070 21490
rect 13090 21420 13160 21490
rect 13180 21420 13250 21490
rect 13270 21420 13340 21490
rect 13360 21420 13430 21490
rect 13450 21420 13520 21490
rect 13540 21420 13610 21490
rect 13670 21420 13740 21490
rect 13760 21420 13830 21490
rect 13850 21420 13920 21490
rect 13940 21420 14010 21490
rect 14030 21420 14100 21490
rect 14120 21420 14190 21490
rect 14210 21420 14280 21490
rect 14300 21420 14370 21490
rect 14390 21420 14460 21490
rect 14480 21420 14550 21490
rect 14570 21420 14640 21490
rect 14660 21420 14730 21490
rect 14750 21420 14820 21490
rect 14840 21420 14910 21490
rect 14930 21420 15000 21490
rect 15020 21420 15090 21490
rect 15110 21420 15180 21490
rect 15200 21420 15270 21490
rect 15290 21420 15360 21490
rect 15380 21420 15450 21490
rect 15470 21420 15540 21490
rect 15560 21420 15630 21490
rect 15650 21420 15720 21490
rect 15740 21420 15810 21490
rect 15830 21420 15900 21490
rect 15920 21420 15990 21490
rect 16010 21420 16080 21490
rect 16100 21420 16170 21490
rect 16190 21420 16260 21490
rect 16280 21420 16350 21490
rect 16370 21420 16440 21490
rect 16460 21420 16530 21490
rect 16550 21420 16620 21490
rect 16680 21420 16750 21490
rect 16770 21420 16840 21490
rect 16860 21420 16930 21490
rect 16950 21420 17020 21490
rect 17040 21420 17110 21490
rect 17130 21420 17200 21490
rect 17220 21420 17290 21490
rect 17310 21420 17380 21490
rect 17400 21420 17470 21490
rect 17490 21420 17560 21490
rect 17580 21420 17650 21490
rect 17670 21420 17740 21490
rect 17760 21420 17830 21490
rect 17850 21420 17920 21490
rect 17940 21420 18010 21490
rect 18030 21420 18100 21490
rect 18120 21420 18190 21490
rect 18210 21420 18280 21490
rect 18300 21420 18370 21490
rect 18390 21420 18460 21490
rect 18480 21420 18550 21490
rect 18570 21420 18640 21490
rect 18660 21420 18730 21490
rect 18750 21420 18820 21490
rect 18840 21420 18910 21490
rect 18930 21420 19000 21490
rect 19020 21420 19090 21490
rect 19110 21420 19180 21490
rect 19200 21420 19270 21490
rect 19290 21420 19360 21490
rect 19380 21420 19450 21490
rect 19470 21420 19540 21490
rect 19560 21420 19630 21490
rect 7650 21330 7720 21400
rect 7740 21330 7810 21400
rect 7830 21330 7900 21400
rect 7920 21330 7990 21400
rect 8010 21330 8080 21400
rect 8100 21330 8170 21400
rect 8190 21330 8260 21400
rect 8280 21330 8350 21400
rect 8370 21330 8440 21400
rect 8460 21330 8530 21400
rect 8550 21330 8620 21400
rect 8640 21330 8710 21400
rect 8730 21330 8800 21400
rect 8820 21330 8890 21400
rect 8910 21330 8980 21400
rect 9000 21330 9070 21400
rect 9090 21330 9160 21400
rect 9180 21330 9250 21400
rect 9270 21330 9340 21400
rect 9360 21330 9430 21400
rect 9450 21330 9520 21400
rect 9540 21330 9610 21400
rect 9630 21330 9700 21400
rect 9720 21330 9790 21400
rect 9810 21330 9880 21400
rect 9900 21330 9970 21400
rect 9990 21330 10060 21400
rect 10080 21330 10150 21400
rect 10170 21330 10240 21400
rect 10260 21330 10330 21400
rect 10350 21330 10420 21400
rect 10440 21330 10510 21400
rect 10530 21330 10600 21400
rect 10660 21330 10730 21400
rect 10750 21330 10820 21400
rect 10840 21330 10910 21400
rect 10930 21330 11000 21400
rect 11020 21330 11090 21400
rect 11110 21330 11180 21400
rect 11200 21330 11270 21400
rect 11290 21330 11360 21400
rect 11380 21330 11450 21400
rect 11470 21330 11540 21400
rect 11560 21330 11630 21400
rect 11650 21330 11720 21400
rect 11740 21330 11810 21400
rect 11830 21330 11900 21400
rect 11920 21330 11990 21400
rect 12010 21330 12080 21400
rect 12100 21330 12170 21400
rect 12190 21330 12260 21400
rect 12280 21330 12350 21400
rect 12370 21330 12440 21400
rect 12460 21330 12530 21400
rect 12550 21330 12620 21400
rect 12640 21330 12710 21400
rect 12730 21330 12800 21400
rect 12820 21330 12890 21400
rect 12910 21330 12980 21400
rect 13000 21330 13070 21400
rect 13090 21330 13160 21400
rect 13180 21330 13250 21400
rect 13270 21330 13340 21400
rect 13360 21330 13430 21400
rect 13450 21330 13520 21400
rect 13540 21330 13610 21400
rect 13670 21330 13740 21400
rect 13760 21330 13830 21400
rect 13850 21330 13920 21400
rect 13940 21330 14010 21400
rect 14030 21330 14100 21400
rect 14120 21330 14190 21400
rect 14210 21330 14280 21400
rect 14300 21330 14370 21400
rect 14390 21330 14460 21400
rect 14480 21330 14550 21400
rect 14570 21330 14640 21400
rect 14660 21330 14730 21400
rect 14750 21330 14820 21400
rect 14840 21330 14910 21400
rect 14930 21330 15000 21400
rect 15020 21330 15090 21400
rect 15110 21330 15180 21400
rect 15200 21330 15270 21400
rect 15290 21330 15360 21400
rect 15380 21330 15450 21400
rect 15470 21330 15540 21400
rect 15560 21330 15630 21400
rect 15650 21330 15720 21400
rect 15740 21330 15810 21400
rect 15830 21330 15900 21400
rect 15920 21330 15990 21400
rect 16010 21330 16080 21400
rect 16100 21330 16170 21400
rect 16190 21330 16260 21400
rect 16280 21330 16350 21400
rect 16370 21330 16440 21400
rect 16460 21330 16530 21400
rect 16550 21330 16620 21400
rect 16680 21330 16750 21400
rect 16770 21330 16840 21400
rect 16860 21330 16930 21400
rect 16950 21330 17020 21400
rect 17040 21330 17110 21400
rect 17130 21330 17200 21400
rect 17220 21330 17290 21400
rect 17310 21330 17380 21400
rect 17400 21330 17470 21400
rect 17490 21330 17560 21400
rect 17580 21330 17650 21400
rect 17670 21330 17740 21400
rect 17760 21330 17830 21400
rect 17850 21330 17920 21400
rect 17940 21330 18010 21400
rect 18030 21330 18100 21400
rect 18120 21330 18190 21400
rect 18210 21330 18280 21400
rect 18300 21330 18370 21400
rect 18390 21330 18460 21400
rect 18480 21330 18550 21400
rect 18570 21330 18640 21400
rect 18660 21330 18730 21400
rect 18750 21330 18820 21400
rect 18840 21330 18910 21400
rect 18930 21330 19000 21400
rect 19020 21330 19090 21400
rect 19110 21330 19180 21400
rect 19200 21330 19270 21400
rect 19290 21330 19360 21400
rect 19380 21330 19450 21400
rect 19470 21330 19540 21400
rect 19560 21330 19630 21400
rect 7040 8340 7140 8410
rect 7170 8340 7270 8410
rect 7040 8250 7140 8320
rect 7170 8250 7270 8320
rect 1570 6780 1640 6850
rect 1680 6780 1750 6850
rect 1790 6780 1860 6850
rect 1900 6780 1970 6850
rect 2010 6780 2080 6850
rect 2120 6780 2190 6850
rect 2230 6780 2300 6850
rect 2340 6780 2410 6850
rect 2450 6780 2520 6850
rect 2560 6780 2630 6850
rect 2670 6780 2740 6850
rect 2780 6780 2850 6850
rect 2890 6780 2960 6850
rect 3000 6780 3070 6850
rect 1570 6670 1640 6740
rect 1680 6670 1750 6740
rect 1790 6670 1860 6740
rect 1900 6670 1970 6740
rect 2010 6670 2080 6740
rect 2120 6670 2190 6740
rect 2230 6670 2300 6740
rect 2340 6670 2410 6740
rect 2450 6670 2520 6740
rect 2560 6670 2630 6740
rect 2670 6670 2740 6740
rect 2780 6670 2850 6740
rect 2890 6670 2960 6740
rect 3000 6670 3070 6740
rect 7630 8340 7730 8410
rect 7760 8340 7860 8410
rect 7630 8250 7730 8320
rect 7760 8250 7860 8320
rect 7410 5320 7480 5390
rect 7410 5210 7480 5280
rect 7410 5100 7480 5170
rect 7410 4990 7480 5060
rect 7410 4880 7480 4950
rect 38190 7750 38260 7820
rect 38280 7750 38350 7820
rect 38370 7750 38440 7820
rect 38190 7660 38260 7730
rect 38280 7660 38350 7730
rect 38370 7660 38440 7730
rect 38190 7570 38260 7640
rect 38280 7570 38350 7640
rect 38370 7570 38440 7640
rect 38190 7480 38260 7550
rect 38280 7480 38350 7550
rect 38370 7480 38440 7550
rect 38190 7390 38260 7460
rect 38280 7390 38350 7460
rect 38370 7390 38440 7460
rect 38190 7300 38260 7370
rect 38280 7300 38350 7370
rect 38370 7300 38440 7370
rect 23490 7140 23560 7210
rect 23600 7140 23670 7210
rect 23710 7140 23780 7210
rect 23820 7140 23890 7210
rect 23490 7030 23560 7100
rect 23600 7030 23670 7100
rect 23710 7030 23780 7100
rect 23820 7030 23890 7100
rect 25890 7140 25960 7210
rect 26000 7140 26070 7210
rect 26110 7140 26180 7210
rect 26220 7140 26290 7210
rect 25890 7030 25960 7100
rect 26000 7030 26070 7100
rect 26110 7030 26180 7100
rect 26220 7030 26290 7100
rect 38190 7210 38260 7280
rect 38280 7210 38350 7280
rect 38370 7210 38440 7280
rect 38190 7080 38260 7150
rect 38280 7080 38350 7150
rect 38370 7080 38440 7150
rect 38190 6990 38260 7060
rect 38280 6990 38350 7060
rect 38370 6990 38440 7060
rect 11790 6810 11860 6880
rect 11900 6810 11970 6880
rect 12010 6810 12080 6880
rect 12120 6810 12190 6880
rect 12230 6810 12300 6880
rect 12340 6810 12410 6880
rect 12450 6810 12520 6880
rect 12560 6810 12630 6880
rect 12670 6810 12740 6880
rect 12780 6810 12850 6880
rect 12890 6810 12960 6880
rect 13000 6810 13070 6880
rect 13110 6810 13180 6880
rect 13220 6810 13290 6880
rect 11790 6700 11860 6770
rect 11900 6700 11970 6770
rect 12010 6700 12080 6770
rect 12120 6700 12190 6770
rect 12230 6700 12300 6770
rect 12340 6700 12410 6770
rect 12450 6700 12520 6770
rect 12560 6700 12630 6770
rect 12670 6700 12740 6770
rect 12780 6700 12850 6770
rect 12890 6700 12960 6770
rect 13000 6700 13070 6770
rect 13110 6700 13180 6770
rect 13220 6700 13290 6770
rect 38190 6900 38260 6970
rect 38280 6900 38350 6970
rect 38370 6900 38440 6970
rect 38190 6810 38260 6880
rect 38280 6810 38350 6880
rect 38370 6810 38440 6880
rect 38190 6720 38260 6790
rect 38280 6720 38350 6790
rect 38370 6720 38440 6790
rect 38190 6630 38260 6700
rect 38280 6630 38350 6700
rect 38370 6630 38440 6700
rect 38190 6540 38260 6610
rect 38280 6540 38350 6610
rect 38370 6540 38440 6610
rect 38190 6450 38260 6520
rect 38280 6450 38350 6520
rect 38370 6450 38440 6520
rect 38190 6360 38260 6430
rect 38280 6360 38350 6430
rect 38370 6360 38440 6430
rect 30740 6230 30810 6300
rect 30850 6230 30920 6300
rect 30740 6100 30810 6170
rect 30850 6100 30920 6170
rect 30740 5970 30810 6040
rect 30850 5970 30920 6040
rect 38190 6270 38260 6340
rect 38280 6270 38350 6340
rect 38370 6270 38440 6340
rect 38190 6180 38260 6250
rect 38280 6180 38350 6250
rect 38370 6180 38440 6250
rect 38190 6090 38260 6160
rect 38280 6090 38350 6160
rect 38370 6090 38440 6160
rect 38190 6000 38260 6070
rect 38280 6000 38350 6070
rect 38370 6000 38440 6070
rect 38190 5910 38260 5980
rect 38280 5910 38350 5980
rect 38370 5910 38440 5980
rect 38190 5820 38260 5890
rect 38280 5820 38350 5890
rect 38370 5820 38440 5890
rect 38190 5730 38260 5800
rect 38280 5730 38350 5800
rect 38370 5730 38440 5800
rect 21820 5600 21890 5670
rect 21930 5600 22000 5670
rect 21820 5490 21890 5560
rect 21930 5490 22000 5560
rect 21820 5380 21890 5450
rect 21930 5380 22000 5450
rect 21820 5270 21890 5340
rect 21930 5270 22000 5340
rect 21820 5160 21890 5230
rect 21930 5160 22000 5230
rect 21820 5050 21890 5120
rect 21930 5050 22000 5120
rect 21820 4940 21890 5010
rect 21930 4940 22000 5010
rect 21820 4830 21890 4900
rect 21930 4830 22000 4900
rect 21820 4720 21890 4790
rect 21930 4720 22000 4790
rect 21820 4610 21890 4680
rect 21930 4610 22000 4680
rect 21820 4500 21890 4570
rect 21930 4500 22000 4570
rect 38190 5640 38260 5710
rect 38280 5640 38350 5710
rect 38370 5640 38440 5710
rect 38190 5550 38260 5620
rect 38280 5550 38350 5620
rect 38370 5550 38440 5620
rect 38190 5460 38260 5530
rect 38280 5460 38350 5530
rect 38370 5460 38440 5530
rect 38190 5370 38260 5440
rect 38280 5370 38350 5440
rect 38370 5370 38440 5440
rect 38190 5280 38260 5350
rect 38280 5280 38350 5350
rect 38370 5280 38440 5350
rect 38190 5190 38260 5260
rect 38280 5190 38350 5260
rect 38370 5190 38440 5260
rect 38190 5100 38260 5170
rect 38280 5100 38350 5170
rect 38370 5100 38440 5170
rect 38190 5010 38260 5080
rect 38280 5010 38350 5080
rect 38370 5010 38440 5080
rect 38190 4920 38260 4990
rect 38280 4920 38350 4990
rect 38370 4920 38440 4990
rect 38190 4830 38260 4900
rect 38280 4830 38350 4900
rect 38370 4830 38440 4900
rect 38190 4740 38260 4810
rect 38280 4740 38350 4810
rect 38370 4740 38440 4810
rect 38190 4650 38260 4720
rect 38280 4650 38350 4720
rect 38370 4650 38440 4720
rect 38190 4560 38260 4630
rect 38280 4560 38350 4630
rect 38370 4560 38440 4630
rect 38190 4470 38260 4540
rect 38280 4470 38350 4540
rect 38370 4470 38440 4540
rect 38190 4380 38260 4450
rect 38280 4380 38350 4450
rect 38370 4380 38440 4450
rect 38190 4290 38260 4360
rect 38280 4290 38350 4360
rect 38370 4290 38440 4360
rect 38190 4200 38260 4270
rect 38280 4200 38350 4270
rect 38370 4200 38440 4270
rect 38190 4070 38260 4140
rect 38280 4070 38350 4140
rect 38370 4070 38440 4140
rect 38190 3980 38260 4050
rect 38280 3980 38350 4050
rect 38370 3980 38440 4050
rect 38190 3890 38260 3960
rect 38280 3890 38350 3960
rect 38370 3890 38440 3960
rect 38190 3800 38260 3870
rect 38280 3800 38350 3870
rect 38370 3800 38440 3870
rect 38190 3710 38260 3780
rect 38280 3710 38350 3780
rect 38370 3710 38440 3780
rect 38190 3620 38260 3690
rect 38280 3620 38350 3690
rect 38370 3620 38440 3690
rect 38190 3530 38260 3600
rect 38280 3530 38350 3600
rect 38370 3530 38440 3600
rect 38190 3440 38260 3510
rect 38280 3440 38350 3510
rect 38370 3440 38440 3510
rect 24720 3290 24790 3360
rect 24830 3290 24900 3360
rect 24940 3290 25010 3360
rect 24720 3180 24790 3250
rect 24830 3180 24900 3250
rect 24940 3180 25010 3250
rect 24720 3070 24790 3140
rect 24830 3070 24900 3140
rect 24940 3070 25010 3140
rect 38190 3350 38260 3420
rect 38280 3350 38350 3420
rect 38370 3350 38440 3420
rect 38190 3260 38260 3330
rect 38280 3260 38350 3330
rect 38370 3260 38440 3330
rect 38190 3170 38260 3240
rect 38280 3170 38350 3240
rect 38370 3170 38440 3240
rect 38190 3080 38260 3150
rect 38280 3080 38350 3150
rect 38370 3080 38440 3150
rect 38190 2990 38260 3060
rect 38280 2990 38350 3060
rect 38370 2990 38440 3060
rect 1150 -860 1220 -790
rect 1260 -860 1330 -790
rect 1370 -860 1440 -790
rect 1480 -860 1550 -790
rect 1590 -860 1660 -790
rect 1700 -860 1770 -790
rect 1810 -860 1880 -790
rect 1920 -860 1990 -790
rect 2030 -860 2100 -790
rect 2140 -860 2210 -790
rect 2250 -860 2320 -790
rect 2360 -860 2430 -790
rect 2470 -860 2540 -790
rect 2580 -860 2650 -790
rect 1150 -970 1220 -900
rect 1260 -970 1330 -900
rect 1370 -970 1440 -900
rect 1480 -970 1550 -900
rect 1590 -970 1660 -900
rect 1700 -970 1770 -900
rect 1810 -970 1880 -900
rect 1920 -970 1990 -900
rect 2030 -970 2100 -900
rect 2140 -970 2210 -900
rect 2250 -970 2320 -900
rect 2360 -970 2430 -900
rect 2470 -970 2540 -900
rect 2580 -970 2650 -900
rect 1570 -2850 1640 -2780
rect 1680 -2850 1750 -2780
rect 1790 -2850 1860 -2780
rect 1900 -2850 1970 -2780
rect 2010 -2850 2080 -2780
rect 2120 -2850 2190 -2780
rect 2230 -2850 2300 -2780
rect 2340 -2850 2410 -2780
rect 2450 -2850 2520 -2780
rect 2560 -2850 2630 -2780
rect 2670 -2850 2740 -2780
rect 2780 -2850 2850 -2780
rect 2890 -2850 2960 -2780
rect 3000 -2850 3070 -2780
rect 1570 -2960 1640 -2890
rect 1680 -2960 1750 -2890
rect 1790 -2960 1860 -2890
rect 1900 -2960 1970 -2890
rect 2010 -2960 2080 -2890
rect 2120 -2960 2190 -2890
rect 2230 -2960 2300 -2890
rect 2340 -2960 2410 -2890
rect 2450 -2960 2520 -2890
rect 2560 -2960 2630 -2890
rect 2670 -2960 2740 -2890
rect 2780 -2960 2850 -2890
rect 2890 -2960 2960 -2890
rect 3000 -2960 3070 -2890
rect 38190 2900 38260 2970
rect 38280 2900 38350 2970
rect 38370 2900 38440 2970
rect 38190 2810 38260 2880
rect 38280 2810 38350 2880
rect 38370 2810 38440 2880
rect 38190 2720 38260 2790
rect 38280 2720 38350 2790
rect 38370 2720 38440 2790
rect 38190 2630 38260 2700
rect 38280 2630 38350 2700
rect 38370 2630 38440 2700
rect 22470 2530 22540 2600
rect 22580 2530 22650 2600
rect 22690 2530 22760 2600
rect 22800 2530 22870 2600
rect 22470 2420 22540 2490
rect 22580 2420 22650 2490
rect 22690 2420 22760 2490
rect 22800 2420 22870 2490
rect 26950 2530 27020 2600
rect 27060 2530 27130 2600
rect 27170 2530 27240 2600
rect 27280 2530 27350 2600
rect 26950 2420 27020 2490
rect 27060 2420 27130 2490
rect 27170 2420 27240 2490
rect 27280 2420 27350 2490
rect 38190 2540 38260 2610
rect 38280 2540 38350 2610
rect 38370 2540 38440 2610
rect 38190 2450 38260 2520
rect 38280 2450 38350 2520
rect 38370 2450 38440 2520
rect 38190 2360 38260 2430
rect 38280 2360 38350 2430
rect 38370 2360 38440 2430
rect 38190 2270 38260 2340
rect 38280 2270 38350 2340
rect 38370 2270 38440 2340
rect 38190 2180 38260 2250
rect 38280 2180 38350 2250
rect 38370 2180 38440 2250
rect 38190 2090 38260 2160
rect 38280 2090 38350 2160
rect 38370 2090 38440 2160
rect 38190 2000 38260 2070
rect 38280 2000 38350 2070
rect 38370 2000 38440 2070
rect 38190 1910 38260 1980
rect 38280 1910 38350 1980
rect 38370 1910 38440 1980
rect 38190 1820 38260 1890
rect 38280 1820 38350 1890
rect 38370 1820 38440 1890
rect 38190 1730 38260 1800
rect 38280 1730 38350 1800
rect 38370 1730 38440 1800
rect 38190 1640 38260 1710
rect 38280 1640 38350 1710
rect 38370 1640 38440 1710
rect 38190 1550 38260 1620
rect 38280 1550 38350 1620
rect 38370 1550 38440 1620
rect 38190 1460 38260 1530
rect 38280 1460 38350 1530
rect 38370 1460 38440 1530
rect 38190 1370 38260 1440
rect 38280 1370 38350 1440
rect 38370 1370 38440 1440
rect 38190 1280 38260 1350
rect 38280 1280 38350 1350
rect 38370 1280 38440 1350
rect 38190 1190 38260 1260
rect 38280 1190 38350 1260
rect 38370 1190 38440 1260
rect 17480 1090 17550 1160
rect 17480 980 17550 1050
rect 17480 870 17550 940
rect 23490 850 23560 920
rect 23600 850 23670 920
rect 23710 850 23780 920
rect 23820 850 23890 920
rect 23490 740 23560 810
rect 23600 740 23670 810
rect 23710 740 23780 810
rect 23820 740 23890 810
rect 25890 850 25960 920
rect 26000 850 26070 920
rect 26110 850 26180 920
rect 26220 850 26290 920
rect 25890 740 25960 810
rect 26000 740 26070 810
rect 26110 740 26180 810
rect 26220 740 26290 810
rect 38190 150 38260 220
rect 38280 150 38350 220
rect 38370 150 38440 220
rect 38190 60 38260 130
rect 38280 60 38350 130
rect 38370 60 38440 130
rect 30740 -70 30810 0
rect 30850 -70 30920 0
rect 30740 -200 30810 -130
rect 30850 -200 30920 -130
rect 30740 -330 30810 -260
rect 30850 -330 30920 -260
rect 38190 -30 38260 40
rect 38280 -30 38350 40
rect 38370 -30 38440 40
rect 38190 -120 38260 -50
rect 38280 -120 38350 -50
rect 38370 -120 38440 -50
rect 38190 -210 38260 -140
rect 38280 -210 38350 -140
rect 38370 -210 38440 -140
rect 38190 -300 38260 -230
rect 38280 -300 38350 -230
rect 38370 -300 38440 -230
rect 7310 -3950 7380 -3880
rect 7420 -3950 7490 -3880
rect 7530 -3950 7600 -3880
rect 7310 -4060 7380 -3990
rect 7420 -4060 7490 -3990
rect 7530 -4060 7600 -3990
rect 7310 -4170 7380 -4100
rect 7420 -4170 7490 -4100
rect 7530 -4170 7600 -4100
rect -1330 -4420 -1260 -4350
rect -1220 -4420 -1150 -4350
rect -1110 -4420 -1040 -4350
rect -1000 -4420 -930 -4350
rect -1330 -4530 -1260 -4460
rect -1220 -4530 -1150 -4460
rect -1110 -4530 -1040 -4460
rect -1000 -4530 -930 -4460
rect -1160 -6400 -1090 -6330
rect -1070 -6400 -1000 -6330
rect -980 -6400 -910 -6330
rect -890 -6400 -820 -6330
rect -800 -6400 -730 -6330
rect -710 -6400 -640 -6330
rect -620 -6400 -550 -6330
rect -530 -6400 -460 -6330
rect -440 -6400 -370 -6330
rect -350 -6400 -280 -6330
rect -260 -6400 -190 -6330
rect -170 -6400 -100 -6330
rect -80 -6400 -10 -6330
rect 10 -6400 80 -6330
rect -1160 -6490 -1090 -6420
rect -1070 -6490 -1000 -6420
rect -980 -6490 -910 -6420
rect -890 -6490 -820 -6420
rect -800 -6490 -730 -6420
rect -710 -6490 -640 -6420
rect -620 -6490 -550 -6420
rect -530 -6490 -460 -6420
rect -440 -6490 -370 -6420
rect -350 -6490 -280 -6420
rect -260 -6490 -190 -6420
rect -170 -6490 -100 -6420
rect -80 -6490 -10 -6420
rect 10 -6490 80 -6420
rect -1160 -6580 -1090 -6510
rect -1070 -6580 -1000 -6510
rect -980 -6580 -910 -6510
rect -890 -6580 -820 -6510
rect -800 -6580 -730 -6510
rect -710 -6580 -640 -6510
rect -620 -6580 -550 -6510
rect -530 -6580 -460 -6510
rect -440 -6580 -370 -6510
rect -350 -6580 -280 -6510
rect -260 -6580 -190 -6510
rect -170 -6580 -100 -6510
rect -80 -6580 -10 -6510
rect 10 -6580 80 -6510
rect 38190 -390 38260 -320
rect 38280 -390 38350 -320
rect 38370 -390 38440 -320
rect 38190 -520 38260 -450
rect 38280 -520 38350 -450
rect 38370 -520 38440 -450
rect 38190 -610 38260 -540
rect 38280 -610 38350 -540
rect 38370 -610 38440 -540
rect 38190 -700 38260 -630
rect 38280 -700 38350 -630
rect 38370 -700 38440 -630
rect 12250 -860 12320 -790
rect 12360 -860 12430 -790
rect 12470 -860 12540 -790
rect 12580 -860 12650 -790
rect 12690 -860 12760 -790
rect 12800 -860 12870 -790
rect 12910 -860 12980 -790
rect 13020 -860 13090 -790
rect 13130 -860 13200 -790
rect 13240 -860 13310 -790
rect 13350 -860 13420 -790
rect 13460 -860 13530 -790
rect 13570 -860 13640 -790
rect 13680 -860 13750 -790
rect 38190 -790 38260 -720
rect 38280 -790 38350 -720
rect 38370 -790 38440 -720
rect 12250 -970 12320 -900
rect 12360 -970 12430 -900
rect 12470 -970 12540 -900
rect 12580 -970 12650 -900
rect 12690 -970 12760 -900
rect 12800 -970 12870 -900
rect 12910 -970 12980 -900
rect 13020 -970 13090 -900
rect 13130 -970 13200 -900
rect 13240 -970 13310 -900
rect 13350 -970 13420 -900
rect 13460 -970 13530 -900
rect 13570 -970 13640 -900
rect 13680 -970 13750 -900
rect 21820 -920 21890 -850
rect 21930 -920 22000 -850
rect 21820 -1030 21890 -960
rect 21930 -1030 22000 -960
rect 21820 -1140 21890 -1070
rect 21930 -1140 22000 -1070
rect 21820 -1250 21890 -1180
rect 21930 -1250 22000 -1180
rect 21820 -1360 21890 -1290
rect 21930 -1360 22000 -1290
rect 21820 -1470 21890 -1400
rect 21930 -1470 22000 -1400
rect 21820 -1580 21890 -1510
rect 21930 -1580 22000 -1510
rect 21820 -1690 21890 -1620
rect 21930 -1690 22000 -1620
rect 21820 -1800 21890 -1730
rect 21930 -1800 22000 -1730
rect 21820 -1910 21890 -1840
rect 21930 -1910 22000 -1840
rect 21820 -2020 21890 -1950
rect 21930 -2020 22000 -1950
rect 38190 -880 38260 -810
rect 38280 -880 38350 -810
rect 38370 -880 38440 -810
rect 38190 -970 38260 -900
rect 38280 -970 38350 -900
rect 38370 -970 38440 -900
rect 38190 -1060 38260 -990
rect 38280 -1060 38350 -990
rect 38370 -1060 38440 -990
rect 38190 -1150 38260 -1080
rect 38280 -1150 38350 -1080
rect 38370 -1150 38440 -1080
rect 38190 -1240 38260 -1170
rect 38280 -1240 38350 -1170
rect 38370 -1240 38440 -1170
rect 38190 -1330 38260 -1260
rect 38280 -1330 38350 -1260
rect 38370 -1330 38440 -1260
rect 38190 -1420 38260 -1350
rect 38280 -1420 38350 -1350
rect 38370 -1420 38440 -1350
rect 38190 -1510 38260 -1440
rect 38280 -1510 38350 -1440
rect 38370 -1510 38440 -1440
rect 38190 -1600 38260 -1530
rect 38280 -1600 38350 -1530
rect 38370 -1600 38440 -1530
rect 38190 -1690 38260 -1620
rect 38280 -1690 38350 -1620
rect 38370 -1690 38440 -1620
rect 38190 -1780 38260 -1710
rect 38280 -1780 38350 -1710
rect 38370 -1780 38440 -1710
rect 38190 -1870 38260 -1800
rect 38280 -1870 38350 -1800
rect 38370 -1870 38440 -1800
rect 38190 -1960 38260 -1890
rect 38280 -1960 38350 -1890
rect 38370 -1960 38440 -1890
rect 38190 -2050 38260 -1980
rect 38280 -2050 38350 -1980
rect 38370 -2050 38440 -1980
rect 38190 -2140 38260 -2070
rect 38280 -2140 38350 -2070
rect 38370 -2140 38440 -2070
rect 38190 -2230 38260 -2160
rect 38280 -2230 38350 -2160
rect 38370 -2230 38440 -2160
rect 38190 -2320 38260 -2250
rect 38280 -2320 38350 -2250
rect 38370 -2320 38440 -2250
rect 38190 -2410 38260 -2340
rect 38280 -2410 38350 -2340
rect 38370 -2410 38440 -2340
rect 38190 -2500 38260 -2430
rect 38280 -2500 38350 -2430
rect 38370 -2500 38440 -2430
rect 38190 -2590 38260 -2520
rect 38280 -2590 38350 -2520
rect 38370 -2590 38440 -2520
rect 38190 -2680 38260 -2610
rect 38280 -2680 38350 -2610
rect 38370 -2680 38440 -2610
rect 11790 -2850 11860 -2780
rect 11900 -2850 11970 -2780
rect 12010 -2850 12080 -2780
rect 12120 -2850 12190 -2780
rect 12230 -2850 12300 -2780
rect 12340 -2850 12410 -2780
rect 12450 -2850 12520 -2780
rect 12560 -2850 12630 -2780
rect 12670 -2850 12740 -2780
rect 12780 -2850 12850 -2780
rect 12890 -2850 12960 -2780
rect 13000 -2850 13070 -2780
rect 13110 -2850 13180 -2780
rect 13220 -2850 13290 -2780
rect 11790 -2960 11860 -2890
rect 11900 -2960 11970 -2890
rect 12010 -2960 12080 -2890
rect 12120 -2960 12190 -2890
rect 12230 -2960 12300 -2890
rect 12340 -2960 12410 -2890
rect 12450 -2960 12520 -2890
rect 12560 -2960 12630 -2890
rect 12670 -2960 12740 -2890
rect 12780 -2960 12850 -2890
rect 12890 -2960 12960 -2890
rect 13000 -2960 13070 -2890
rect 13110 -2960 13180 -2890
rect 13220 -2960 13290 -2890
rect 38190 -2770 38260 -2700
rect 38280 -2770 38350 -2700
rect 38370 -2770 38440 -2700
rect 38190 -2860 38260 -2790
rect 38280 -2860 38350 -2790
rect 38370 -2860 38440 -2790
rect 38190 -2950 38260 -2880
rect 38280 -2950 38350 -2880
rect 38370 -2950 38440 -2880
rect 24740 -3120 24810 -3050
rect 24850 -3120 24920 -3050
rect 24960 -3120 25030 -3050
rect 24740 -3230 24810 -3160
rect 24850 -3230 24920 -3160
rect 24960 -3230 25030 -3160
rect 24740 -3340 24810 -3270
rect 24850 -3340 24920 -3270
rect 24960 -3340 25030 -3270
rect 38190 -3040 38260 -2970
rect 38280 -3040 38350 -2970
rect 38370 -3040 38440 -2970
rect 38190 -3130 38260 -3060
rect 38280 -3130 38350 -3060
rect 38370 -3130 38440 -3060
rect 38190 -3220 38260 -3150
rect 38280 -3220 38350 -3150
rect 38370 -3220 38440 -3150
rect 38190 -3310 38260 -3240
rect 38280 -3310 38350 -3240
rect 38370 -3310 38440 -3240
rect 38190 -3400 38260 -3330
rect 38280 -3400 38350 -3330
rect 38370 -3400 38440 -3330
rect 38190 -3530 38260 -3460
rect 38280 -3530 38350 -3460
rect 38370 -3530 38440 -3460
rect 38190 -3620 38260 -3550
rect 38280 -3620 38350 -3550
rect 38370 -3620 38440 -3550
rect 22470 -3760 22540 -3690
rect 22580 -3760 22650 -3690
rect 22690 -3760 22760 -3690
rect 22800 -3760 22870 -3690
rect 22470 -3870 22540 -3800
rect 22580 -3870 22650 -3800
rect 22690 -3870 22760 -3800
rect 22800 -3870 22870 -3800
rect 26950 -3760 27020 -3690
rect 27060 -3760 27130 -3690
rect 27170 -3760 27240 -3690
rect 27280 -3760 27350 -3690
rect 26950 -3870 27020 -3800
rect 27060 -3870 27130 -3800
rect 27170 -3870 27240 -3800
rect 27280 -3870 27350 -3800
rect 38190 -3710 38260 -3640
rect 38280 -3710 38350 -3640
rect 38370 -3710 38440 -3640
rect 38190 -3800 38260 -3730
rect 38280 -3800 38350 -3730
rect 38370 -3800 38440 -3730
rect 38190 -3890 38260 -3820
rect 38280 -3890 38350 -3820
rect 38370 -3890 38440 -3820
rect 38190 -3980 38260 -3910
rect 38280 -3980 38350 -3910
rect 38370 -3980 38440 -3910
rect 38190 -4070 38260 -4000
rect 38280 -4070 38350 -4000
rect 38370 -4070 38440 -4000
rect 38190 -4160 38260 -4090
rect 38280 -4160 38350 -4090
rect 38370 -4160 38440 -4090
rect 38190 -4250 38260 -4180
rect 38280 -4250 38350 -4180
rect 38370 -4250 38440 -4180
rect 15710 -4420 15780 -4350
rect 15820 -4420 15890 -4350
rect 15930 -4420 16000 -4350
rect 16040 -4420 16110 -4350
rect 15710 -4530 15780 -4460
rect 15820 -4530 15890 -4460
rect 15930 -4530 16000 -4460
rect 16040 -4530 16110 -4460
rect 38190 -4340 38260 -4270
rect 38280 -4340 38350 -4270
rect 38370 -4340 38440 -4270
rect 38190 -4430 38260 -4360
rect 38280 -4430 38350 -4360
rect 38370 -4430 38440 -4360
rect 38190 -4520 38260 -4450
rect 38280 -4520 38350 -4450
rect 38370 -4520 38440 -4450
rect 38190 -4610 38260 -4540
rect 38280 -4610 38350 -4540
rect 38370 -4610 38440 -4540
rect 14700 -6400 14770 -6330
rect 14790 -6400 14860 -6330
rect 14880 -6400 14950 -6330
rect 14970 -6400 15040 -6330
rect 15060 -6400 15130 -6330
rect 15150 -6400 15220 -6330
rect 15240 -6400 15310 -6330
rect 15330 -6400 15400 -6330
rect 15420 -6400 15490 -6330
rect 15510 -6400 15580 -6330
rect 15600 -6400 15670 -6330
rect 15690 -6400 15760 -6330
rect 15780 -6400 15850 -6330
rect 15870 -6400 15940 -6330
rect 14700 -6490 14770 -6420
rect 14790 -6490 14860 -6420
rect 14880 -6490 14950 -6420
rect 14970 -6490 15040 -6420
rect 15060 -6490 15130 -6420
rect 15150 -6490 15220 -6420
rect 15240 -6490 15310 -6420
rect 15330 -6490 15400 -6420
rect 15420 -6490 15490 -6420
rect 15510 -6490 15580 -6420
rect 15600 -6490 15670 -6420
rect 15690 -6490 15760 -6420
rect 15780 -6490 15850 -6420
rect 15870 -6490 15940 -6420
rect 38190 -4700 38260 -4630
rect 38280 -4700 38350 -4630
rect 38370 -4700 38440 -4630
rect 38190 -4790 38260 -4720
rect 38280 -4790 38350 -4720
rect 38370 -4790 38440 -4720
rect 38190 -4880 38260 -4810
rect 38280 -4880 38350 -4810
rect 38370 -4880 38440 -4810
rect 38190 -4970 38260 -4900
rect 38280 -4970 38350 -4900
rect 38370 -4970 38440 -4900
rect 38190 -5060 38260 -4990
rect 38280 -5060 38350 -4990
rect 38370 -5060 38440 -4990
rect 38190 -5150 38260 -5080
rect 38280 -5150 38350 -5080
rect 38370 -5150 38440 -5080
rect 38190 -5240 38260 -5170
rect 38280 -5240 38350 -5170
rect 38370 -5240 38440 -5170
rect 38190 -5330 38260 -5260
rect 38280 -5330 38350 -5260
rect 38370 -5330 38440 -5260
rect 38190 -5420 38260 -5350
rect 38280 -5420 38350 -5350
rect 38370 -5420 38440 -5350
rect 38190 -5510 38260 -5440
rect 38280 -5510 38350 -5440
rect 38370 -5510 38440 -5440
rect 38190 -5600 38260 -5530
rect 38280 -5600 38350 -5530
rect 38370 -5600 38440 -5530
rect 38190 -5690 38260 -5620
rect 38280 -5690 38350 -5620
rect 38370 -5690 38440 -5620
rect 38190 -5780 38260 -5710
rect 38280 -5780 38350 -5710
rect 38370 -5780 38440 -5710
rect 38190 -5870 38260 -5800
rect 38280 -5870 38350 -5800
rect 38370 -5870 38440 -5800
rect 38190 -5960 38260 -5890
rect 38280 -5960 38350 -5890
rect 38370 -5960 38440 -5890
rect 38190 -6050 38260 -5980
rect 38280 -6050 38350 -5980
rect 38370 -6050 38440 -5980
rect 38190 -6140 38260 -6070
rect 38280 -6140 38350 -6070
rect 38370 -6140 38440 -6070
rect 38190 -6230 38260 -6160
rect 38280 -6230 38350 -6160
rect 38370 -6230 38440 -6160
rect 38190 -6320 38260 -6250
rect 38280 -6320 38350 -6250
rect 38370 -6320 38440 -6250
rect 38190 -6410 38260 -6340
rect 38280 -6410 38350 -6340
rect 38370 -6410 38440 -6340
rect 14700 -6580 14770 -6510
rect 14790 -6580 14860 -6510
rect 14880 -6580 14950 -6510
rect 14970 -6580 15040 -6510
rect 15060 -6580 15130 -6510
rect 15150 -6580 15220 -6510
rect 15240 -6580 15310 -6510
rect 15330 -6580 15400 -6510
rect 15420 -6580 15490 -6510
rect 15510 -6580 15580 -6510
rect 15600 -6580 15670 -6510
rect 15690 -6580 15760 -6510
rect 15780 -6580 15850 -6510
rect 15870 -6580 15940 -6510
rect 1150 -10410 1220 -10340
rect 1260 -10410 1330 -10340
rect 1370 -10410 1440 -10340
rect 1480 -10410 1550 -10340
rect 1590 -10410 1660 -10340
rect 1700 -10410 1770 -10340
rect 1810 -10410 1880 -10340
rect 1920 -10410 1990 -10340
rect 2030 -10410 2100 -10340
rect 2140 -10410 2210 -10340
rect 2250 -10410 2320 -10340
rect 2360 -10410 2430 -10340
rect 2470 -10410 2540 -10340
rect 2580 -10410 2650 -10340
rect 1150 -10520 1220 -10450
rect 1260 -10520 1330 -10450
rect 1370 -10520 1440 -10450
rect 1480 -10520 1550 -10450
rect 1590 -10520 1660 -10450
rect 1700 -10520 1770 -10450
rect 1810 -10520 1880 -10450
rect 1920 -10520 1990 -10450
rect 2030 -10520 2100 -10450
rect 2140 -10520 2210 -10450
rect 2250 -10520 2320 -10450
rect 2360 -10520 2430 -10450
rect 2470 -10520 2540 -10450
rect 2580 -10520 2650 -10450
rect 2240 -12370 2310 -12300
rect 2350 -12370 2420 -12300
rect 2460 -12370 2530 -12300
rect 2570 -12370 2640 -12300
rect 2680 -12370 2750 -12300
rect 2790 -12370 2860 -12300
rect 2900 -12370 2970 -12300
rect 3010 -12370 3080 -12300
rect 3120 -12370 3190 -12300
rect 3230 -12370 3300 -12300
rect 3340 -12370 3410 -12300
rect 3450 -12370 3520 -12300
rect 3560 -12370 3630 -12300
rect 3670 -12370 3740 -12300
rect 2240 -12480 2310 -12410
rect 2350 -12480 2420 -12410
rect 2460 -12480 2530 -12410
rect 2570 -12480 2640 -12410
rect 2680 -12480 2750 -12410
rect 2790 -12480 2860 -12410
rect 2900 -12480 2970 -12410
rect 3010 -12480 3080 -12410
rect 3120 -12480 3190 -12410
rect 3230 -12480 3300 -12410
rect 3340 -12480 3410 -12410
rect 3450 -12480 3520 -12410
rect 3560 -12480 3630 -12410
rect 3670 -12480 3740 -12410
rect 14600 -8300 14670 -8230
rect 14700 -8300 14770 -8230
rect 14810 -8300 14880 -8230
rect 14600 -8410 14670 -8340
rect 14700 -8410 14770 -8340
rect 14810 -8410 14880 -8340
rect 14600 -8520 14670 -8450
rect 14700 -8520 14770 -8450
rect 14810 -8520 14880 -8450
rect 21630 -8430 21700 -8360
rect 21730 -8430 21800 -8360
rect 21830 -8430 21900 -8360
rect 21630 -8530 21700 -8460
rect 21730 -8530 21800 -8460
rect 21830 -8530 21900 -8460
rect 21630 -8630 21700 -8560
rect 21730 -8630 21800 -8560
rect 21830 -8630 21900 -8560
rect 22650 -9080 22720 -9010
rect 22750 -9080 22820 -9010
rect 22850 -9080 22920 -9010
rect 22650 -9180 22720 -9110
rect 22750 -9180 22820 -9110
rect 22850 -9180 22920 -9110
rect 22650 -9280 22720 -9210
rect 22750 -9280 22820 -9210
rect 22850 -9280 22920 -9210
rect 12290 -10440 12360 -10370
rect 12400 -10440 12470 -10370
rect 12510 -10440 12580 -10370
rect 12620 -10440 12690 -10370
rect 12730 -10440 12800 -10370
rect 12840 -10440 12910 -10370
rect 12950 -10440 13020 -10370
rect 13060 -10440 13130 -10370
rect 13170 -10440 13240 -10370
rect 13280 -10440 13350 -10370
rect 13390 -10440 13460 -10370
rect 13500 -10440 13570 -10370
rect 13610 -10440 13680 -10370
rect 13720 -10440 13790 -10370
rect 12290 -10550 12360 -10480
rect 12400 -10550 12470 -10480
rect 12510 -10550 12580 -10480
rect 12620 -10550 12690 -10480
rect 12730 -10550 12800 -10480
rect 12840 -10550 12910 -10480
rect 12950 -10550 13020 -10480
rect 13060 -10550 13130 -10480
rect 13170 -10550 13240 -10480
rect 13280 -10550 13350 -10480
rect 13390 -10550 13460 -10480
rect 13500 -10550 13570 -10480
rect 13610 -10550 13680 -10480
rect 13720 -10550 13790 -10480
rect 29990 -10590 30060 -10520
rect 30700 -10590 30770 -10520
rect 29990 -10700 30060 -10630
rect 30700 -10700 30770 -10630
rect 29990 -10810 30060 -10740
rect 30700 -10810 30770 -10740
rect 11120 -12370 11190 -12300
rect 11230 -12370 11300 -12300
rect 11340 -12370 11410 -12300
rect 11450 -12370 11520 -12300
rect 11560 -12370 11630 -12300
rect 11670 -12370 11740 -12300
rect 11780 -12370 11850 -12300
rect 11890 -12370 11960 -12300
rect 12000 -12370 12070 -12300
rect 12110 -12370 12180 -12300
rect 12220 -12370 12290 -12300
rect 12330 -12370 12400 -12300
rect 12440 -12370 12510 -12300
rect 12550 -12370 12620 -12300
rect 11120 -12480 11190 -12410
rect 11230 -12480 11300 -12410
rect 11340 -12480 11410 -12410
rect 11450 -12480 11520 -12410
rect 11560 -12480 11630 -12410
rect 11670 -12480 11740 -12410
rect 11780 -12480 11850 -12410
rect 11890 -12480 11960 -12410
rect 12000 -12480 12070 -12410
rect 12110 -12480 12180 -12410
rect 12220 -12480 12290 -12410
rect 12330 -12480 12400 -12410
rect 12440 -12480 12510 -12410
rect 12550 -12480 12620 -12410
rect 21630 -14090 21700 -14020
rect 21730 -14090 21800 -14020
rect 21830 -14090 21900 -14020
rect 21630 -14190 21700 -14120
rect 21730 -14190 21800 -14120
rect 21830 -14190 21900 -14120
rect 21630 -14290 21700 -14220
rect 21730 -14290 21800 -14220
rect 21830 -14290 21900 -14220
rect 22920 -14940 22990 -14870
rect 23020 -14940 23090 -14870
rect 23120 -14940 23190 -14870
rect 22920 -15040 22990 -14970
rect 23020 -15040 23090 -14970
rect 23120 -15040 23190 -14970
rect 22920 -15140 22990 -15070
rect 23020 -15140 23090 -15070
rect 23120 -15140 23190 -15070
rect 2280 -22730 2350 -22660
rect 2390 -22730 2460 -22660
rect 2500 -22730 2570 -22660
rect 2610 -22730 2680 -22660
rect 2720 -22730 2790 -22660
rect 2830 -22730 2900 -22660
rect 2940 -22730 3010 -22660
rect 3050 -22730 3120 -22660
rect 3160 -22730 3230 -22660
rect 3270 -22730 3340 -22660
rect 3380 -22730 3450 -22660
rect 3490 -22730 3560 -22660
rect 3600 -22730 3670 -22660
rect 3710 -22730 3780 -22660
rect 2280 -22840 2350 -22770
rect 2390 -22840 2460 -22770
rect 2500 -22840 2570 -22770
rect 2610 -22840 2680 -22770
rect 2720 -22840 2790 -22770
rect 2830 -22840 2900 -22770
rect 2940 -22840 3010 -22770
rect 3050 -22840 3120 -22770
rect 3160 -22840 3230 -22770
rect 3270 -22840 3340 -22770
rect 3380 -22840 3450 -22770
rect 3490 -22840 3560 -22770
rect 3600 -22840 3670 -22770
rect 3710 -22840 3780 -22770
rect 7230 -17670 7300 -17600
rect 7340 -17670 7410 -17600
rect 7450 -17670 7520 -17600
rect 7560 -17670 7630 -17600
rect 7230 -17780 7300 -17710
rect 7340 -17780 7410 -17710
rect 7450 -17780 7520 -17710
rect 7560 -17780 7630 -17710
rect 7230 -17890 7300 -17820
rect 7340 -17890 7410 -17820
rect 7450 -17890 7520 -17820
rect 7560 -17890 7630 -17820
rect 7230 -18000 7300 -17930
rect 7340 -18000 7410 -17930
rect 7450 -18000 7520 -17930
rect 7560 -18000 7630 -17930
rect 21630 -20170 21700 -20100
rect 21730 -20170 21800 -20100
rect 21830 -20170 21900 -20100
rect 21630 -20270 21700 -20200
rect 21730 -20270 21800 -20200
rect 21830 -20270 21900 -20200
rect 21630 -20370 21700 -20300
rect 21730 -20370 21800 -20300
rect 21830 -20370 21900 -20300
rect 22700 -20800 22770 -20730
rect 22800 -20800 22870 -20730
rect 22900 -20800 22970 -20730
rect 22700 -20900 22770 -20830
rect 22800 -20900 22870 -20830
rect 22900 -20900 22970 -20830
rect 22700 -21000 22770 -20930
rect 22800 -21000 22870 -20930
rect 22900 -21000 22970 -20930
rect 11160 -22730 11230 -22660
rect 11270 -22730 11340 -22660
rect 11380 -22730 11450 -22660
rect 11490 -22730 11560 -22660
rect 11600 -22730 11670 -22660
rect 11710 -22730 11780 -22660
rect 11820 -22730 11890 -22660
rect 11930 -22730 12000 -22660
rect 12040 -22730 12110 -22660
rect 12150 -22730 12220 -22660
rect 12260 -22730 12330 -22660
rect 12370 -22730 12440 -22660
rect 12480 -22730 12550 -22660
rect 12590 -22730 12660 -22660
rect 11160 -22840 11230 -22770
rect 11270 -22840 11340 -22770
rect 11380 -22840 11450 -22770
rect 11490 -22840 11560 -22770
rect 11600 -22840 11670 -22770
rect 11710 -22840 11780 -22770
rect 11820 -22840 11890 -22770
rect 11930 -22840 12000 -22770
rect 12040 -22840 12110 -22770
rect 12150 -22840 12220 -22770
rect 12260 -22840 12330 -22770
rect 12370 -22840 12440 -22770
rect 12480 -22840 12550 -22770
rect 12590 -22840 12660 -22770
<< mimcap >>
rect -4980 20830 7260 20960
rect -4980 20590 -4670 20830
rect -4430 20590 -4340 20830
rect -4100 20590 -4010 20830
rect -3770 20590 -3680 20830
rect -3440 20590 -3350 20830
rect -3110 20590 -3020 20830
rect -2780 20590 -2690 20830
rect -2450 20590 -2360 20830
rect -2120 20590 -2030 20830
rect -1790 20590 -1700 20830
rect -1460 20590 -1370 20830
rect -1130 20590 -1040 20830
rect -800 20590 -710 20830
rect -470 20590 -380 20830
rect -140 20590 -50 20830
rect 190 20590 280 20830
rect 520 20590 610 20830
rect 850 20590 940 20830
rect 1180 20590 1270 20830
rect 1510 20590 1600 20830
rect 1840 20590 1930 20830
rect 2170 20590 2260 20830
rect 2500 20590 2590 20830
rect 2830 20590 2920 20830
rect 3160 20590 3250 20830
rect 3490 20590 3580 20830
rect 3820 20590 3910 20830
rect 4150 20590 4240 20830
rect 4480 20590 4570 20830
rect 4810 20590 4900 20830
rect 5140 20590 5230 20830
rect 5470 20590 5560 20830
rect 5800 20590 5890 20830
rect 6130 20590 6220 20830
rect 6460 20590 6550 20830
rect 6790 20590 6880 20830
rect 7120 20590 7260 20830
rect -4980 20500 7260 20590
rect -4980 20260 -4670 20500
rect -4430 20260 -4340 20500
rect -4100 20260 -4010 20500
rect -3770 20260 -3680 20500
rect -3440 20260 -3350 20500
rect -3110 20260 -3020 20500
rect -2780 20260 -2690 20500
rect -2450 20260 -2360 20500
rect -2120 20260 -2030 20500
rect -1790 20260 -1700 20500
rect -1460 20260 -1370 20500
rect -1130 20260 -1040 20500
rect -800 20260 -710 20500
rect -470 20260 -380 20500
rect -140 20260 -50 20500
rect 190 20260 280 20500
rect 520 20260 610 20500
rect 850 20260 940 20500
rect 1180 20260 1270 20500
rect 1510 20260 1600 20500
rect 1840 20260 1930 20500
rect 2170 20260 2260 20500
rect 2500 20260 2590 20500
rect 2830 20260 2920 20500
rect 3160 20260 3250 20500
rect 3490 20260 3580 20500
rect 3820 20260 3910 20500
rect 4150 20260 4240 20500
rect 4480 20260 4570 20500
rect 4810 20260 4900 20500
rect 5140 20260 5230 20500
rect 5470 20260 5560 20500
rect 5800 20260 5890 20500
rect 6130 20260 6220 20500
rect 6460 20260 6550 20500
rect 6790 20260 6880 20500
rect 7120 20260 7260 20500
rect -4980 20170 7260 20260
rect -4980 19930 -4670 20170
rect -4430 19930 -4340 20170
rect -4100 19930 -4010 20170
rect -3770 19930 -3680 20170
rect -3440 19930 -3350 20170
rect -3110 19930 -3020 20170
rect -2780 19930 -2690 20170
rect -2450 19930 -2360 20170
rect -2120 19930 -2030 20170
rect -1790 19930 -1700 20170
rect -1460 19930 -1370 20170
rect -1130 19930 -1040 20170
rect -800 19930 -710 20170
rect -470 19930 -380 20170
rect -140 19930 -50 20170
rect 190 19930 280 20170
rect 520 19930 610 20170
rect 850 19930 940 20170
rect 1180 19930 1270 20170
rect 1510 19930 1600 20170
rect 1840 19930 1930 20170
rect 2170 19930 2260 20170
rect 2500 19930 2590 20170
rect 2830 19930 2920 20170
rect 3160 19930 3250 20170
rect 3490 19930 3580 20170
rect 3820 19930 3910 20170
rect 4150 19930 4240 20170
rect 4480 19930 4570 20170
rect 4810 19930 4900 20170
rect 5140 19930 5230 20170
rect 5470 19930 5560 20170
rect 5800 19930 5890 20170
rect 6130 19930 6220 20170
rect 6460 19930 6550 20170
rect 6790 19930 6880 20170
rect 7120 19930 7260 20170
rect -4980 19840 7260 19930
rect -4980 19600 -4670 19840
rect -4430 19600 -4340 19840
rect -4100 19600 -4010 19840
rect -3770 19600 -3680 19840
rect -3440 19600 -3350 19840
rect -3110 19600 -3020 19840
rect -2780 19600 -2690 19840
rect -2450 19600 -2360 19840
rect -2120 19600 -2030 19840
rect -1790 19600 -1700 19840
rect -1460 19600 -1370 19840
rect -1130 19600 -1040 19840
rect -800 19600 -710 19840
rect -470 19600 -380 19840
rect -140 19600 -50 19840
rect 190 19600 280 19840
rect 520 19600 610 19840
rect 850 19600 940 19840
rect 1180 19600 1270 19840
rect 1510 19600 1600 19840
rect 1840 19600 1930 19840
rect 2170 19600 2260 19840
rect 2500 19600 2590 19840
rect 2830 19600 2920 19840
rect 3160 19600 3250 19840
rect 3490 19600 3580 19840
rect 3820 19600 3910 19840
rect 4150 19600 4240 19840
rect 4480 19600 4570 19840
rect 4810 19600 4900 19840
rect 5140 19600 5230 19840
rect 5470 19600 5560 19840
rect 5800 19600 5890 19840
rect 6130 19600 6220 19840
rect 6460 19600 6550 19840
rect 6790 19600 6880 19840
rect 7120 19600 7260 19840
rect -4980 19510 7260 19600
rect -4980 19270 -4670 19510
rect -4430 19270 -4340 19510
rect -4100 19270 -4010 19510
rect -3770 19270 -3680 19510
rect -3440 19270 -3350 19510
rect -3110 19270 -3020 19510
rect -2780 19270 -2690 19510
rect -2450 19270 -2360 19510
rect -2120 19270 -2030 19510
rect -1790 19270 -1700 19510
rect -1460 19270 -1370 19510
rect -1130 19270 -1040 19510
rect -800 19270 -710 19510
rect -470 19270 -380 19510
rect -140 19270 -50 19510
rect 190 19270 280 19510
rect 520 19270 610 19510
rect 850 19270 940 19510
rect 1180 19270 1270 19510
rect 1510 19270 1600 19510
rect 1840 19270 1930 19510
rect 2170 19270 2260 19510
rect 2500 19270 2590 19510
rect 2830 19270 2920 19510
rect 3160 19270 3250 19510
rect 3490 19270 3580 19510
rect 3820 19270 3910 19510
rect 4150 19270 4240 19510
rect 4480 19270 4570 19510
rect 4810 19270 4900 19510
rect 5140 19270 5230 19510
rect 5470 19270 5560 19510
rect 5800 19270 5890 19510
rect 6130 19270 6220 19510
rect 6460 19270 6550 19510
rect 6790 19270 6880 19510
rect 7120 19270 7260 19510
rect -4980 19180 7260 19270
rect -4980 18940 -4670 19180
rect -4430 18940 -4340 19180
rect -4100 18940 -4010 19180
rect -3770 18940 -3680 19180
rect -3440 18940 -3350 19180
rect -3110 18940 -3020 19180
rect -2780 18940 -2690 19180
rect -2450 18940 -2360 19180
rect -2120 18940 -2030 19180
rect -1790 18940 -1700 19180
rect -1460 18940 -1370 19180
rect -1130 18940 -1040 19180
rect -800 18940 -710 19180
rect -470 18940 -380 19180
rect -140 18940 -50 19180
rect 190 18940 280 19180
rect 520 18940 610 19180
rect 850 18940 940 19180
rect 1180 18940 1270 19180
rect 1510 18940 1600 19180
rect 1840 18940 1930 19180
rect 2170 18940 2260 19180
rect 2500 18940 2590 19180
rect 2830 18940 2920 19180
rect 3160 18940 3250 19180
rect 3490 18940 3580 19180
rect 3820 18940 3910 19180
rect 4150 18940 4240 19180
rect 4480 18940 4570 19180
rect 4810 18940 4900 19180
rect 5140 18940 5230 19180
rect 5470 18940 5560 19180
rect 5800 18940 5890 19180
rect 6130 18940 6220 19180
rect 6460 18940 6550 19180
rect 6790 18940 6880 19180
rect 7120 18940 7260 19180
rect -4980 18850 7260 18940
rect -4980 18610 -4670 18850
rect -4430 18610 -4340 18850
rect -4100 18610 -4010 18850
rect -3770 18610 -3680 18850
rect -3440 18610 -3350 18850
rect -3110 18610 -3020 18850
rect -2780 18610 -2690 18850
rect -2450 18610 -2360 18850
rect -2120 18610 -2030 18850
rect -1790 18610 -1700 18850
rect -1460 18610 -1370 18850
rect -1130 18610 -1040 18850
rect -800 18610 -710 18850
rect -470 18610 -380 18850
rect -140 18610 -50 18850
rect 190 18610 280 18850
rect 520 18610 610 18850
rect 850 18610 940 18850
rect 1180 18610 1270 18850
rect 1510 18610 1600 18850
rect 1840 18610 1930 18850
rect 2170 18610 2260 18850
rect 2500 18610 2590 18850
rect 2830 18610 2920 18850
rect 3160 18610 3250 18850
rect 3490 18610 3580 18850
rect 3820 18610 3910 18850
rect 4150 18610 4240 18850
rect 4480 18610 4570 18850
rect 4810 18610 4900 18850
rect 5140 18610 5230 18850
rect 5470 18610 5560 18850
rect 5800 18610 5890 18850
rect 6130 18610 6220 18850
rect 6460 18610 6550 18850
rect 6790 18610 6880 18850
rect 7120 18610 7260 18850
rect -4980 18520 7260 18610
rect -4980 18280 -4670 18520
rect -4430 18280 -4340 18520
rect -4100 18280 -4010 18520
rect -3770 18280 -3680 18520
rect -3440 18280 -3350 18520
rect -3110 18280 -3020 18520
rect -2780 18280 -2690 18520
rect -2450 18280 -2360 18520
rect -2120 18280 -2030 18520
rect -1790 18280 -1700 18520
rect -1460 18280 -1370 18520
rect -1130 18280 -1040 18520
rect -800 18280 -710 18520
rect -470 18280 -380 18520
rect -140 18280 -50 18520
rect 190 18280 280 18520
rect 520 18280 610 18520
rect 850 18280 940 18520
rect 1180 18280 1270 18520
rect 1510 18280 1600 18520
rect 1840 18280 1930 18520
rect 2170 18280 2260 18520
rect 2500 18280 2590 18520
rect 2830 18280 2920 18520
rect 3160 18280 3250 18520
rect 3490 18280 3580 18520
rect 3820 18280 3910 18520
rect 4150 18280 4240 18520
rect 4480 18280 4570 18520
rect 4810 18280 4900 18520
rect 5140 18280 5230 18520
rect 5470 18280 5560 18520
rect 5800 18280 5890 18520
rect 6130 18280 6220 18520
rect 6460 18280 6550 18520
rect 6790 18280 6880 18520
rect 7120 18280 7260 18520
rect -4980 18190 7260 18280
rect -4980 17950 -4670 18190
rect -4430 17950 -4340 18190
rect -4100 17950 -4010 18190
rect -3770 17950 -3680 18190
rect -3440 17950 -3350 18190
rect -3110 17950 -3020 18190
rect -2780 17950 -2690 18190
rect -2450 17950 -2360 18190
rect -2120 17950 -2030 18190
rect -1790 17950 -1700 18190
rect -1460 17950 -1370 18190
rect -1130 17950 -1040 18190
rect -800 17950 -710 18190
rect -470 17950 -380 18190
rect -140 17950 -50 18190
rect 190 17950 280 18190
rect 520 17950 610 18190
rect 850 17950 940 18190
rect 1180 17950 1270 18190
rect 1510 17950 1600 18190
rect 1840 17950 1930 18190
rect 2170 17950 2260 18190
rect 2500 17950 2590 18190
rect 2830 17950 2920 18190
rect 3160 17950 3250 18190
rect 3490 17950 3580 18190
rect 3820 17950 3910 18190
rect 4150 17950 4240 18190
rect 4480 17950 4570 18190
rect 4810 17950 4900 18190
rect 5140 17950 5230 18190
rect 5470 17950 5560 18190
rect 5800 17950 5890 18190
rect 6130 17950 6220 18190
rect 6460 17950 6550 18190
rect 6790 17950 6880 18190
rect 7120 17950 7260 18190
rect -4980 17860 7260 17950
rect -4980 17620 -4670 17860
rect -4430 17620 -4340 17860
rect -4100 17620 -4010 17860
rect -3770 17620 -3680 17860
rect -3440 17620 -3350 17860
rect -3110 17620 -3020 17860
rect -2780 17620 -2690 17860
rect -2450 17620 -2360 17860
rect -2120 17620 -2030 17860
rect -1790 17620 -1700 17860
rect -1460 17620 -1370 17860
rect -1130 17620 -1040 17860
rect -800 17620 -710 17860
rect -470 17620 -380 17860
rect -140 17620 -50 17860
rect 190 17620 280 17860
rect 520 17620 610 17860
rect 850 17620 940 17860
rect 1180 17620 1270 17860
rect 1510 17620 1600 17860
rect 1840 17620 1930 17860
rect 2170 17620 2260 17860
rect 2500 17620 2590 17860
rect 2830 17620 2920 17860
rect 3160 17620 3250 17860
rect 3490 17620 3580 17860
rect 3820 17620 3910 17860
rect 4150 17620 4240 17860
rect 4480 17620 4570 17860
rect 4810 17620 4900 17860
rect 5140 17620 5230 17860
rect 5470 17620 5560 17860
rect 5800 17620 5890 17860
rect 6130 17620 6220 17860
rect 6460 17620 6550 17860
rect 6790 17620 6880 17860
rect 7120 17620 7260 17860
rect -4980 17530 7260 17620
rect -4980 17290 -4670 17530
rect -4430 17290 -4340 17530
rect -4100 17290 -4010 17530
rect -3770 17290 -3680 17530
rect -3440 17290 -3350 17530
rect -3110 17290 -3020 17530
rect -2780 17290 -2690 17530
rect -2450 17290 -2360 17530
rect -2120 17290 -2030 17530
rect -1790 17290 -1700 17530
rect -1460 17290 -1370 17530
rect -1130 17290 -1040 17530
rect -800 17290 -710 17530
rect -470 17290 -380 17530
rect -140 17290 -50 17530
rect 190 17290 280 17530
rect 520 17290 610 17530
rect 850 17290 940 17530
rect 1180 17290 1270 17530
rect 1510 17290 1600 17530
rect 1840 17290 1930 17530
rect 2170 17290 2260 17530
rect 2500 17290 2590 17530
rect 2830 17290 2920 17530
rect 3160 17290 3250 17530
rect 3490 17290 3580 17530
rect 3820 17290 3910 17530
rect 4150 17290 4240 17530
rect 4480 17290 4570 17530
rect 4810 17290 4900 17530
rect 5140 17290 5230 17530
rect 5470 17290 5560 17530
rect 5800 17290 5890 17530
rect 6130 17290 6220 17530
rect 6460 17290 6550 17530
rect 6790 17290 6880 17530
rect 7120 17290 7260 17530
rect -4980 17200 7260 17290
rect -4980 16960 -4670 17200
rect -4430 16960 -4340 17200
rect -4100 16960 -4010 17200
rect -3770 16960 -3680 17200
rect -3440 16960 -3350 17200
rect -3110 16960 -3020 17200
rect -2780 16960 -2690 17200
rect -2450 16960 -2360 17200
rect -2120 16960 -2030 17200
rect -1790 16960 -1700 17200
rect -1460 16960 -1370 17200
rect -1130 16960 -1040 17200
rect -800 16960 -710 17200
rect -470 16960 -380 17200
rect -140 16960 -50 17200
rect 190 16960 280 17200
rect 520 16960 610 17200
rect 850 16960 940 17200
rect 1180 16960 1270 17200
rect 1510 16960 1600 17200
rect 1840 16960 1930 17200
rect 2170 16960 2260 17200
rect 2500 16960 2590 17200
rect 2830 16960 2920 17200
rect 3160 16960 3250 17200
rect 3490 16960 3580 17200
rect 3820 16960 3910 17200
rect 4150 16960 4240 17200
rect 4480 16960 4570 17200
rect 4810 16960 4900 17200
rect 5140 16960 5230 17200
rect 5470 16960 5560 17200
rect 5800 16960 5890 17200
rect 6130 16960 6220 17200
rect 6460 16960 6550 17200
rect 6790 16960 6880 17200
rect 7120 16960 7260 17200
rect -4980 16870 7260 16960
rect -4980 16630 -4670 16870
rect -4430 16630 -4340 16870
rect -4100 16630 -4010 16870
rect -3770 16630 -3680 16870
rect -3440 16630 -3350 16870
rect -3110 16630 -3020 16870
rect -2780 16630 -2690 16870
rect -2450 16630 -2360 16870
rect -2120 16630 -2030 16870
rect -1790 16630 -1700 16870
rect -1460 16630 -1370 16870
rect -1130 16630 -1040 16870
rect -800 16630 -710 16870
rect -470 16630 -380 16870
rect -140 16630 -50 16870
rect 190 16630 280 16870
rect 520 16630 610 16870
rect 850 16630 940 16870
rect 1180 16630 1270 16870
rect 1510 16630 1600 16870
rect 1840 16630 1930 16870
rect 2170 16630 2260 16870
rect 2500 16630 2590 16870
rect 2830 16630 2920 16870
rect 3160 16630 3250 16870
rect 3490 16630 3580 16870
rect 3820 16630 3910 16870
rect 4150 16630 4240 16870
rect 4480 16630 4570 16870
rect 4810 16630 4900 16870
rect 5140 16630 5230 16870
rect 5470 16630 5560 16870
rect 5800 16630 5890 16870
rect 6130 16630 6220 16870
rect 6460 16630 6550 16870
rect 6790 16630 6880 16870
rect 7120 16630 7260 16870
rect -4980 16540 7260 16630
rect -4980 16300 -4670 16540
rect -4430 16300 -4340 16540
rect -4100 16300 -4010 16540
rect -3770 16300 -3680 16540
rect -3440 16300 -3350 16540
rect -3110 16300 -3020 16540
rect -2780 16300 -2690 16540
rect -2450 16300 -2360 16540
rect -2120 16300 -2030 16540
rect -1790 16300 -1700 16540
rect -1460 16300 -1370 16540
rect -1130 16300 -1040 16540
rect -800 16300 -710 16540
rect -470 16300 -380 16540
rect -140 16300 -50 16540
rect 190 16300 280 16540
rect 520 16300 610 16540
rect 850 16300 940 16540
rect 1180 16300 1270 16540
rect 1510 16300 1600 16540
rect 1840 16300 1930 16540
rect 2170 16300 2260 16540
rect 2500 16300 2590 16540
rect 2830 16300 2920 16540
rect 3160 16300 3250 16540
rect 3490 16300 3580 16540
rect 3820 16300 3910 16540
rect 4150 16300 4240 16540
rect 4480 16300 4570 16540
rect 4810 16300 4900 16540
rect 5140 16300 5230 16540
rect 5470 16300 5560 16540
rect 5800 16300 5890 16540
rect 6130 16300 6220 16540
rect 6460 16300 6550 16540
rect 6790 16300 6880 16540
rect 7120 16300 7260 16540
rect -4980 16210 7260 16300
rect -4980 15970 -4670 16210
rect -4430 15970 -4340 16210
rect -4100 15970 -4010 16210
rect -3770 15970 -3680 16210
rect -3440 15970 -3350 16210
rect -3110 15970 -3020 16210
rect -2780 15970 -2690 16210
rect -2450 15970 -2360 16210
rect -2120 15970 -2030 16210
rect -1790 15970 -1700 16210
rect -1460 15970 -1370 16210
rect -1130 15970 -1040 16210
rect -800 15970 -710 16210
rect -470 15970 -380 16210
rect -140 15970 -50 16210
rect 190 15970 280 16210
rect 520 15970 610 16210
rect 850 15970 940 16210
rect 1180 15970 1270 16210
rect 1510 15970 1600 16210
rect 1840 15970 1930 16210
rect 2170 15970 2260 16210
rect 2500 15970 2590 16210
rect 2830 15970 2920 16210
rect 3160 15970 3250 16210
rect 3490 15970 3580 16210
rect 3820 15970 3910 16210
rect 4150 15970 4240 16210
rect 4480 15970 4570 16210
rect 4810 15970 4900 16210
rect 5140 15970 5230 16210
rect 5470 15970 5560 16210
rect 5800 15970 5890 16210
rect 6130 15970 6220 16210
rect 6460 15970 6550 16210
rect 6790 15970 6880 16210
rect 7120 15970 7260 16210
rect -4980 15880 7260 15970
rect -4980 15640 -4670 15880
rect -4430 15640 -4340 15880
rect -4100 15640 -4010 15880
rect -3770 15640 -3680 15880
rect -3440 15640 -3350 15880
rect -3110 15640 -3020 15880
rect -2780 15640 -2690 15880
rect -2450 15640 -2360 15880
rect -2120 15640 -2030 15880
rect -1790 15640 -1700 15880
rect -1460 15640 -1370 15880
rect -1130 15640 -1040 15880
rect -800 15640 -710 15880
rect -470 15640 -380 15880
rect -140 15640 -50 15880
rect 190 15640 280 15880
rect 520 15640 610 15880
rect 850 15640 940 15880
rect 1180 15640 1270 15880
rect 1510 15640 1600 15880
rect 1840 15640 1930 15880
rect 2170 15640 2260 15880
rect 2500 15640 2590 15880
rect 2830 15640 2920 15880
rect 3160 15640 3250 15880
rect 3490 15640 3580 15880
rect 3820 15640 3910 15880
rect 4150 15640 4240 15880
rect 4480 15640 4570 15880
rect 4810 15640 4900 15880
rect 5140 15640 5230 15880
rect 5470 15640 5560 15880
rect 5800 15640 5890 15880
rect 6130 15640 6220 15880
rect 6460 15640 6550 15880
rect 6790 15640 6880 15880
rect 7120 15640 7260 15880
rect -4980 15550 7260 15640
rect -4980 15310 -4670 15550
rect -4430 15310 -4340 15550
rect -4100 15310 -4010 15550
rect -3770 15310 -3680 15550
rect -3440 15310 -3350 15550
rect -3110 15310 -3020 15550
rect -2780 15310 -2690 15550
rect -2450 15310 -2360 15550
rect -2120 15310 -2030 15550
rect -1790 15310 -1700 15550
rect -1460 15310 -1370 15550
rect -1130 15310 -1040 15550
rect -800 15310 -710 15550
rect -470 15310 -380 15550
rect -140 15310 -50 15550
rect 190 15310 280 15550
rect 520 15310 610 15550
rect 850 15310 940 15550
rect 1180 15310 1270 15550
rect 1510 15310 1600 15550
rect 1840 15310 1930 15550
rect 2170 15310 2260 15550
rect 2500 15310 2590 15550
rect 2830 15310 2920 15550
rect 3160 15310 3250 15550
rect 3490 15310 3580 15550
rect 3820 15310 3910 15550
rect 4150 15310 4240 15550
rect 4480 15310 4570 15550
rect 4810 15310 4900 15550
rect 5140 15310 5230 15550
rect 5470 15310 5560 15550
rect 5800 15310 5890 15550
rect 6130 15310 6220 15550
rect 6460 15310 6550 15550
rect 6790 15310 6880 15550
rect 7120 15310 7260 15550
rect -4980 15220 7260 15310
rect -4980 14980 -4670 15220
rect -4430 14980 -4340 15220
rect -4100 14980 -4010 15220
rect -3770 14980 -3680 15220
rect -3440 14980 -3350 15220
rect -3110 14980 -3020 15220
rect -2780 14980 -2690 15220
rect -2450 14980 -2360 15220
rect -2120 14980 -2030 15220
rect -1790 14980 -1700 15220
rect -1460 14980 -1370 15220
rect -1130 14980 -1040 15220
rect -800 14980 -710 15220
rect -470 14980 -380 15220
rect -140 14980 -50 15220
rect 190 14980 280 15220
rect 520 14980 610 15220
rect 850 14980 940 15220
rect 1180 14980 1270 15220
rect 1510 14980 1600 15220
rect 1840 14980 1930 15220
rect 2170 14980 2260 15220
rect 2500 14980 2590 15220
rect 2830 14980 2920 15220
rect 3160 14980 3250 15220
rect 3490 14980 3580 15220
rect 3820 14980 3910 15220
rect 4150 14980 4240 15220
rect 4480 14980 4570 15220
rect 4810 14980 4900 15220
rect 5140 14980 5230 15220
rect 5470 14980 5560 15220
rect 5800 14980 5890 15220
rect 6130 14980 6220 15220
rect 6460 14980 6550 15220
rect 6790 14980 6880 15220
rect 7120 14980 7260 15220
rect -4980 14890 7260 14980
rect -4980 14650 -4670 14890
rect -4430 14650 -4340 14890
rect -4100 14650 -4010 14890
rect -3770 14650 -3680 14890
rect -3440 14650 -3350 14890
rect -3110 14650 -3020 14890
rect -2780 14650 -2690 14890
rect -2450 14650 -2360 14890
rect -2120 14650 -2030 14890
rect -1790 14650 -1700 14890
rect -1460 14650 -1370 14890
rect -1130 14650 -1040 14890
rect -800 14650 -710 14890
rect -470 14650 -380 14890
rect -140 14650 -50 14890
rect 190 14650 280 14890
rect 520 14650 610 14890
rect 850 14650 940 14890
rect 1180 14650 1270 14890
rect 1510 14650 1600 14890
rect 1840 14650 1930 14890
rect 2170 14650 2260 14890
rect 2500 14650 2590 14890
rect 2830 14650 2920 14890
rect 3160 14650 3250 14890
rect 3490 14650 3580 14890
rect 3820 14650 3910 14890
rect 4150 14650 4240 14890
rect 4480 14650 4570 14890
rect 4810 14650 4900 14890
rect 5140 14650 5230 14890
rect 5470 14650 5560 14890
rect 5800 14650 5890 14890
rect 6130 14650 6220 14890
rect 6460 14650 6550 14890
rect 6790 14650 6880 14890
rect 7120 14650 7260 14890
rect -4980 14560 7260 14650
rect -4980 14320 -4670 14560
rect -4430 14320 -4340 14560
rect -4100 14320 -4010 14560
rect -3770 14320 -3680 14560
rect -3440 14320 -3350 14560
rect -3110 14320 -3020 14560
rect -2780 14320 -2690 14560
rect -2450 14320 -2360 14560
rect -2120 14320 -2030 14560
rect -1790 14320 -1700 14560
rect -1460 14320 -1370 14560
rect -1130 14320 -1040 14560
rect -800 14320 -710 14560
rect -470 14320 -380 14560
rect -140 14320 -50 14560
rect 190 14320 280 14560
rect 520 14320 610 14560
rect 850 14320 940 14560
rect 1180 14320 1270 14560
rect 1510 14320 1600 14560
rect 1840 14320 1930 14560
rect 2170 14320 2260 14560
rect 2500 14320 2590 14560
rect 2830 14320 2920 14560
rect 3160 14320 3250 14560
rect 3490 14320 3580 14560
rect 3820 14320 3910 14560
rect 4150 14320 4240 14560
rect 4480 14320 4570 14560
rect 4810 14320 4900 14560
rect 5140 14320 5230 14560
rect 5470 14320 5560 14560
rect 5800 14320 5890 14560
rect 6130 14320 6220 14560
rect 6460 14320 6550 14560
rect 6790 14320 6880 14560
rect 7120 14320 7260 14560
rect -4980 14230 7260 14320
rect -4980 13990 -4670 14230
rect -4430 13990 -4340 14230
rect -4100 13990 -4010 14230
rect -3770 13990 -3680 14230
rect -3440 13990 -3350 14230
rect -3110 13990 -3020 14230
rect -2780 13990 -2690 14230
rect -2450 13990 -2360 14230
rect -2120 13990 -2030 14230
rect -1790 13990 -1700 14230
rect -1460 13990 -1370 14230
rect -1130 13990 -1040 14230
rect -800 13990 -710 14230
rect -470 13990 -380 14230
rect -140 13990 -50 14230
rect 190 13990 280 14230
rect 520 13990 610 14230
rect 850 13990 940 14230
rect 1180 13990 1270 14230
rect 1510 13990 1600 14230
rect 1840 13990 1930 14230
rect 2170 13990 2260 14230
rect 2500 13990 2590 14230
rect 2830 13990 2920 14230
rect 3160 13990 3250 14230
rect 3490 13990 3580 14230
rect 3820 13990 3910 14230
rect 4150 13990 4240 14230
rect 4480 13990 4570 14230
rect 4810 13990 4900 14230
rect 5140 13990 5230 14230
rect 5470 13990 5560 14230
rect 5800 13990 5890 14230
rect 6130 13990 6220 14230
rect 6460 13990 6550 14230
rect 6790 13990 6880 14230
rect 7120 13990 7260 14230
rect -4980 13900 7260 13990
rect -4980 13660 -4670 13900
rect -4430 13660 -4340 13900
rect -4100 13660 -4010 13900
rect -3770 13660 -3680 13900
rect -3440 13660 -3350 13900
rect -3110 13660 -3020 13900
rect -2780 13660 -2690 13900
rect -2450 13660 -2360 13900
rect -2120 13660 -2030 13900
rect -1790 13660 -1700 13900
rect -1460 13660 -1370 13900
rect -1130 13660 -1040 13900
rect -800 13660 -710 13900
rect -470 13660 -380 13900
rect -140 13660 -50 13900
rect 190 13660 280 13900
rect 520 13660 610 13900
rect 850 13660 940 13900
rect 1180 13660 1270 13900
rect 1510 13660 1600 13900
rect 1840 13660 1930 13900
rect 2170 13660 2260 13900
rect 2500 13660 2590 13900
rect 2830 13660 2920 13900
rect 3160 13660 3250 13900
rect 3490 13660 3580 13900
rect 3820 13660 3910 13900
rect 4150 13660 4240 13900
rect 4480 13660 4570 13900
rect 4810 13660 4900 13900
rect 5140 13660 5230 13900
rect 5470 13660 5560 13900
rect 5800 13660 5890 13900
rect 6130 13660 6220 13900
rect 6460 13660 6550 13900
rect 6790 13660 6880 13900
rect 7120 13660 7260 13900
rect -4980 13570 7260 13660
rect -4980 13330 -4670 13570
rect -4430 13330 -4340 13570
rect -4100 13330 -4010 13570
rect -3770 13330 -3680 13570
rect -3440 13330 -3350 13570
rect -3110 13330 -3020 13570
rect -2780 13330 -2690 13570
rect -2450 13330 -2360 13570
rect -2120 13330 -2030 13570
rect -1790 13330 -1700 13570
rect -1460 13330 -1370 13570
rect -1130 13330 -1040 13570
rect -800 13330 -710 13570
rect -470 13330 -380 13570
rect -140 13330 -50 13570
rect 190 13330 280 13570
rect 520 13330 610 13570
rect 850 13330 940 13570
rect 1180 13330 1270 13570
rect 1510 13330 1600 13570
rect 1840 13330 1930 13570
rect 2170 13330 2260 13570
rect 2500 13330 2590 13570
rect 2830 13330 2920 13570
rect 3160 13330 3250 13570
rect 3490 13330 3580 13570
rect 3820 13330 3910 13570
rect 4150 13330 4240 13570
rect 4480 13330 4570 13570
rect 4810 13330 4900 13570
rect 5140 13330 5230 13570
rect 5470 13330 5560 13570
rect 5800 13330 5890 13570
rect 6130 13330 6220 13570
rect 6460 13330 6550 13570
rect 6790 13330 6880 13570
rect 7120 13330 7260 13570
rect -4980 13240 7260 13330
rect -4980 13000 -4670 13240
rect -4430 13000 -4340 13240
rect -4100 13000 -4010 13240
rect -3770 13000 -3680 13240
rect -3440 13000 -3350 13240
rect -3110 13000 -3020 13240
rect -2780 13000 -2690 13240
rect -2450 13000 -2360 13240
rect -2120 13000 -2030 13240
rect -1790 13000 -1700 13240
rect -1460 13000 -1370 13240
rect -1130 13000 -1040 13240
rect -800 13000 -710 13240
rect -470 13000 -380 13240
rect -140 13000 -50 13240
rect 190 13000 280 13240
rect 520 13000 610 13240
rect 850 13000 940 13240
rect 1180 13000 1270 13240
rect 1510 13000 1600 13240
rect 1840 13000 1930 13240
rect 2170 13000 2260 13240
rect 2500 13000 2590 13240
rect 2830 13000 2920 13240
rect 3160 13000 3250 13240
rect 3490 13000 3580 13240
rect 3820 13000 3910 13240
rect 4150 13000 4240 13240
rect 4480 13000 4570 13240
rect 4810 13000 4900 13240
rect 5140 13000 5230 13240
rect 5470 13000 5560 13240
rect 5800 13000 5890 13240
rect 6130 13000 6220 13240
rect 6460 13000 6550 13240
rect 6790 13000 6880 13240
rect 7120 13000 7260 13240
rect -4980 12910 7260 13000
rect -4980 12670 -4670 12910
rect -4430 12670 -4340 12910
rect -4100 12670 -4010 12910
rect -3770 12670 -3680 12910
rect -3440 12670 -3350 12910
rect -3110 12670 -3020 12910
rect -2780 12670 -2690 12910
rect -2450 12670 -2360 12910
rect -2120 12670 -2030 12910
rect -1790 12670 -1700 12910
rect -1460 12670 -1370 12910
rect -1130 12670 -1040 12910
rect -800 12670 -710 12910
rect -470 12670 -380 12910
rect -140 12670 -50 12910
rect 190 12670 280 12910
rect 520 12670 610 12910
rect 850 12670 940 12910
rect 1180 12670 1270 12910
rect 1510 12670 1600 12910
rect 1840 12670 1930 12910
rect 2170 12670 2260 12910
rect 2500 12670 2590 12910
rect 2830 12670 2920 12910
rect 3160 12670 3250 12910
rect 3490 12670 3580 12910
rect 3820 12670 3910 12910
rect 4150 12670 4240 12910
rect 4480 12670 4570 12910
rect 4810 12670 4900 12910
rect 5140 12670 5230 12910
rect 5470 12670 5560 12910
rect 5800 12670 5890 12910
rect 6130 12670 6220 12910
rect 6460 12670 6550 12910
rect 6790 12670 6880 12910
rect 7120 12670 7260 12910
rect -4980 12580 7260 12670
rect -4980 12340 -4670 12580
rect -4430 12340 -4340 12580
rect -4100 12340 -4010 12580
rect -3770 12340 -3680 12580
rect -3440 12340 -3350 12580
rect -3110 12340 -3020 12580
rect -2780 12340 -2690 12580
rect -2450 12340 -2360 12580
rect -2120 12340 -2030 12580
rect -1790 12340 -1700 12580
rect -1460 12340 -1370 12580
rect -1130 12340 -1040 12580
rect -800 12340 -710 12580
rect -470 12340 -380 12580
rect -140 12340 -50 12580
rect 190 12340 280 12580
rect 520 12340 610 12580
rect 850 12340 940 12580
rect 1180 12340 1270 12580
rect 1510 12340 1600 12580
rect 1840 12340 1930 12580
rect 2170 12340 2260 12580
rect 2500 12340 2590 12580
rect 2830 12340 2920 12580
rect 3160 12340 3250 12580
rect 3490 12340 3580 12580
rect 3820 12340 3910 12580
rect 4150 12340 4240 12580
rect 4480 12340 4570 12580
rect 4810 12340 4900 12580
rect 5140 12340 5230 12580
rect 5470 12340 5560 12580
rect 5800 12340 5890 12580
rect 6130 12340 6220 12580
rect 6460 12340 6550 12580
rect 6790 12340 6880 12580
rect 7120 12340 7260 12580
rect -4980 12250 7260 12340
rect -4980 12010 -4670 12250
rect -4430 12010 -4340 12250
rect -4100 12010 -4010 12250
rect -3770 12010 -3680 12250
rect -3440 12010 -3350 12250
rect -3110 12010 -3020 12250
rect -2780 12010 -2690 12250
rect -2450 12010 -2360 12250
rect -2120 12010 -2030 12250
rect -1790 12010 -1700 12250
rect -1460 12010 -1370 12250
rect -1130 12010 -1040 12250
rect -800 12010 -710 12250
rect -470 12010 -380 12250
rect -140 12010 -50 12250
rect 190 12010 280 12250
rect 520 12010 610 12250
rect 850 12010 940 12250
rect 1180 12010 1270 12250
rect 1510 12010 1600 12250
rect 1840 12010 1930 12250
rect 2170 12010 2260 12250
rect 2500 12010 2590 12250
rect 2830 12010 2920 12250
rect 3160 12010 3250 12250
rect 3490 12010 3580 12250
rect 3820 12010 3910 12250
rect 4150 12010 4240 12250
rect 4480 12010 4570 12250
rect 4810 12010 4900 12250
rect 5140 12010 5230 12250
rect 5470 12010 5560 12250
rect 5800 12010 5890 12250
rect 6130 12010 6220 12250
rect 6460 12010 6550 12250
rect 6790 12010 6880 12250
rect 7120 12010 7260 12250
rect -4980 11920 7260 12010
rect -4980 11680 -4670 11920
rect -4430 11680 -4340 11920
rect -4100 11680 -4010 11920
rect -3770 11680 -3680 11920
rect -3440 11680 -3350 11920
rect -3110 11680 -3020 11920
rect -2780 11680 -2690 11920
rect -2450 11680 -2360 11920
rect -2120 11680 -2030 11920
rect -1790 11680 -1700 11920
rect -1460 11680 -1370 11920
rect -1130 11680 -1040 11920
rect -800 11680 -710 11920
rect -470 11680 -380 11920
rect -140 11680 -50 11920
rect 190 11680 280 11920
rect 520 11680 610 11920
rect 850 11680 940 11920
rect 1180 11680 1270 11920
rect 1510 11680 1600 11920
rect 1840 11680 1930 11920
rect 2170 11680 2260 11920
rect 2500 11680 2590 11920
rect 2830 11680 2920 11920
rect 3160 11680 3250 11920
rect 3490 11680 3580 11920
rect 3820 11680 3910 11920
rect 4150 11680 4240 11920
rect 4480 11680 4570 11920
rect 4810 11680 4900 11920
rect 5140 11680 5230 11920
rect 5470 11680 5560 11920
rect 5800 11680 5890 11920
rect 6130 11680 6220 11920
rect 6460 11680 6550 11920
rect 6790 11680 6880 11920
rect 7120 11680 7260 11920
rect -4980 11590 7260 11680
rect -4980 11350 -4670 11590
rect -4430 11350 -4340 11590
rect -4100 11350 -4010 11590
rect -3770 11350 -3680 11590
rect -3440 11350 -3350 11590
rect -3110 11350 -3020 11590
rect -2780 11350 -2690 11590
rect -2450 11350 -2360 11590
rect -2120 11350 -2030 11590
rect -1790 11350 -1700 11590
rect -1460 11350 -1370 11590
rect -1130 11350 -1040 11590
rect -800 11350 -710 11590
rect -470 11350 -380 11590
rect -140 11350 -50 11590
rect 190 11350 280 11590
rect 520 11350 610 11590
rect 850 11350 940 11590
rect 1180 11350 1270 11590
rect 1510 11350 1600 11590
rect 1840 11350 1930 11590
rect 2170 11350 2260 11590
rect 2500 11350 2590 11590
rect 2830 11350 2920 11590
rect 3160 11350 3250 11590
rect 3490 11350 3580 11590
rect 3820 11350 3910 11590
rect 4150 11350 4240 11590
rect 4480 11350 4570 11590
rect 4810 11350 4900 11590
rect 5140 11350 5230 11590
rect 5470 11350 5560 11590
rect 5800 11350 5890 11590
rect 6130 11350 6220 11590
rect 6460 11350 6550 11590
rect 6790 11350 6880 11590
rect 7120 11350 7260 11590
rect -4980 11260 7260 11350
rect -4980 11020 -4670 11260
rect -4430 11020 -4340 11260
rect -4100 11020 -4010 11260
rect -3770 11020 -3680 11260
rect -3440 11020 -3350 11260
rect -3110 11020 -3020 11260
rect -2780 11020 -2690 11260
rect -2450 11020 -2360 11260
rect -2120 11020 -2030 11260
rect -1790 11020 -1700 11260
rect -1460 11020 -1370 11260
rect -1130 11020 -1040 11260
rect -800 11020 -710 11260
rect -470 11020 -380 11260
rect -140 11020 -50 11260
rect 190 11020 280 11260
rect 520 11020 610 11260
rect 850 11020 940 11260
rect 1180 11020 1270 11260
rect 1510 11020 1600 11260
rect 1840 11020 1930 11260
rect 2170 11020 2260 11260
rect 2500 11020 2590 11260
rect 2830 11020 2920 11260
rect 3160 11020 3250 11260
rect 3490 11020 3580 11260
rect 3820 11020 3910 11260
rect 4150 11020 4240 11260
rect 4480 11020 4570 11260
rect 4810 11020 4900 11260
rect 5140 11020 5230 11260
rect 5470 11020 5560 11260
rect 5800 11020 5890 11260
rect 6130 11020 6220 11260
rect 6460 11020 6550 11260
rect 6790 11020 6880 11260
rect 7120 11020 7260 11260
rect -4980 10930 7260 11020
rect -4980 10690 -4670 10930
rect -4430 10690 -4340 10930
rect -4100 10690 -4010 10930
rect -3770 10690 -3680 10930
rect -3440 10690 -3350 10930
rect -3110 10690 -3020 10930
rect -2780 10690 -2690 10930
rect -2450 10690 -2360 10930
rect -2120 10690 -2030 10930
rect -1790 10690 -1700 10930
rect -1460 10690 -1370 10930
rect -1130 10690 -1040 10930
rect -800 10690 -710 10930
rect -470 10690 -380 10930
rect -140 10690 -50 10930
rect 190 10690 280 10930
rect 520 10690 610 10930
rect 850 10690 940 10930
rect 1180 10690 1270 10930
rect 1510 10690 1600 10930
rect 1840 10690 1930 10930
rect 2170 10690 2260 10930
rect 2500 10690 2590 10930
rect 2830 10690 2920 10930
rect 3160 10690 3250 10930
rect 3490 10690 3580 10930
rect 3820 10690 3910 10930
rect 4150 10690 4240 10930
rect 4480 10690 4570 10930
rect 4810 10690 4900 10930
rect 5140 10690 5230 10930
rect 5470 10690 5560 10930
rect 5800 10690 5890 10930
rect 6130 10690 6220 10930
rect 6460 10690 6550 10930
rect 6790 10690 6880 10930
rect 7120 10690 7260 10930
rect -4980 10600 7260 10690
rect -4980 10360 -4670 10600
rect -4430 10360 -4340 10600
rect -4100 10360 -4010 10600
rect -3770 10360 -3680 10600
rect -3440 10360 -3350 10600
rect -3110 10360 -3020 10600
rect -2780 10360 -2690 10600
rect -2450 10360 -2360 10600
rect -2120 10360 -2030 10600
rect -1790 10360 -1700 10600
rect -1460 10360 -1370 10600
rect -1130 10360 -1040 10600
rect -800 10360 -710 10600
rect -470 10360 -380 10600
rect -140 10360 -50 10600
rect 190 10360 280 10600
rect 520 10360 610 10600
rect 850 10360 940 10600
rect 1180 10360 1270 10600
rect 1510 10360 1600 10600
rect 1840 10360 1930 10600
rect 2170 10360 2260 10600
rect 2500 10360 2590 10600
rect 2830 10360 2920 10600
rect 3160 10360 3250 10600
rect 3490 10360 3580 10600
rect 3820 10360 3910 10600
rect 4150 10360 4240 10600
rect 4480 10360 4570 10600
rect 4810 10360 4900 10600
rect 5140 10360 5230 10600
rect 5470 10360 5560 10600
rect 5800 10360 5890 10600
rect 6130 10360 6220 10600
rect 6460 10360 6550 10600
rect 6790 10360 6880 10600
rect 7120 10360 7260 10600
rect -4980 10270 7260 10360
rect -4980 10030 -4670 10270
rect -4430 10030 -4340 10270
rect -4100 10030 -4010 10270
rect -3770 10030 -3680 10270
rect -3440 10030 -3350 10270
rect -3110 10030 -3020 10270
rect -2780 10030 -2690 10270
rect -2450 10030 -2360 10270
rect -2120 10030 -2030 10270
rect -1790 10030 -1700 10270
rect -1460 10030 -1370 10270
rect -1130 10030 -1040 10270
rect -800 10030 -710 10270
rect -470 10030 -380 10270
rect -140 10030 -50 10270
rect 190 10030 280 10270
rect 520 10030 610 10270
rect 850 10030 940 10270
rect 1180 10030 1270 10270
rect 1510 10030 1600 10270
rect 1840 10030 1930 10270
rect 2170 10030 2260 10270
rect 2500 10030 2590 10270
rect 2830 10030 2920 10270
rect 3160 10030 3250 10270
rect 3490 10030 3580 10270
rect 3820 10030 3910 10270
rect 4150 10030 4240 10270
rect 4480 10030 4570 10270
rect 4810 10030 4900 10270
rect 5140 10030 5230 10270
rect 5470 10030 5560 10270
rect 5800 10030 5890 10270
rect 6130 10030 6220 10270
rect 6460 10030 6550 10270
rect 6790 10030 6880 10270
rect 7120 10030 7260 10270
rect -4980 9940 7260 10030
rect -4980 9700 -4670 9940
rect -4430 9700 -4340 9940
rect -4100 9700 -4010 9940
rect -3770 9700 -3680 9940
rect -3440 9700 -3350 9940
rect -3110 9700 -3020 9940
rect -2780 9700 -2690 9940
rect -2450 9700 -2360 9940
rect -2120 9700 -2030 9940
rect -1790 9700 -1700 9940
rect -1460 9700 -1370 9940
rect -1130 9700 -1040 9940
rect -800 9700 -710 9940
rect -470 9700 -380 9940
rect -140 9700 -50 9940
rect 190 9700 280 9940
rect 520 9700 610 9940
rect 850 9700 940 9940
rect 1180 9700 1270 9940
rect 1510 9700 1600 9940
rect 1840 9700 1930 9940
rect 2170 9700 2260 9940
rect 2500 9700 2590 9940
rect 2830 9700 2920 9940
rect 3160 9700 3250 9940
rect 3490 9700 3580 9940
rect 3820 9700 3910 9940
rect 4150 9700 4240 9940
rect 4480 9700 4570 9940
rect 4810 9700 4900 9940
rect 5140 9700 5230 9940
rect 5470 9700 5560 9940
rect 5800 9700 5890 9940
rect 6130 9700 6220 9940
rect 6460 9700 6550 9940
rect 6790 9700 6880 9940
rect 7120 9700 7260 9940
rect -4980 9610 7260 9700
rect -4980 9370 -4670 9610
rect -4430 9370 -4340 9610
rect -4100 9370 -4010 9610
rect -3770 9370 -3680 9610
rect -3440 9370 -3350 9610
rect -3110 9370 -3020 9610
rect -2780 9370 -2690 9610
rect -2450 9370 -2360 9610
rect -2120 9370 -2030 9610
rect -1790 9370 -1700 9610
rect -1460 9370 -1370 9610
rect -1130 9370 -1040 9610
rect -800 9370 -710 9610
rect -470 9370 -380 9610
rect -140 9370 -50 9610
rect 190 9370 280 9610
rect 520 9370 610 9610
rect 850 9370 940 9610
rect 1180 9370 1270 9610
rect 1510 9370 1600 9610
rect 1840 9370 1930 9610
rect 2170 9370 2260 9610
rect 2500 9370 2590 9610
rect 2830 9370 2920 9610
rect 3160 9370 3250 9610
rect 3490 9370 3580 9610
rect 3820 9370 3910 9610
rect 4150 9370 4240 9610
rect 4480 9370 4570 9610
rect 4810 9370 4900 9610
rect 5140 9370 5230 9610
rect 5470 9370 5560 9610
rect 5800 9370 5890 9610
rect 6130 9370 6220 9610
rect 6460 9370 6550 9610
rect 6790 9370 6880 9610
rect 7120 9370 7260 9610
rect -4980 9280 7260 9370
rect -4980 9040 -4670 9280
rect -4430 9040 -4340 9280
rect -4100 9040 -4010 9280
rect -3770 9040 -3680 9280
rect -3440 9040 -3350 9280
rect -3110 9040 -3020 9280
rect -2780 9040 -2690 9280
rect -2450 9040 -2360 9280
rect -2120 9040 -2030 9280
rect -1790 9040 -1700 9280
rect -1460 9040 -1370 9280
rect -1130 9040 -1040 9280
rect -800 9040 -710 9280
rect -470 9040 -380 9280
rect -140 9040 -50 9280
rect 190 9040 280 9280
rect 520 9040 610 9280
rect 850 9040 940 9280
rect 1180 9040 1270 9280
rect 1510 9040 1600 9280
rect 1840 9040 1930 9280
rect 2170 9040 2260 9280
rect 2500 9040 2590 9280
rect 2830 9040 2920 9280
rect 3160 9040 3250 9280
rect 3490 9040 3580 9280
rect 3820 9040 3910 9280
rect 4150 9040 4240 9280
rect 4480 9040 4570 9280
rect 4810 9040 4900 9280
rect 5140 9040 5230 9280
rect 5470 9040 5560 9280
rect 5800 9040 5890 9280
rect 6130 9040 6220 9280
rect 6460 9040 6550 9280
rect 6790 9040 6880 9280
rect 7120 9040 7260 9280
rect -4980 8720 7260 9040
rect 7640 20830 19880 20960
rect 7640 20590 7780 20830
rect 8020 20590 8110 20830
rect 8350 20590 8440 20830
rect 8680 20590 8770 20830
rect 9010 20590 9100 20830
rect 9340 20590 9430 20830
rect 9670 20590 9760 20830
rect 10000 20590 10090 20830
rect 10330 20590 10420 20830
rect 10660 20590 10750 20830
rect 10990 20590 11080 20830
rect 11320 20590 11410 20830
rect 11650 20590 11740 20830
rect 11980 20590 12070 20830
rect 12310 20590 12400 20830
rect 12640 20590 12730 20830
rect 12970 20590 13060 20830
rect 13300 20590 13390 20830
rect 13630 20590 13720 20830
rect 13960 20590 14050 20830
rect 14290 20590 14380 20830
rect 14620 20590 14710 20830
rect 14950 20590 15040 20830
rect 15280 20590 15370 20830
rect 15610 20590 15700 20830
rect 15940 20590 16030 20830
rect 16270 20590 16360 20830
rect 16600 20590 16690 20830
rect 16930 20590 17020 20830
rect 17260 20590 17350 20830
rect 17590 20590 17680 20830
rect 17920 20590 18010 20830
rect 18250 20590 18340 20830
rect 18580 20590 18670 20830
rect 18910 20590 19000 20830
rect 19240 20590 19330 20830
rect 19570 20590 19880 20830
rect 7640 20500 19880 20590
rect 7640 20260 7780 20500
rect 8020 20260 8110 20500
rect 8350 20260 8440 20500
rect 8680 20260 8770 20500
rect 9010 20260 9100 20500
rect 9340 20260 9430 20500
rect 9670 20260 9760 20500
rect 10000 20260 10090 20500
rect 10330 20260 10420 20500
rect 10660 20260 10750 20500
rect 10990 20260 11080 20500
rect 11320 20260 11410 20500
rect 11650 20260 11740 20500
rect 11980 20260 12070 20500
rect 12310 20260 12400 20500
rect 12640 20260 12730 20500
rect 12970 20260 13060 20500
rect 13300 20260 13390 20500
rect 13630 20260 13720 20500
rect 13960 20260 14050 20500
rect 14290 20260 14380 20500
rect 14620 20260 14710 20500
rect 14950 20260 15040 20500
rect 15280 20260 15370 20500
rect 15610 20260 15700 20500
rect 15940 20260 16030 20500
rect 16270 20260 16360 20500
rect 16600 20260 16690 20500
rect 16930 20260 17020 20500
rect 17260 20260 17350 20500
rect 17590 20260 17680 20500
rect 17920 20260 18010 20500
rect 18250 20260 18340 20500
rect 18580 20260 18670 20500
rect 18910 20260 19000 20500
rect 19240 20260 19330 20500
rect 19570 20260 19880 20500
rect 7640 20170 19880 20260
rect 7640 19930 7780 20170
rect 8020 19930 8110 20170
rect 8350 19930 8440 20170
rect 8680 19930 8770 20170
rect 9010 19930 9100 20170
rect 9340 19930 9430 20170
rect 9670 19930 9760 20170
rect 10000 19930 10090 20170
rect 10330 19930 10420 20170
rect 10660 19930 10750 20170
rect 10990 19930 11080 20170
rect 11320 19930 11410 20170
rect 11650 19930 11740 20170
rect 11980 19930 12070 20170
rect 12310 19930 12400 20170
rect 12640 19930 12730 20170
rect 12970 19930 13060 20170
rect 13300 19930 13390 20170
rect 13630 19930 13720 20170
rect 13960 19930 14050 20170
rect 14290 19930 14380 20170
rect 14620 19930 14710 20170
rect 14950 19930 15040 20170
rect 15280 19930 15370 20170
rect 15610 19930 15700 20170
rect 15940 19930 16030 20170
rect 16270 19930 16360 20170
rect 16600 19930 16690 20170
rect 16930 19930 17020 20170
rect 17260 19930 17350 20170
rect 17590 19930 17680 20170
rect 17920 19930 18010 20170
rect 18250 19930 18340 20170
rect 18580 19930 18670 20170
rect 18910 19930 19000 20170
rect 19240 19930 19330 20170
rect 19570 19930 19880 20170
rect 7640 19840 19880 19930
rect 7640 19600 7780 19840
rect 8020 19600 8110 19840
rect 8350 19600 8440 19840
rect 8680 19600 8770 19840
rect 9010 19600 9100 19840
rect 9340 19600 9430 19840
rect 9670 19600 9760 19840
rect 10000 19600 10090 19840
rect 10330 19600 10420 19840
rect 10660 19600 10750 19840
rect 10990 19600 11080 19840
rect 11320 19600 11410 19840
rect 11650 19600 11740 19840
rect 11980 19600 12070 19840
rect 12310 19600 12400 19840
rect 12640 19600 12730 19840
rect 12970 19600 13060 19840
rect 13300 19600 13390 19840
rect 13630 19600 13720 19840
rect 13960 19600 14050 19840
rect 14290 19600 14380 19840
rect 14620 19600 14710 19840
rect 14950 19600 15040 19840
rect 15280 19600 15370 19840
rect 15610 19600 15700 19840
rect 15940 19600 16030 19840
rect 16270 19600 16360 19840
rect 16600 19600 16690 19840
rect 16930 19600 17020 19840
rect 17260 19600 17350 19840
rect 17590 19600 17680 19840
rect 17920 19600 18010 19840
rect 18250 19600 18340 19840
rect 18580 19600 18670 19840
rect 18910 19600 19000 19840
rect 19240 19600 19330 19840
rect 19570 19600 19880 19840
rect 7640 19510 19880 19600
rect 7640 19270 7780 19510
rect 8020 19270 8110 19510
rect 8350 19270 8440 19510
rect 8680 19270 8770 19510
rect 9010 19270 9100 19510
rect 9340 19270 9430 19510
rect 9670 19270 9760 19510
rect 10000 19270 10090 19510
rect 10330 19270 10420 19510
rect 10660 19270 10750 19510
rect 10990 19270 11080 19510
rect 11320 19270 11410 19510
rect 11650 19270 11740 19510
rect 11980 19270 12070 19510
rect 12310 19270 12400 19510
rect 12640 19270 12730 19510
rect 12970 19270 13060 19510
rect 13300 19270 13390 19510
rect 13630 19270 13720 19510
rect 13960 19270 14050 19510
rect 14290 19270 14380 19510
rect 14620 19270 14710 19510
rect 14950 19270 15040 19510
rect 15280 19270 15370 19510
rect 15610 19270 15700 19510
rect 15940 19270 16030 19510
rect 16270 19270 16360 19510
rect 16600 19270 16690 19510
rect 16930 19270 17020 19510
rect 17260 19270 17350 19510
rect 17590 19270 17680 19510
rect 17920 19270 18010 19510
rect 18250 19270 18340 19510
rect 18580 19270 18670 19510
rect 18910 19270 19000 19510
rect 19240 19270 19330 19510
rect 19570 19270 19880 19510
rect 7640 19180 19880 19270
rect 7640 18940 7780 19180
rect 8020 18940 8110 19180
rect 8350 18940 8440 19180
rect 8680 18940 8770 19180
rect 9010 18940 9100 19180
rect 9340 18940 9430 19180
rect 9670 18940 9760 19180
rect 10000 18940 10090 19180
rect 10330 18940 10420 19180
rect 10660 18940 10750 19180
rect 10990 18940 11080 19180
rect 11320 18940 11410 19180
rect 11650 18940 11740 19180
rect 11980 18940 12070 19180
rect 12310 18940 12400 19180
rect 12640 18940 12730 19180
rect 12970 18940 13060 19180
rect 13300 18940 13390 19180
rect 13630 18940 13720 19180
rect 13960 18940 14050 19180
rect 14290 18940 14380 19180
rect 14620 18940 14710 19180
rect 14950 18940 15040 19180
rect 15280 18940 15370 19180
rect 15610 18940 15700 19180
rect 15940 18940 16030 19180
rect 16270 18940 16360 19180
rect 16600 18940 16690 19180
rect 16930 18940 17020 19180
rect 17260 18940 17350 19180
rect 17590 18940 17680 19180
rect 17920 18940 18010 19180
rect 18250 18940 18340 19180
rect 18580 18940 18670 19180
rect 18910 18940 19000 19180
rect 19240 18940 19330 19180
rect 19570 18940 19880 19180
rect 7640 18850 19880 18940
rect 7640 18610 7780 18850
rect 8020 18610 8110 18850
rect 8350 18610 8440 18850
rect 8680 18610 8770 18850
rect 9010 18610 9100 18850
rect 9340 18610 9430 18850
rect 9670 18610 9760 18850
rect 10000 18610 10090 18850
rect 10330 18610 10420 18850
rect 10660 18610 10750 18850
rect 10990 18610 11080 18850
rect 11320 18610 11410 18850
rect 11650 18610 11740 18850
rect 11980 18610 12070 18850
rect 12310 18610 12400 18850
rect 12640 18610 12730 18850
rect 12970 18610 13060 18850
rect 13300 18610 13390 18850
rect 13630 18610 13720 18850
rect 13960 18610 14050 18850
rect 14290 18610 14380 18850
rect 14620 18610 14710 18850
rect 14950 18610 15040 18850
rect 15280 18610 15370 18850
rect 15610 18610 15700 18850
rect 15940 18610 16030 18850
rect 16270 18610 16360 18850
rect 16600 18610 16690 18850
rect 16930 18610 17020 18850
rect 17260 18610 17350 18850
rect 17590 18610 17680 18850
rect 17920 18610 18010 18850
rect 18250 18610 18340 18850
rect 18580 18610 18670 18850
rect 18910 18610 19000 18850
rect 19240 18610 19330 18850
rect 19570 18610 19880 18850
rect 7640 18520 19880 18610
rect 7640 18280 7780 18520
rect 8020 18280 8110 18520
rect 8350 18280 8440 18520
rect 8680 18280 8770 18520
rect 9010 18280 9100 18520
rect 9340 18280 9430 18520
rect 9670 18280 9760 18520
rect 10000 18280 10090 18520
rect 10330 18280 10420 18520
rect 10660 18280 10750 18520
rect 10990 18280 11080 18520
rect 11320 18280 11410 18520
rect 11650 18280 11740 18520
rect 11980 18280 12070 18520
rect 12310 18280 12400 18520
rect 12640 18280 12730 18520
rect 12970 18280 13060 18520
rect 13300 18280 13390 18520
rect 13630 18280 13720 18520
rect 13960 18280 14050 18520
rect 14290 18280 14380 18520
rect 14620 18280 14710 18520
rect 14950 18280 15040 18520
rect 15280 18280 15370 18520
rect 15610 18280 15700 18520
rect 15940 18280 16030 18520
rect 16270 18280 16360 18520
rect 16600 18280 16690 18520
rect 16930 18280 17020 18520
rect 17260 18280 17350 18520
rect 17590 18280 17680 18520
rect 17920 18280 18010 18520
rect 18250 18280 18340 18520
rect 18580 18280 18670 18520
rect 18910 18280 19000 18520
rect 19240 18280 19330 18520
rect 19570 18280 19880 18520
rect 7640 18190 19880 18280
rect 7640 17950 7780 18190
rect 8020 17950 8110 18190
rect 8350 17950 8440 18190
rect 8680 17950 8770 18190
rect 9010 17950 9100 18190
rect 9340 17950 9430 18190
rect 9670 17950 9760 18190
rect 10000 17950 10090 18190
rect 10330 17950 10420 18190
rect 10660 17950 10750 18190
rect 10990 17950 11080 18190
rect 11320 17950 11410 18190
rect 11650 17950 11740 18190
rect 11980 17950 12070 18190
rect 12310 17950 12400 18190
rect 12640 17950 12730 18190
rect 12970 17950 13060 18190
rect 13300 17950 13390 18190
rect 13630 17950 13720 18190
rect 13960 17950 14050 18190
rect 14290 17950 14380 18190
rect 14620 17950 14710 18190
rect 14950 17950 15040 18190
rect 15280 17950 15370 18190
rect 15610 17950 15700 18190
rect 15940 17950 16030 18190
rect 16270 17950 16360 18190
rect 16600 17950 16690 18190
rect 16930 17950 17020 18190
rect 17260 17950 17350 18190
rect 17590 17950 17680 18190
rect 17920 17950 18010 18190
rect 18250 17950 18340 18190
rect 18580 17950 18670 18190
rect 18910 17950 19000 18190
rect 19240 17950 19330 18190
rect 19570 17950 19880 18190
rect 7640 17860 19880 17950
rect 7640 17620 7780 17860
rect 8020 17620 8110 17860
rect 8350 17620 8440 17860
rect 8680 17620 8770 17860
rect 9010 17620 9100 17860
rect 9340 17620 9430 17860
rect 9670 17620 9760 17860
rect 10000 17620 10090 17860
rect 10330 17620 10420 17860
rect 10660 17620 10750 17860
rect 10990 17620 11080 17860
rect 11320 17620 11410 17860
rect 11650 17620 11740 17860
rect 11980 17620 12070 17860
rect 12310 17620 12400 17860
rect 12640 17620 12730 17860
rect 12970 17620 13060 17860
rect 13300 17620 13390 17860
rect 13630 17620 13720 17860
rect 13960 17620 14050 17860
rect 14290 17620 14380 17860
rect 14620 17620 14710 17860
rect 14950 17620 15040 17860
rect 15280 17620 15370 17860
rect 15610 17620 15700 17860
rect 15940 17620 16030 17860
rect 16270 17620 16360 17860
rect 16600 17620 16690 17860
rect 16930 17620 17020 17860
rect 17260 17620 17350 17860
rect 17590 17620 17680 17860
rect 17920 17620 18010 17860
rect 18250 17620 18340 17860
rect 18580 17620 18670 17860
rect 18910 17620 19000 17860
rect 19240 17620 19330 17860
rect 19570 17620 19880 17860
rect 7640 17530 19880 17620
rect 7640 17290 7780 17530
rect 8020 17290 8110 17530
rect 8350 17290 8440 17530
rect 8680 17290 8770 17530
rect 9010 17290 9100 17530
rect 9340 17290 9430 17530
rect 9670 17290 9760 17530
rect 10000 17290 10090 17530
rect 10330 17290 10420 17530
rect 10660 17290 10750 17530
rect 10990 17290 11080 17530
rect 11320 17290 11410 17530
rect 11650 17290 11740 17530
rect 11980 17290 12070 17530
rect 12310 17290 12400 17530
rect 12640 17290 12730 17530
rect 12970 17290 13060 17530
rect 13300 17290 13390 17530
rect 13630 17290 13720 17530
rect 13960 17290 14050 17530
rect 14290 17290 14380 17530
rect 14620 17290 14710 17530
rect 14950 17290 15040 17530
rect 15280 17290 15370 17530
rect 15610 17290 15700 17530
rect 15940 17290 16030 17530
rect 16270 17290 16360 17530
rect 16600 17290 16690 17530
rect 16930 17290 17020 17530
rect 17260 17290 17350 17530
rect 17590 17290 17680 17530
rect 17920 17290 18010 17530
rect 18250 17290 18340 17530
rect 18580 17290 18670 17530
rect 18910 17290 19000 17530
rect 19240 17290 19330 17530
rect 19570 17290 19880 17530
rect 7640 17200 19880 17290
rect 7640 16960 7780 17200
rect 8020 16960 8110 17200
rect 8350 16960 8440 17200
rect 8680 16960 8770 17200
rect 9010 16960 9100 17200
rect 9340 16960 9430 17200
rect 9670 16960 9760 17200
rect 10000 16960 10090 17200
rect 10330 16960 10420 17200
rect 10660 16960 10750 17200
rect 10990 16960 11080 17200
rect 11320 16960 11410 17200
rect 11650 16960 11740 17200
rect 11980 16960 12070 17200
rect 12310 16960 12400 17200
rect 12640 16960 12730 17200
rect 12970 16960 13060 17200
rect 13300 16960 13390 17200
rect 13630 16960 13720 17200
rect 13960 16960 14050 17200
rect 14290 16960 14380 17200
rect 14620 16960 14710 17200
rect 14950 16960 15040 17200
rect 15280 16960 15370 17200
rect 15610 16960 15700 17200
rect 15940 16960 16030 17200
rect 16270 16960 16360 17200
rect 16600 16960 16690 17200
rect 16930 16960 17020 17200
rect 17260 16960 17350 17200
rect 17590 16960 17680 17200
rect 17920 16960 18010 17200
rect 18250 16960 18340 17200
rect 18580 16960 18670 17200
rect 18910 16960 19000 17200
rect 19240 16960 19330 17200
rect 19570 16960 19880 17200
rect 7640 16870 19880 16960
rect 7640 16630 7780 16870
rect 8020 16630 8110 16870
rect 8350 16630 8440 16870
rect 8680 16630 8770 16870
rect 9010 16630 9100 16870
rect 9340 16630 9430 16870
rect 9670 16630 9760 16870
rect 10000 16630 10090 16870
rect 10330 16630 10420 16870
rect 10660 16630 10750 16870
rect 10990 16630 11080 16870
rect 11320 16630 11410 16870
rect 11650 16630 11740 16870
rect 11980 16630 12070 16870
rect 12310 16630 12400 16870
rect 12640 16630 12730 16870
rect 12970 16630 13060 16870
rect 13300 16630 13390 16870
rect 13630 16630 13720 16870
rect 13960 16630 14050 16870
rect 14290 16630 14380 16870
rect 14620 16630 14710 16870
rect 14950 16630 15040 16870
rect 15280 16630 15370 16870
rect 15610 16630 15700 16870
rect 15940 16630 16030 16870
rect 16270 16630 16360 16870
rect 16600 16630 16690 16870
rect 16930 16630 17020 16870
rect 17260 16630 17350 16870
rect 17590 16630 17680 16870
rect 17920 16630 18010 16870
rect 18250 16630 18340 16870
rect 18580 16630 18670 16870
rect 18910 16630 19000 16870
rect 19240 16630 19330 16870
rect 19570 16630 19880 16870
rect 7640 16540 19880 16630
rect 7640 16300 7780 16540
rect 8020 16300 8110 16540
rect 8350 16300 8440 16540
rect 8680 16300 8770 16540
rect 9010 16300 9100 16540
rect 9340 16300 9430 16540
rect 9670 16300 9760 16540
rect 10000 16300 10090 16540
rect 10330 16300 10420 16540
rect 10660 16300 10750 16540
rect 10990 16300 11080 16540
rect 11320 16300 11410 16540
rect 11650 16300 11740 16540
rect 11980 16300 12070 16540
rect 12310 16300 12400 16540
rect 12640 16300 12730 16540
rect 12970 16300 13060 16540
rect 13300 16300 13390 16540
rect 13630 16300 13720 16540
rect 13960 16300 14050 16540
rect 14290 16300 14380 16540
rect 14620 16300 14710 16540
rect 14950 16300 15040 16540
rect 15280 16300 15370 16540
rect 15610 16300 15700 16540
rect 15940 16300 16030 16540
rect 16270 16300 16360 16540
rect 16600 16300 16690 16540
rect 16930 16300 17020 16540
rect 17260 16300 17350 16540
rect 17590 16300 17680 16540
rect 17920 16300 18010 16540
rect 18250 16300 18340 16540
rect 18580 16300 18670 16540
rect 18910 16300 19000 16540
rect 19240 16300 19330 16540
rect 19570 16300 19880 16540
rect 7640 16210 19880 16300
rect 7640 15970 7780 16210
rect 8020 15970 8110 16210
rect 8350 15970 8440 16210
rect 8680 15970 8770 16210
rect 9010 15970 9100 16210
rect 9340 15970 9430 16210
rect 9670 15970 9760 16210
rect 10000 15970 10090 16210
rect 10330 15970 10420 16210
rect 10660 15970 10750 16210
rect 10990 15970 11080 16210
rect 11320 15970 11410 16210
rect 11650 15970 11740 16210
rect 11980 15970 12070 16210
rect 12310 15970 12400 16210
rect 12640 15970 12730 16210
rect 12970 15970 13060 16210
rect 13300 15970 13390 16210
rect 13630 15970 13720 16210
rect 13960 15970 14050 16210
rect 14290 15970 14380 16210
rect 14620 15970 14710 16210
rect 14950 15970 15040 16210
rect 15280 15970 15370 16210
rect 15610 15970 15700 16210
rect 15940 15970 16030 16210
rect 16270 15970 16360 16210
rect 16600 15970 16690 16210
rect 16930 15970 17020 16210
rect 17260 15970 17350 16210
rect 17590 15970 17680 16210
rect 17920 15970 18010 16210
rect 18250 15970 18340 16210
rect 18580 15970 18670 16210
rect 18910 15970 19000 16210
rect 19240 15970 19330 16210
rect 19570 15970 19880 16210
rect 7640 15880 19880 15970
rect 7640 15640 7780 15880
rect 8020 15640 8110 15880
rect 8350 15640 8440 15880
rect 8680 15640 8770 15880
rect 9010 15640 9100 15880
rect 9340 15640 9430 15880
rect 9670 15640 9760 15880
rect 10000 15640 10090 15880
rect 10330 15640 10420 15880
rect 10660 15640 10750 15880
rect 10990 15640 11080 15880
rect 11320 15640 11410 15880
rect 11650 15640 11740 15880
rect 11980 15640 12070 15880
rect 12310 15640 12400 15880
rect 12640 15640 12730 15880
rect 12970 15640 13060 15880
rect 13300 15640 13390 15880
rect 13630 15640 13720 15880
rect 13960 15640 14050 15880
rect 14290 15640 14380 15880
rect 14620 15640 14710 15880
rect 14950 15640 15040 15880
rect 15280 15640 15370 15880
rect 15610 15640 15700 15880
rect 15940 15640 16030 15880
rect 16270 15640 16360 15880
rect 16600 15640 16690 15880
rect 16930 15640 17020 15880
rect 17260 15640 17350 15880
rect 17590 15640 17680 15880
rect 17920 15640 18010 15880
rect 18250 15640 18340 15880
rect 18580 15640 18670 15880
rect 18910 15640 19000 15880
rect 19240 15640 19330 15880
rect 19570 15640 19880 15880
rect 7640 15550 19880 15640
rect 7640 15310 7780 15550
rect 8020 15310 8110 15550
rect 8350 15310 8440 15550
rect 8680 15310 8770 15550
rect 9010 15310 9100 15550
rect 9340 15310 9430 15550
rect 9670 15310 9760 15550
rect 10000 15310 10090 15550
rect 10330 15310 10420 15550
rect 10660 15310 10750 15550
rect 10990 15310 11080 15550
rect 11320 15310 11410 15550
rect 11650 15310 11740 15550
rect 11980 15310 12070 15550
rect 12310 15310 12400 15550
rect 12640 15310 12730 15550
rect 12970 15310 13060 15550
rect 13300 15310 13390 15550
rect 13630 15310 13720 15550
rect 13960 15310 14050 15550
rect 14290 15310 14380 15550
rect 14620 15310 14710 15550
rect 14950 15310 15040 15550
rect 15280 15310 15370 15550
rect 15610 15310 15700 15550
rect 15940 15310 16030 15550
rect 16270 15310 16360 15550
rect 16600 15310 16690 15550
rect 16930 15310 17020 15550
rect 17260 15310 17350 15550
rect 17590 15310 17680 15550
rect 17920 15310 18010 15550
rect 18250 15310 18340 15550
rect 18580 15310 18670 15550
rect 18910 15310 19000 15550
rect 19240 15310 19330 15550
rect 19570 15310 19880 15550
rect 7640 15220 19880 15310
rect 7640 14980 7780 15220
rect 8020 14980 8110 15220
rect 8350 14980 8440 15220
rect 8680 14980 8770 15220
rect 9010 14980 9100 15220
rect 9340 14980 9430 15220
rect 9670 14980 9760 15220
rect 10000 14980 10090 15220
rect 10330 14980 10420 15220
rect 10660 14980 10750 15220
rect 10990 14980 11080 15220
rect 11320 14980 11410 15220
rect 11650 14980 11740 15220
rect 11980 14980 12070 15220
rect 12310 14980 12400 15220
rect 12640 14980 12730 15220
rect 12970 14980 13060 15220
rect 13300 14980 13390 15220
rect 13630 14980 13720 15220
rect 13960 14980 14050 15220
rect 14290 14980 14380 15220
rect 14620 14980 14710 15220
rect 14950 14980 15040 15220
rect 15280 14980 15370 15220
rect 15610 14980 15700 15220
rect 15940 14980 16030 15220
rect 16270 14980 16360 15220
rect 16600 14980 16690 15220
rect 16930 14980 17020 15220
rect 17260 14980 17350 15220
rect 17590 14980 17680 15220
rect 17920 14980 18010 15220
rect 18250 14980 18340 15220
rect 18580 14980 18670 15220
rect 18910 14980 19000 15220
rect 19240 14980 19330 15220
rect 19570 14980 19880 15220
rect 7640 14890 19880 14980
rect 7640 14650 7780 14890
rect 8020 14650 8110 14890
rect 8350 14650 8440 14890
rect 8680 14650 8770 14890
rect 9010 14650 9100 14890
rect 9340 14650 9430 14890
rect 9670 14650 9760 14890
rect 10000 14650 10090 14890
rect 10330 14650 10420 14890
rect 10660 14650 10750 14890
rect 10990 14650 11080 14890
rect 11320 14650 11410 14890
rect 11650 14650 11740 14890
rect 11980 14650 12070 14890
rect 12310 14650 12400 14890
rect 12640 14650 12730 14890
rect 12970 14650 13060 14890
rect 13300 14650 13390 14890
rect 13630 14650 13720 14890
rect 13960 14650 14050 14890
rect 14290 14650 14380 14890
rect 14620 14650 14710 14890
rect 14950 14650 15040 14890
rect 15280 14650 15370 14890
rect 15610 14650 15700 14890
rect 15940 14650 16030 14890
rect 16270 14650 16360 14890
rect 16600 14650 16690 14890
rect 16930 14650 17020 14890
rect 17260 14650 17350 14890
rect 17590 14650 17680 14890
rect 17920 14650 18010 14890
rect 18250 14650 18340 14890
rect 18580 14650 18670 14890
rect 18910 14650 19000 14890
rect 19240 14650 19330 14890
rect 19570 14650 19880 14890
rect 7640 14560 19880 14650
rect 7640 14320 7780 14560
rect 8020 14320 8110 14560
rect 8350 14320 8440 14560
rect 8680 14320 8770 14560
rect 9010 14320 9100 14560
rect 9340 14320 9430 14560
rect 9670 14320 9760 14560
rect 10000 14320 10090 14560
rect 10330 14320 10420 14560
rect 10660 14320 10750 14560
rect 10990 14320 11080 14560
rect 11320 14320 11410 14560
rect 11650 14320 11740 14560
rect 11980 14320 12070 14560
rect 12310 14320 12400 14560
rect 12640 14320 12730 14560
rect 12970 14320 13060 14560
rect 13300 14320 13390 14560
rect 13630 14320 13720 14560
rect 13960 14320 14050 14560
rect 14290 14320 14380 14560
rect 14620 14320 14710 14560
rect 14950 14320 15040 14560
rect 15280 14320 15370 14560
rect 15610 14320 15700 14560
rect 15940 14320 16030 14560
rect 16270 14320 16360 14560
rect 16600 14320 16690 14560
rect 16930 14320 17020 14560
rect 17260 14320 17350 14560
rect 17590 14320 17680 14560
rect 17920 14320 18010 14560
rect 18250 14320 18340 14560
rect 18580 14320 18670 14560
rect 18910 14320 19000 14560
rect 19240 14320 19330 14560
rect 19570 14320 19880 14560
rect 7640 14230 19880 14320
rect 7640 13990 7780 14230
rect 8020 13990 8110 14230
rect 8350 13990 8440 14230
rect 8680 13990 8770 14230
rect 9010 13990 9100 14230
rect 9340 13990 9430 14230
rect 9670 13990 9760 14230
rect 10000 13990 10090 14230
rect 10330 13990 10420 14230
rect 10660 13990 10750 14230
rect 10990 13990 11080 14230
rect 11320 13990 11410 14230
rect 11650 13990 11740 14230
rect 11980 13990 12070 14230
rect 12310 13990 12400 14230
rect 12640 13990 12730 14230
rect 12970 13990 13060 14230
rect 13300 13990 13390 14230
rect 13630 13990 13720 14230
rect 13960 13990 14050 14230
rect 14290 13990 14380 14230
rect 14620 13990 14710 14230
rect 14950 13990 15040 14230
rect 15280 13990 15370 14230
rect 15610 13990 15700 14230
rect 15940 13990 16030 14230
rect 16270 13990 16360 14230
rect 16600 13990 16690 14230
rect 16930 13990 17020 14230
rect 17260 13990 17350 14230
rect 17590 13990 17680 14230
rect 17920 13990 18010 14230
rect 18250 13990 18340 14230
rect 18580 13990 18670 14230
rect 18910 13990 19000 14230
rect 19240 13990 19330 14230
rect 19570 13990 19880 14230
rect 7640 13900 19880 13990
rect 7640 13660 7780 13900
rect 8020 13660 8110 13900
rect 8350 13660 8440 13900
rect 8680 13660 8770 13900
rect 9010 13660 9100 13900
rect 9340 13660 9430 13900
rect 9670 13660 9760 13900
rect 10000 13660 10090 13900
rect 10330 13660 10420 13900
rect 10660 13660 10750 13900
rect 10990 13660 11080 13900
rect 11320 13660 11410 13900
rect 11650 13660 11740 13900
rect 11980 13660 12070 13900
rect 12310 13660 12400 13900
rect 12640 13660 12730 13900
rect 12970 13660 13060 13900
rect 13300 13660 13390 13900
rect 13630 13660 13720 13900
rect 13960 13660 14050 13900
rect 14290 13660 14380 13900
rect 14620 13660 14710 13900
rect 14950 13660 15040 13900
rect 15280 13660 15370 13900
rect 15610 13660 15700 13900
rect 15940 13660 16030 13900
rect 16270 13660 16360 13900
rect 16600 13660 16690 13900
rect 16930 13660 17020 13900
rect 17260 13660 17350 13900
rect 17590 13660 17680 13900
rect 17920 13660 18010 13900
rect 18250 13660 18340 13900
rect 18580 13660 18670 13900
rect 18910 13660 19000 13900
rect 19240 13660 19330 13900
rect 19570 13660 19880 13900
rect 7640 13570 19880 13660
rect 7640 13330 7780 13570
rect 8020 13330 8110 13570
rect 8350 13330 8440 13570
rect 8680 13330 8770 13570
rect 9010 13330 9100 13570
rect 9340 13330 9430 13570
rect 9670 13330 9760 13570
rect 10000 13330 10090 13570
rect 10330 13330 10420 13570
rect 10660 13330 10750 13570
rect 10990 13330 11080 13570
rect 11320 13330 11410 13570
rect 11650 13330 11740 13570
rect 11980 13330 12070 13570
rect 12310 13330 12400 13570
rect 12640 13330 12730 13570
rect 12970 13330 13060 13570
rect 13300 13330 13390 13570
rect 13630 13330 13720 13570
rect 13960 13330 14050 13570
rect 14290 13330 14380 13570
rect 14620 13330 14710 13570
rect 14950 13330 15040 13570
rect 15280 13330 15370 13570
rect 15610 13330 15700 13570
rect 15940 13330 16030 13570
rect 16270 13330 16360 13570
rect 16600 13330 16690 13570
rect 16930 13330 17020 13570
rect 17260 13330 17350 13570
rect 17590 13330 17680 13570
rect 17920 13330 18010 13570
rect 18250 13330 18340 13570
rect 18580 13330 18670 13570
rect 18910 13330 19000 13570
rect 19240 13330 19330 13570
rect 19570 13330 19880 13570
rect 7640 13240 19880 13330
rect 7640 13000 7780 13240
rect 8020 13000 8110 13240
rect 8350 13000 8440 13240
rect 8680 13000 8770 13240
rect 9010 13000 9100 13240
rect 9340 13000 9430 13240
rect 9670 13000 9760 13240
rect 10000 13000 10090 13240
rect 10330 13000 10420 13240
rect 10660 13000 10750 13240
rect 10990 13000 11080 13240
rect 11320 13000 11410 13240
rect 11650 13000 11740 13240
rect 11980 13000 12070 13240
rect 12310 13000 12400 13240
rect 12640 13000 12730 13240
rect 12970 13000 13060 13240
rect 13300 13000 13390 13240
rect 13630 13000 13720 13240
rect 13960 13000 14050 13240
rect 14290 13000 14380 13240
rect 14620 13000 14710 13240
rect 14950 13000 15040 13240
rect 15280 13000 15370 13240
rect 15610 13000 15700 13240
rect 15940 13000 16030 13240
rect 16270 13000 16360 13240
rect 16600 13000 16690 13240
rect 16930 13000 17020 13240
rect 17260 13000 17350 13240
rect 17590 13000 17680 13240
rect 17920 13000 18010 13240
rect 18250 13000 18340 13240
rect 18580 13000 18670 13240
rect 18910 13000 19000 13240
rect 19240 13000 19330 13240
rect 19570 13000 19880 13240
rect 7640 12910 19880 13000
rect 7640 12670 7780 12910
rect 8020 12670 8110 12910
rect 8350 12670 8440 12910
rect 8680 12670 8770 12910
rect 9010 12670 9100 12910
rect 9340 12670 9430 12910
rect 9670 12670 9760 12910
rect 10000 12670 10090 12910
rect 10330 12670 10420 12910
rect 10660 12670 10750 12910
rect 10990 12670 11080 12910
rect 11320 12670 11410 12910
rect 11650 12670 11740 12910
rect 11980 12670 12070 12910
rect 12310 12670 12400 12910
rect 12640 12670 12730 12910
rect 12970 12670 13060 12910
rect 13300 12670 13390 12910
rect 13630 12670 13720 12910
rect 13960 12670 14050 12910
rect 14290 12670 14380 12910
rect 14620 12670 14710 12910
rect 14950 12670 15040 12910
rect 15280 12670 15370 12910
rect 15610 12670 15700 12910
rect 15940 12670 16030 12910
rect 16270 12670 16360 12910
rect 16600 12670 16690 12910
rect 16930 12670 17020 12910
rect 17260 12670 17350 12910
rect 17590 12670 17680 12910
rect 17920 12670 18010 12910
rect 18250 12670 18340 12910
rect 18580 12670 18670 12910
rect 18910 12670 19000 12910
rect 19240 12670 19330 12910
rect 19570 12670 19880 12910
rect 7640 12580 19880 12670
rect 7640 12340 7780 12580
rect 8020 12340 8110 12580
rect 8350 12340 8440 12580
rect 8680 12340 8770 12580
rect 9010 12340 9100 12580
rect 9340 12340 9430 12580
rect 9670 12340 9760 12580
rect 10000 12340 10090 12580
rect 10330 12340 10420 12580
rect 10660 12340 10750 12580
rect 10990 12340 11080 12580
rect 11320 12340 11410 12580
rect 11650 12340 11740 12580
rect 11980 12340 12070 12580
rect 12310 12340 12400 12580
rect 12640 12340 12730 12580
rect 12970 12340 13060 12580
rect 13300 12340 13390 12580
rect 13630 12340 13720 12580
rect 13960 12340 14050 12580
rect 14290 12340 14380 12580
rect 14620 12340 14710 12580
rect 14950 12340 15040 12580
rect 15280 12340 15370 12580
rect 15610 12340 15700 12580
rect 15940 12340 16030 12580
rect 16270 12340 16360 12580
rect 16600 12340 16690 12580
rect 16930 12340 17020 12580
rect 17260 12340 17350 12580
rect 17590 12340 17680 12580
rect 17920 12340 18010 12580
rect 18250 12340 18340 12580
rect 18580 12340 18670 12580
rect 18910 12340 19000 12580
rect 19240 12340 19330 12580
rect 19570 12340 19880 12580
rect 7640 12250 19880 12340
rect 7640 12010 7780 12250
rect 8020 12010 8110 12250
rect 8350 12010 8440 12250
rect 8680 12010 8770 12250
rect 9010 12010 9100 12250
rect 9340 12010 9430 12250
rect 9670 12010 9760 12250
rect 10000 12010 10090 12250
rect 10330 12010 10420 12250
rect 10660 12010 10750 12250
rect 10990 12010 11080 12250
rect 11320 12010 11410 12250
rect 11650 12010 11740 12250
rect 11980 12010 12070 12250
rect 12310 12010 12400 12250
rect 12640 12010 12730 12250
rect 12970 12010 13060 12250
rect 13300 12010 13390 12250
rect 13630 12010 13720 12250
rect 13960 12010 14050 12250
rect 14290 12010 14380 12250
rect 14620 12010 14710 12250
rect 14950 12010 15040 12250
rect 15280 12010 15370 12250
rect 15610 12010 15700 12250
rect 15940 12010 16030 12250
rect 16270 12010 16360 12250
rect 16600 12010 16690 12250
rect 16930 12010 17020 12250
rect 17260 12010 17350 12250
rect 17590 12010 17680 12250
rect 17920 12010 18010 12250
rect 18250 12010 18340 12250
rect 18580 12010 18670 12250
rect 18910 12010 19000 12250
rect 19240 12010 19330 12250
rect 19570 12010 19880 12250
rect 7640 11920 19880 12010
rect 7640 11680 7780 11920
rect 8020 11680 8110 11920
rect 8350 11680 8440 11920
rect 8680 11680 8770 11920
rect 9010 11680 9100 11920
rect 9340 11680 9430 11920
rect 9670 11680 9760 11920
rect 10000 11680 10090 11920
rect 10330 11680 10420 11920
rect 10660 11680 10750 11920
rect 10990 11680 11080 11920
rect 11320 11680 11410 11920
rect 11650 11680 11740 11920
rect 11980 11680 12070 11920
rect 12310 11680 12400 11920
rect 12640 11680 12730 11920
rect 12970 11680 13060 11920
rect 13300 11680 13390 11920
rect 13630 11680 13720 11920
rect 13960 11680 14050 11920
rect 14290 11680 14380 11920
rect 14620 11680 14710 11920
rect 14950 11680 15040 11920
rect 15280 11680 15370 11920
rect 15610 11680 15700 11920
rect 15940 11680 16030 11920
rect 16270 11680 16360 11920
rect 16600 11680 16690 11920
rect 16930 11680 17020 11920
rect 17260 11680 17350 11920
rect 17590 11680 17680 11920
rect 17920 11680 18010 11920
rect 18250 11680 18340 11920
rect 18580 11680 18670 11920
rect 18910 11680 19000 11920
rect 19240 11680 19330 11920
rect 19570 11680 19880 11920
rect 7640 11590 19880 11680
rect 7640 11350 7780 11590
rect 8020 11350 8110 11590
rect 8350 11350 8440 11590
rect 8680 11350 8770 11590
rect 9010 11350 9100 11590
rect 9340 11350 9430 11590
rect 9670 11350 9760 11590
rect 10000 11350 10090 11590
rect 10330 11350 10420 11590
rect 10660 11350 10750 11590
rect 10990 11350 11080 11590
rect 11320 11350 11410 11590
rect 11650 11350 11740 11590
rect 11980 11350 12070 11590
rect 12310 11350 12400 11590
rect 12640 11350 12730 11590
rect 12970 11350 13060 11590
rect 13300 11350 13390 11590
rect 13630 11350 13720 11590
rect 13960 11350 14050 11590
rect 14290 11350 14380 11590
rect 14620 11350 14710 11590
rect 14950 11350 15040 11590
rect 15280 11350 15370 11590
rect 15610 11350 15700 11590
rect 15940 11350 16030 11590
rect 16270 11350 16360 11590
rect 16600 11350 16690 11590
rect 16930 11350 17020 11590
rect 17260 11350 17350 11590
rect 17590 11350 17680 11590
rect 17920 11350 18010 11590
rect 18250 11350 18340 11590
rect 18580 11350 18670 11590
rect 18910 11350 19000 11590
rect 19240 11350 19330 11590
rect 19570 11350 19880 11590
rect 7640 11260 19880 11350
rect 7640 11020 7780 11260
rect 8020 11020 8110 11260
rect 8350 11020 8440 11260
rect 8680 11020 8770 11260
rect 9010 11020 9100 11260
rect 9340 11020 9430 11260
rect 9670 11020 9760 11260
rect 10000 11020 10090 11260
rect 10330 11020 10420 11260
rect 10660 11020 10750 11260
rect 10990 11020 11080 11260
rect 11320 11020 11410 11260
rect 11650 11020 11740 11260
rect 11980 11020 12070 11260
rect 12310 11020 12400 11260
rect 12640 11020 12730 11260
rect 12970 11020 13060 11260
rect 13300 11020 13390 11260
rect 13630 11020 13720 11260
rect 13960 11020 14050 11260
rect 14290 11020 14380 11260
rect 14620 11020 14710 11260
rect 14950 11020 15040 11260
rect 15280 11020 15370 11260
rect 15610 11020 15700 11260
rect 15940 11020 16030 11260
rect 16270 11020 16360 11260
rect 16600 11020 16690 11260
rect 16930 11020 17020 11260
rect 17260 11020 17350 11260
rect 17590 11020 17680 11260
rect 17920 11020 18010 11260
rect 18250 11020 18340 11260
rect 18580 11020 18670 11260
rect 18910 11020 19000 11260
rect 19240 11020 19330 11260
rect 19570 11020 19880 11260
rect 7640 10930 19880 11020
rect 7640 10690 7780 10930
rect 8020 10690 8110 10930
rect 8350 10690 8440 10930
rect 8680 10690 8770 10930
rect 9010 10690 9100 10930
rect 9340 10690 9430 10930
rect 9670 10690 9760 10930
rect 10000 10690 10090 10930
rect 10330 10690 10420 10930
rect 10660 10690 10750 10930
rect 10990 10690 11080 10930
rect 11320 10690 11410 10930
rect 11650 10690 11740 10930
rect 11980 10690 12070 10930
rect 12310 10690 12400 10930
rect 12640 10690 12730 10930
rect 12970 10690 13060 10930
rect 13300 10690 13390 10930
rect 13630 10690 13720 10930
rect 13960 10690 14050 10930
rect 14290 10690 14380 10930
rect 14620 10690 14710 10930
rect 14950 10690 15040 10930
rect 15280 10690 15370 10930
rect 15610 10690 15700 10930
rect 15940 10690 16030 10930
rect 16270 10690 16360 10930
rect 16600 10690 16690 10930
rect 16930 10690 17020 10930
rect 17260 10690 17350 10930
rect 17590 10690 17680 10930
rect 17920 10690 18010 10930
rect 18250 10690 18340 10930
rect 18580 10690 18670 10930
rect 18910 10690 19000 10930
rect 19240 10690 19330 10930
rect 19570 10690 19880 10930
rect 7640 10600 19880 10690
rect 7640 10360 7780 10600
rect 8020 10360 8110 10600
rect 8350 10360 8440 10600
rect 8680 10360 8770 10600
rect 9010 10360 9100 10600
rect 9340 10360 9430 10600
rect 9670 10360 9760 10600
rect 10000 10360 10090 10600
rect 10330 10360 10420 10600
rect 10660 10360 10750 10600
rect 10990 10360 11080 10600
rect 11320 10360 11410 10600
rect 11650 10360 11740 10600
rect 11980 10360 12070 10600
rect 12310 10360 12400 10600
rect 12640 10360 12730 10600
rect 12970 10360 13060 10600
rect 13300 10360 13390 10600
rect 13630 10360 13720 10600
rect 13960 10360 14050 10600
rect 14290 10360 14380 10600
rect 14620 10360 14710 10600
rect 14950 10360 15040 10600
rect 15280 10360 15370 10600
rect 15610 10360 15700 10600
rect 15940 10360 16030 10600
rect 16270 10360 16360 10600
rect 16600 10360 16690 10600
rect 16930 10360 17020 10600
rect 17260 10360 17350 10600
rect 17590 10360 17680 10600
rect 17920 10360 18010 10600
rect 18250 10360 18340 10600
rect 18580 10360 18670 10600
rect 18910 10360 19000 10600
rect 19240 10360 19330 10600
rect 19570 10360 19880 10600
rect 7640 10270 19880 10360
rect 7640 10030 7780 10270
rect 8020 10030 8110 10270
rect 8350 10030 8440 10270
rect 8680 10030 8770 10270
rect 9010 10030 9100 10270
rect 9340 10030 9430 10270
rect 9670 10030 9760 10270
rect 10000 10030 10090 10270
rect 10330 10030 10420 10270
rect 10660 10030 10750 10270
rect 10990 10030 11080 10270
rect 11320 10030 11410 10270
rect 11650 10030 11740 10270
rect 11980 10030 12070 10270
rect 12310 10030 12400 10270
rect 12640 10030 12730 10270
rect 12970 10030 13060 10270
rect 13300 10030 13390 10270
rect 13630 10030 13720 10270
rect 13960 10030 14050 10270
rect 14290 10030 14380 10270
rect 14620 10030 14710 10270
rect 14950 10030 15040 10270
rect 15280 10030 15370 10270
rect 15610 10030 15700 10270
rect 15940 10030 16030 10270
rect 16270 10030 16360 10270
rect 16600 10030 16690 10270
rect 16930 10030 17020 10270
rect 17260 10030 17350 10270
rect 17590 10030 17680 10270
rect 17920 10030 18010 10270
rect 18250 10030 18340 10270
rect 18580 10030 18670 10270
rect 18910 10030 19000 10270
rect 19240 10030 19330 10270
rect 19570 10030 19880 10270
rect 7640 9940 19880 10030
rect 7640 9700 7780 9940
rect 8020 9700 8110 9940
rect 8350 9700 8440 9940
rect 8680 9700 8770 9940
rect 9010 9700 9100 9940
rect 9340 9700 9430 9940
rect 9670 9700 9760 9940
rect 10000 9700 10090 9940
rect 10330 9700 10420 9940
rect 10660 9700 10750 9940
rect 10990 9700 11080 9940
rect 11320 9700 11410 9940
rect 11650 9700 11740 9940
rect 11980 9700 12070 9940
rect 12310 9700 12400 9940
rect 12640 9700 12730 9940
rect 12970 9700 13060 9940
rect 13300 9700 13390 9940
rect 13630 9700 13720 9940
rect 13960 9700 14050 9940
rect 14290 9700 14380 9940
rect 14620 9700 14710 9940
rect 14950 9700 15040 9940
rect 15280 9700 15370 9940
rect 15610 9700 15700 9940
rect 15940 9700 16030 9940
rect 16270 9700 16360 9940
rect 16600 9700 16690 9940
rect 16930 9700 17020 9940
rect 17260 9700 17350 9940
rect 17590 9700 17680 9940
rect 17920 9700 18010 9940
rect 18250 9700 18340 9940
rect 18580 9700 18670 9940
rect 18910 9700 19000 9940
rect 19240 9700 19330 9940
rect 19570 9700 19880 9940
rect 7640 9610 19880 9700
rect 7640 9370 7780 9610
rect 8020 9370 8110 9610
rect 8350 9370 8440 9610
rect 8680 9370 8770 9610
rect 9010 9370 9100 9610
rect 9340 9370 9430 9610
rect 9670 9370 9760 9610
rect 10000 9370 10090 9610
rect 10330 9370 10420 9610
rect 10660 9370 10750 9610
rect 10990 9370 11080 9610
rect 11320 9370 11410 9610
rect 11650 9370 11740 9610
rect 11980 9370 12070 9610
rect 12310 9370 12400 9610
rect 12640 9370 12730 9610
rect 12970 9370 13060 9610
rect 13300 9370 13390 9610
rect 13630 9370 13720 9610
rect 13960 9370 14050 9610
rect 14290 9370 14380 9610
rect 14620 9370 14710 9610
rect 14950 9370 15040 9610
rect 15280 9370 15370 9610
rect 15610 9370 15700 9610
rect 15940 9370 16030 9610
rect 16270 9370 16360 9610
rect 16600 9370 16690 9610
rect 16930 9370 17020 9610
rect 17260 9370 17350 9610
rect 17590 9370 17680 9610
rect 17920 9370 18010 9610
rect 18250 9370 18340 9610
rect 18580 9370 18670 9610
rect 18910 9370 19000 9610
rect 19240 9370 19330 9610
rect 19570 9370 19880 9610
rect 7640 9280 19880 9370
rect 7640 9040 7780 9280
rect 8020 9040 8110 9280
rect 8350 9040 8440 9280
rect 8680 9040 8770 9280
rect 9010 9040 9100 9280
rect 9340 9040 9430 9280
rect 9670 9040 9760 9280
rect 10000 9040 10090 9280
rect 10330 9040 10420 9280
rect 10660 9040 10750 9280
rect 10990 9040 11080 9280
rect 11320 9040 11410 9280
rect 11650 9040 11740 9280
rect 11980 9040 12070 9280
rect 12310 9040 12400 9280
rect 12640 9040 12730 9280
rect 12970 9040 13060 9280
rect 13300 9040 13390 9280
rect 13630 9040 13720 9280
rect 13960 9040 14050 9280
rect 14290 9040 14380 9280
rect 14620 9040 14710 9280
rect 14950 9040 15040 9280
rect 15280 9040 15370 9280
rect 15610 9040 15700 9280
rect 15940 9040 16030 9280
rect 16270 9040 16360 9280
rect 16600 9040 16690 9280
rect 16930 9040 17020 9280
rect 17260 9040 17350 9280
rect 17590 9040 17680 9280
rect 17920 9040 18010 9280
rect 18250 9040 18340 9280
rect 18580 9040 18670 9280
rect 18910 9040 19000 9280
rect 19240 9040 19330 9280
rect 19570 9040 19880 9280
rect 7640 8720 19880 9040
rect 31130 7830 37830 7880
rect 31130 7590 31180 7830
rect 31420 7590 31510 7830
rect 31750 7590 31840 7830
rect 32080 7590 32170 7830
rect 32410 7590 32500 7830
rect 32740 7590 32830 7830
rect 33070 7590 33160 7830
rect 33400 7590 33490 7830
rect 33730 7590 33820 7830
rect 34060 7590 34150 7830
rect 34390 7590 34480 7830
rect 34720 7590 34810 7830
rect 35050 7590 35140 7830
rect 35380 7590 35470 7830
rect 35710 7590 35800 7830
rect 36040 7590 36130 7830
rect 36370 7590 36460 7830
rect 36700 7590 36790 7830
rect 37030 7590 37120 7830
rect 37360 7590 37450 7830
rect 37690 7590 37830 7830
rect 31130 7500 37830 7590
rect 31130 7260 31180 7500
rect 31420 7260 31510 7500
rect 31750 7260 31840 7500
rect 32080 7260 32170 7500
rect 32410 7260 32500 7500
rect 32740 7260 32830 7500
rect 33070 7260 33160 7500
rect 33400 7260 33490 7500
rect 33730 7260 33820 7500
rect 34060 7260 34150 7500
rect 34390 7260 34480 7500
rect 34720 7260 34810 7500
rect 35050 7260 35140 7500
rect 35380 7260 35470 7500
rect 35710 7260 35800 7500
rect 36040 7260 36130 7500
rect 36370 7260 36460 7500
rect 36700 7260 36790 7500
rect 37030 7260 37120 7500
rect 37360 7260 37450 7500
rect 37690 7260 37830 7500
rect 31130 7170 37830 7260
rect 31130 6930 31180 7170
rect 31420 6930 31510 7170
rect 31750 6930 31840 7170
rect 32080 6930 32170 7170
rect 32410 6930 32500 7170
rect 32740 6930 32830 7170
rect 33070 6930 33160 7170
rect 33400 6930 33490 7170
rect 33730 6930 33820 7170
rect 34060 6930 34150 7170
rect 34390 6930 34480 7170
rect 34720 6930 34810 7170
rect 35050 6930 35140 7170
rect 35380 6930 35470 7170
rect 35710 6930 35800 7170
rect 36040 6930 36130 7170
rect 36370 6930 36460 7170
rect 36700 6930 36790 7170
rect 37030 6930 37120 7170
rect 37360 6930 37450 7170
rect 37690 6930 37830 7170
rect 31130 6840 37830 6930
rect 31130 6600 31180 6840
rect 31420 6600 31510 6840
rect 31750 6600 31840 6840
rect 32080 6600 32170 6840
rect 32410 6600 32500 6840
rect 32740 6600 32830 6840
rect 33070 6600 33160 6840
rect 33400 6600 33490 6840
rect 33730 6600 33820 6840
rect 34060 6600 34150 6840
rect 34390 6600 34480 6840
rect 34720 6600 34810 6840
rect 35050 6600 35140 6840
rect 35380 6600 35470 6840
rect 35710 6600 35800 6840
rect 36040 6600 36130 6840
rect 36370 6600 36460 6840
rect 36700 6600 36790 6840
rect 37030 6600 37120 6840
rect 37360 6600 37450 6840
rect 37690 6600 37830 6840
rect 31130 6510 37830 6600
rect 31130 6270 31180 6510
rect 31420 6270 31510 6510
rect 31750 6270 31840 6510
rect 32080 6270 32170 6510
rect 32410 6270 32500 6510
rect 32740 6270 32830 6510
rect 33070 6270 33160 6510
rect 33400 6270 33490 6510
rect 33730 6270 33820 6510
rect 34060 6270 34150 6510
rect 34390 6270 34480 6510
rect 34720 6270 34810 6510
rect 35050 6270 35140 6510
rect 35380 6270 35470 6510
rect 35710 6270 35800 6510
rect 36040 6270 36130 6510
rect 36370 6270 36460 6510
rect 36700 6270 36790 6510
rect 37030 6270 37120 6510
rect 37360 6270 37450 6510
rect 37690 6270 37830 6510
rect 31130 6180 37830 6270
rect 31130 5940 31180 6180
rect 31420 5940 31510 6180
rect 31750 5940 31840 6180
rect 32080 5940 32170 6180
rect 32410 5940 32500 6180
rect 32740 5940 32830 6180
rect 33070 5940 33160 6180
rect 33400 5940 33490 6180
rect 33730 5940 33820 6180
rect 34060 5940 34150 6180
rect 34390 5940 34480 6180
rect 34720 5940 34810 6180
rect 35050 5940 35140 6180
rect 35380 5940 35470 6180
rect 35710 5940 35800 6180
rect 36040 5940 36130 6180
rect 36370 5940 36460 6180
rect 36700 5940 36790 6180
rect 37030 5940 37120 6180
rect 37360 5940 37450 6180
rect 37690 5940 37830 6180
rect 31130 5850 37830 5940
rect 31130 5610 31180 5850
rect 31420 5610 31510 5850
rect 31750 5610 31840 5850
rect 32080 5610 32170 5850
rect 32410 5610 32500 5850
rect 32740 5610 32830 5850
rect 33070 5610 33160 5850
rect 33400 5610 33490 5850
rect 33730 5610 33820 5850
rect 34060 5610 34150 5850
rect 34390 5610 34480 5850
rect 34720 5610 34810 5850
rect 35050 5610 35140 5850
rect 35380 5610 35470 5850
rect 35710 5610 35800 5850
rect 36040 5610 36130 5850
rect 36370 5610 36460 5850
rect 36700 5610 36790 5850
rect 37030 5610 37120 5850
rect 37360 5610 37450 5850
rect 37690 5610 37830 5850
rect 31130 5520 37830 5610
rect 31130 5280 31180 5520
rect 31420 5280 31510 5520
rect 31750 5280 31840 5520
rect 32080 5280 32170 5520
rect 32410 5280 32500 5520
rect 32740 5280 32830 5520
rect 33070 5280 33160 5520
rect 33400 5280 33490 5520
rect 33730 5280 33820 5520
rect 34060 5280 34150 5520
rect 34390 5280 34480 5520
rect 34720 5280 34810 5520
rect 35050 5280 35140 5520
rect 35380 5280 35470 5520
rect 35710 5280 35800 5520
rect 36040 5280 36130 5520
rect 36370 5280 36460 5520
rect 36700 5280 36790 5520
rect 37030 5280 37120 5520
rect 37360 5280 37450 5520
rect 37690 5280 37830 5520
rect 31130 5190 37830 5280
rect 31130 4950 31180 5190
rect 31420 4950 31510 5190
rect 31750 4950 31840 5190
rect 32080 4950 32170 5190
rect 32410 4950 32500 5190
rect 32740 4950 32830 5190
rect 33070 4950 33160 5190
rect 33400 4950 33490 5190
rect 33730 4950 33820 5190
rect 34060 4950 34150 5190
rect 34390 4950 34480 5190
rect 34720 4950 34810 5190
rect 35050 4950 35140 5190
rect 35380 4950 35470 5190
rect 35710 4950 35800 5190
rect 36040 4950 36130 5190
rect 36370 4950 36460 5190
rect 36700 4950 36790 5190
rect 37030 4950 37120 5190
rect 37360 4950 37450 5190
rect 37690 4950 37830 5190
rect 31130 4860 37830 4950
rect 31130 4620 31180 4860
rect 31420 4620 31510 4860
rect 31750 4620 31840 4860
rect 32080 4620 32170 4860
rect 32410 4620 32500 4860
rect 32740 4620 32830 4860
rect 33070 4620 33160 4860
rect 33400 4620 33490 4860
rect 33730 4620 33820 4860
rect 34060 4620 34150 4860
rect 34390 4620 34480 4860
rect 34720 4620 34810 4860
rect 35050 4620 35140 4860
rect 35380 4620 35470 4860
rect 35710 4620 35800 4860
rect 36040 4620 36130 4860
rect 36370 4620 36460 4860
rect 36700 4620 36790 4860
rect 37030 4620 37120 4860
rect 37360 4620 37450 4860
rect 37690 4620 37830 4860
rect 31130 4530 37830 4620
rect 31130 4290 31180 4530
rect 31420 4290 31510 4530
rect 31750 4290 31840 4530
rect 32080 4290 32170 4530
rect 32410 4290 32500 4530
rect 32740 4290 32830 4530
rect 33070 4290 33160 4530
rect 33400 4290 33490 4530
rect 33730 4290 33820 4530
rect 34060 4290 34150 4530
rect 34390 4290 34480 4530
rect 34720 4290 34810 4530
rect 35050 4290 35140 4530
rect 35380 4290 35470 4530
rect 35710 4290 35800 4530
rect 36040 4290 36130 4530
rect 36370 4290 36460 4530
rect 36700 4290 36790 4530
rect 37030 4290 37120 4530
rect 37360 4290 37450 4530
rect 37690 4290 37830 4530
rect 31130 4200 37830 4290
rect 31130 3960 31180 4200
rect 31420 3960 31510 4200
rect 31750 3960 31840 4200
rect 32080 3960 32170 4200
rect 32410 3960 32500 4200
rect 32740 3960 32830 4200
rect 33070 3960 33160 4200
rect 33400 3960 33490 4200
rect 33730 3960 33820 4200
rect 34060 3960 34150 4200
rect 34390 3960 34480 4200
rect 34720 3960 34810 4200
rect 35050 3960 35140 4200
rect 35380 3960 35470 4200
rect 35710 3960 35800 4200
rect 36040 3960 36130 4200
rect 36370 3960 36460 4200
rect 36700 3960 36790 4200
rect 37030 3960 37120 4200
rect 37360 3960 37450 4200
rect 37690 3960 37830 4200
rect 31130 3870 37830 3960
rect 31130 3630 31180 3870
rect 31420 3630 31510 3870
rect 31750 3630 31840 3870
rect 32080 3630 32170 3870
rect 32410 3630 32500 3870
rect 32740 3630 32830 3870
rect 33070 3630 33160 3870
rect 33400 3630 33490 3870
rect 33730 3630 33820 3870
rect 34060 3630 34150 3870
rect 34390 3630 34480 3870
rect 34720 3630 34810 3870
rect 35050 3630 35140 3870
rect 35380 3630 35470 3870
rect 35710 3630 35800 3870
rect 36040 3630 36130 3870
rect 36370 3630 36460 3870
rect 36700 3630 36790 3870
rect 37030 3630 37120 3870
rect 37360 3630 37450 3870
rect 37690 3630 37830 3870
rect 31130 3540 37830 3630
rect 31130 3300 31180 3540
rect 31420 3300 31510 3540
rect 31750 3300 31840 3540
rect 32080 3300 32170 3540
rect 32410 3300 32500 3540
rect 32740 3300 32830 3540
rect 33070 3300 33160 3540
rect 33400 3300 33490 3540
rect 33730 3300 33820 3540
rect 34060 3300 34150 3540
rect 34390 3300 34480 3540
rect 34720 3300 34810 3540
rect 35050 3300 35140 3540
rect 35380 3300 35470 3540
rect 35710 3300 35800 3540
rect 36040 3300 36130 3540
rect 36370 3300 36460 3540
rect 36700 3300 36790 3540
rect 37030 3300 37120 3540
rect 37360 3300 37450 3540
rect 37690 3300 37830 3540
rect 31130 3210 37830 3300
rect 31130 2970 31180 3210
rect 31420 2970 31510 3210
rect 31750 2970 31840 3210
rect 32080 2970 32170 3210
rect 32410 2970 32500 3210
rect 32740 2970 32830 3210
rect 33070 2970 33160 3210
rect 33400 2970 33490 3210
rect 33730 2970 33820 3210
rect 34060 2970 34150 3210
rect 34390 2970 34480 3210
rect 34720 2970 34810 3210
rect 35050 2970 35140 3210
rect 35380 2970 35470 3210
rect 35710 2970 35800 3210
rect 36040 2970 36130 3210
rect 36370 2970 36460 3210
rect 36700 2970 36790 3210
rect 37030 2970 37120 3210
rect 37360 2970 37450 3210
rect 37690 2970 37830 3210
rect 31130 2880 37830 2970
rect 31130 2640 31180 2880
rect 31420 2640 31510 2880
rect 31750 2640 31840 2880
rect 32080 2640 32170 2880
rect 32410 2640 32500 2880
rect 32740 2640 32830 2880
rect 33070 2640 33160 2880
rect 33400 2640 33490 2880
rect 33730 2640 33820 2880
rect 34060 2640 34150 2880
rect 34390 2640 34480 2880
rect 34720 2640 34810 2880
rect 35050 2640 35140 2880
rect 35380 2640 35470 2880
rect 35710 2640 35800 2880
rect 36040 2640 36130 2880
rect 36370 2640 36460 2880
rect 36700 2640 36790 2880
rect 37030 2640 37120 2880
rect 37360 2640 37450 2880
rect 37690 2640 37830 2880
rect 31130 2550 37830 2640
rect 31130 2310 31180 2550
rect 31420 2310 31510 2550
rect 31750 2310 31840 2550
rect 32080 2310 32170 2550
rect 32410 2310 32500 2550
rect 32740 2310 32830 2550
rect 33070 2310 33160 2550
rect 33400 2310 33490 2550
rect 33730 2310 33820 2550
rect 34060 2310 34150 2550
rect 34390 2310 34480 2550
rect 34720 2310 34810 2550
rect 35050 2310 35140 2550
rect 35380 2310 35470 2550
rect 35710 2310 35800 2550
rect 36040 2310 36130 2550
rect 36370 2310 36460 2550
rect 36700 2310 36790 2550
rect 37030 2310 37120 2550
rect 37360 2310 37450 2550
rect 37690 2310 37830 2550
rect 31130 2220 37830 2310
rect 31130 1980 31180 2220
rect 31420 1980 31510 2220
rect 31750 1980 31840 2220
rect 32080 1980 32170 2220
rect 32410 1980 32500 2220
rect 32740 1980 32830 2220
rect 33070 1980 33160 2220
rect 33400 1980 33490 2220
rect 33730 1980 33820 2220
rect 34060 1980 34150 2220
rect 34390 1980 34480 2220
rect 34720 1980 34810 2220
rect 35050 1980 35140 2220
rect 35380 1980 35470 2220
rect 35710 1980 35800 2220
rect 36040 1980 36130 2220
rect 36370 1980 36460 2220
rect 36700 1980 36790 2220
rect 37030 1980 37120 2220
rect 37360 1980 37450 2220
rect 37690 1980 37830 2220
rect 31130 1890 37830 1980
rect 31130 1650 31180 1890
rect 31420 1650 31510 1890
rect 31750 1650 31840 1890
rect 32080 1650 32170 1890
rect 32410 1650 32500 1890
rect 32740 1650 32830 1890
rect 33070 1650 33160 1890
rect 33400 1650 33490 1890
rect 33730 1650 33820 1890
rect 34060 1650 34150 1890
rect 34390 1650 34480 1890
rect 34720 1650 34810 1890
rect 35050 1650 35140 1890
rect 35380 1650 35470 1890
rect 35710 1650 35800 1890
rect 36040 1650 36130 1890
rect 36370 1650 36460 1890
rect 36700 1650 36790 1890
rect 37030 1650 37120 1890
rect 37360 1650 37450 1890
rect 37690 1650 37830 1890
rect 31130 1560 37830 1650
rect 31130 1320 31180 1560
rect 31420 1320 31510 1560
rect 31750 1320 31840 1560
rect 32080 1320 32170 1560
rect 32410 1320 32500 1560
rect 32740 1320 32830 1560
rect 33070 1320 33160 1560
rect 33400 1320 33490 1560
rect 33730 1320 33820 1560
rect 34060 1320 34150 1560
rect 34390 1320 34480 1560
rect 34720 1320 34810 1560
rect 35050 1320 35140 1560
rect 35380 1320 35470 1560
rect 35710 1320 35800 1560
rect 36040 1320 36130 1560
rect 36370 1320 36460 1560
rect 36700 1320 36790 1560
rect 37030 1320 37120 1560
rect 37360 1320 37450 1560
rect 37690 1320 37830 1560
rect 31130 1180 37830 1320
rect 31130 230 37830 280
rect 31130 -10 31180 230
rect 31420 -10 31510 230
rect 31750 -10 31840 230
rect 32080 -10 32170 230
rect 32410 -10 32500 230
rect 32740 -10 32830 230
rect 33070 -10 33160 230
rect 33400 -10 33490 230
rect 33730 -10 33820 230
rect 34060 -10 34150 230
rect 34390 -10 34480 230
rect 34720 -10 34810 230
rect 35050 -10 35140 230
rect 35380 -10 35470 230
rect 35710 -10 35800 230
rect 36040 -10 36130 230
rect 36370 -10 36460 230
rect 36700 -10 36790 230
rect 37030 -10 37120 230
rect 37360 -10 37450 230
rect 37690 -10 37830 230
rect 31130 -100 37830 -10
rect 31130 -340 31180 -100
rect 31420 -340 31510 -100
rect 31750 -340 31840 -100
rect 32080 -340 32170 -100
rect 32410 -340 32500 -100
rect 32740 -340 32830 -100
rect 33070 -340 33160 -100
rect 33400 -340 33490 -100
rect 33730 -340 33820 -100
rect 34060 -340 34150 -100
rect 34390 -340 34480 -100
rect 34720 -340 34810 -100
rect 35050 -340 35140 -100
rect 35380 -340 35470 -100
rect 35710 -340 35800 -100
rect 36040 -340 36130 -100
rect 36370 -340 36460 -100
rect 36700 -340 36790 -100
rect 37030 -340 37120 -100
rect 37360 -340 37450 -100
rect 37690 -340 37830 -100
rect 31130 -430 37830 -340
rect 31130 -670 31180 -430
rect 31420 -670 31510 -430
rect 31750 -670 31840 -430
rect 32080 -670 32170 -430
rect 32410 -670 32500 -430
rect 32740 -670 32830 -430
rect 33070 -670 33160 -430
rect 33400 -670 33490 -430
rect 33730 -670 33820 -430
rect 34060 -670 34150 -430
rect 34390 -670 34480 -430
rect 34720 -670 34810 -430
rect 35050 -670 35140 -430
rect 35380 -670 35470 -430
rect 35710 -670 35800 -430
rect 36040 -670 36130 -430
rect 36370 -670 36460 -430
rect 36700 -670 36790 -430
rect 37030 -670 37120 -430
rect 37360 -670 37450 -430
rect 37690 -670 37830 -430
rect 31130 -760 37830 -670
rect 31130 -1000 31180 -760
rect 31420 -1000 31510 -760
rect 31750 -1000 31840 -760
rect 32080 -1000 32170 -760
rect 32410 -1000 32500 -760
rect 32740 -1000 32830 -760
rect 33070 -1000 33160 -760
rect 33400 -1000 33490 -760
rect 33730 -1000 33820 -760
rect 34060 -1000 34150 -760
rect 34390 -1000 34480 -760
rect 34720 -1000 34810 -760
rect 35050 -1000 35140 -760
rect 35380 -1000 35470 -760
rect 35710 -1000 35800 -760
rect 36040 -1000 36130 -760
rect 36370 -1000 36460 -760
rect 36700 -1000 36790 -760
rect 37030 -1000 37120 -760
rect 37360 -1000 37450 -760
rect 37690 -1000 37830 -760
rect 31130 -1090 37830 -1000
rect 31130 -1330 31180 -1090
rect 31420 -1330 31510 -1090
rect 31750 -1330 31840 -1090
rect 32080 -1330 32170 -1090
rect 32410 -1330 32500 -1090
rect 32740 -1330 32830 -1090
rect 33070 -1330 33160 -1090
rect 33400 -1330 33490 -1090
rect 33730 -1330 33820 -1090
rect 34060 -1330 34150 -1090
rect 34390 -1330 34480 -1090
rect 34720 -1330 34810 -1090
rect 35050 -1330 35140 -1090
rect 35380 -1330 35470 -1090
rect 35710 -1330 35800 -1090
rect 36040 -1330 36130 -1090
rect 36370 -1330 36460 -1090
rect 36700 -1330 36790 -1090
rect 37030 -1330 37120 -1090
rect 37360 -1330 37450 -1090
rect 37690 -1330 37830 -1090
rect 31130 -1420 37830 -1330
rect 31130 -1660 31180 -1420
rect 31420 -1660 31510 -1420
rect 31750 -1660 31840 -1420
rect 32080 -1660 32170 -1420
rect 32410 -1660 32500 -1420
rect 32740 -1660 32830 -1420
rect 33070 -1660 33160 -1420
rect 33400 -1660 33490 -1420
rect 33730 -1660 33820 -1420
rect 34060 -1660 34150 -1420
rect 34390 -1660 34480 -1420
rect 34720 -1660 34810 -1420
rect 35050 -1660 35140 -1420
rect 35380 -1660 35470 -1420
rect 35710 -1660 35800 -1420
rect 36040 -1660 36130 -1420
rect 36370 -1660 36460 -1420
rect 36700 -1660 36790 -1420
rect 37030 -1660 37120 -1420
rect 37360 -1660 37450 -1420
rect 37690 -1660 37830 -1420
rect 31130 -1750 37830 -1660
rect 31130 -1990 31180 -1750
rect 31420 -1990 31510 -1750
rect 31750 -1990 31840 -1750
rect 32080 -1990 32170 -1750
rect 32410 -1990 32500 -1750
rect 32740 -1990 32830 -1750
rect 33070 -1990 33160 -1750
rect 33400 -1990 33490 -1750
rect 33730 -1990 33820 -1750
rect 34060 -1990 34150 -1750
rect 34390 -1990 34480 -1750
rect 34720 -1990 34810 -1750
rect 35050 -1990 35140 -1750
rect 35380 -1990 35470 -1750
rect 35710 -1990 35800 -1750
rect 36040 -1990 36130 -1750
rect 36370 -1990 36460 -1750
rect 36700 -1990 36790 -1750
rect 37030 -1990 37120 -1750
rect 37360 -1990 37450 -1750
rect 37690 -1990 37830 -1750
rect 31130 -2080 37830 -1990
rect 31130 -2320 31180 -2080
rect 31420 -2320 31510 -2080
rect 31750 -2320 31840 -2080
rect 32080 -2320 32170 -2080
rect 32410 -2320 32500 -2080
rect 32740 -2320 32830 -2080
rect 33070 -2320 33160 -2080
rect 33400 -2320 33490 -2080
rect 33730 -2320 33820 -2080
rect 34060 -2320 34150 -2080
rect 34390 -2320 34480 -2080
rect 34720 -2320 34810 -2080
rect 35050 -2320 35140 -2080
rect 35380 -2320 35470 -2080
rect 35710 -2320 35800 -2080
rect 36040 -2320 36130 -2080
rect 36370 -2320 36460 -2080
rect 36700 -2320 36790 -2080
rect 37030 -2320 37120 -2080
rect 37360 -2320 37450 -2080
rect 37690 -2320 37830 -2080
rect 31130 -2410 37830 -2320
rect 31130 -2650 31180 -2410
rect 31420 -2650 31510 -2410
rect 31750 -2650 31840 -2410
rect 32080 -2650 32170 -2410
rect 32410 -2650 32500 -2410
rect 32740 -2650 32830 -2410
rect 33070 -2650 33160 -2410
rect 33400 -2650 33490 -2410
rect 33730 -2650 33820 -2410
rect 34060 -2650 34150 -2410
rect 34390 -2650 34480 -2410
rect 34720 -2650 34810 -2410
rect 35050 -2650 35140 -2410
rect 35380 -2650 35470 -2410
rect 35710 -2650 35800 -2410
rect 36040 -2650 36130 -2410
rect 36370 -2650 36460 -2410
rect 36700 -2650 36790 -2410
rect 37030 -2650 37120 -2410
rect 37360 -2650 37450 -2410
rect 37690 -2650 37830 -2410
rect 31130 -2740 37830 -2650
rect 31130 -2980 31180 -2740
rect 31420 -2980 31510 -2740
rect 31750 -2980 31840 -2740
rect 32080 -2980 32170 -2740
rect 32410 -2980 32500 -2740
rect 32740 -2980 32830 -2740
rect 33070 -2980 33160 -2740
rect 33400 -2980 33490 -2740
rect 33730 -2980 33820 -2740
rect 34060 -2980 34150 -2740
rect 34390 -2980 34480 -2740
rect 34720 -2980 34810 -2740
rect 35050 -2980 35140 -2740
rect 35380 -2980 35470 -2740
rect 35710 -2980 35800 -2740
rect 36040 -2980 36130 -2740
rect 36370 -2980 36460 -2740
rect 36700 -2980 36790 -2740
rect 37030 -2980 37120 -2740
rect 37360 -2980 37450 -2740
rect 37690 -2980 37830 -2740
rect 31130 -3070 37830 -2980
rect 31130 -3310 31180 -3070
rect 31420 -3310 31510 -3070
rect 31750 -3310 31840 -3070
rect 32080 -3310 32170 -3070
rect 32410 -3310 32500 -3070
rect 32740 -3310 32830 -3070
rect 33070 -3310 33160 -3070
rect 33400 -3310 33490 -3070
rect 33730 -3310 33820 -3070
rect 34060 -3310 34150 -3070
rect 34390 -3310 34480 -3070
rect 34720 -3310 34810 -3070
rect 35050 -3310 35140 -3070
rect 35380 -3310 35470 -3070
rect 35710 -3310 35800 -3070
rect 36040 -3310 36130 -3070
rect 36370 -3310 36460 -3070
rect 36700 -3310 36790 -3070
rect 37030 -3310 37120 -3070
rect 37360 -3310 37450 -3070
rect 37690 -3310 37830 -3070
rect 31130 -3400 37830 -3310
rect 31130 -3640 31180 -3400
rect 31420 -3640 31510 -3400
rect 31750 -3640 31840 -3400
rect 32080 -3640 32170 -3400
rect 32410 -3640 32500 -3400
rect 32740 -3640 32830 -3400
rect 33070 -3640 33160 -3400
rect 33400 -3640 33490 -3400
rect 33730 -3640 33820 -3400
rect 34060 -3640 34150 -3400
rect 34390 -3640 34480 -3400
rect 34720 -3640 34810 -3400
rect 35050 -3640 35140 -3400
rect 35380 -3640 35470 -3400
rect 35710 -3640 35800 -3400
rect 36040 -3640 36130 -3400
rect 36370 -3640 36460 -3400
rect 36700 -3640 36790 -3400
rect 37030 -3640 37120 -3400
rect 37360 -3640 37450 -3400
rect 37690 -3640 37830 -3400
rect 31130 -3730 37830 -3640
rect 31130 -3970 31180 -3730
rect 31420 -3970 31510 -3730
rect 31750 -3970 31840 -3730
rect 32080 -3970 32170 -3730
rect 32410 -3970 32500 -3730
rect 32740 -3970 32830 -3730
rect 33070 -3970 33160 -3730
rect 33400 -3970 33490 -3730
rect 33730 -3970 33820 -3730
rect 34060 -3970 34150 -3730
rect 34390 -3970 34480 -3730
rect 34720 -3970 34810 -3730
rect 35050 -3970 35140 -3730
rect 35380 -3970 35470 -3730
rect 35710 -3970 35800 -3730
rect 36040 -3970 36130 -3730
rect 36370 -3970 36460 -3730
rect 36700 -3970 36790 -3730
rect 37030 -3970 37120 -3730
rect 37360 -3970 37450 -3730
rect 37690 -3970 37830 -3730
rect 31130 -4060 37830 -3970
rect 31130 -4300 31180 -4060
rect 31420 -4300 31510 -4060
rect 31750 -4300 31840 -4060
rect 32080 -4300 32170 -4060
rect 32410 -4300 32500 -4060
rect 32740 -4300 32830 -4060
rect 33070 -4300 33160 -4060
rect 33400 -4300 33490 -4060
rect 33730 -4300 33820 -4060
rect 34060 -4300 34150 -4060
rect 34390 -4300 34480 -4060
rect 34720 -4300 34810 -4060
rect 35050 -4300 35140 -4060
rect 35380 -4300 35470 -4060
rect 35710 -4300 35800 -4060
rect 36040 -4300 36130 -4060
rect 36370 -4300 36460 -4060
rect 36700 -4300 36790 -4060
rect 37030 -4300 37120 -4060
rect 37360 -4300 37450 -4060
rect 37690 -4300 37830 -4060
rect 31130 -4390 37830 -4300
rect 31130 -4630 31180 -4390
rect 31420 -4630 31510 -4390
rect 31750 -4630 31840 -4390
rect 32080 -4630 32170 -4390
rect 32410 -4630 32500 -4390
rect 32740 -4630 32830 -4390
rect 33070 -4630 33160 -4390
rect 33400 -4630 33490 -4390
rect 33730 -4630 33820 -4390
rect 34060 -4630 34150 -4390
rect 34390 -4630 34480 -4390
rect 34720 -4630 34810 -4390
rect 35050 -4630 35140 -4390
rect 35380 -4630 35470 -4390
rect 35710 -4630 35800 -4390
rect 36040 -4630 36130 -4390
rect 36370 -4630 36460 -4390
rect 36700 -4630 36790 -4390
rect 37030 -4630 37120 -4390
rect 37360 -4630 37450 -4390
rect 37690 -4630 37830 -4390
rect -1320 -4840 230 -4660
rect -1320 -5080 -1180 -4840
rect -940 -5080 -850 -4840
rect -610 -5080 -520 -4840
rect -280 -5080 -190 -4840
rect 50 -5080 230 -4840
rect -1320 -5170 230 -5080
rect -1320 -5410 -1180 -5170
rect -940 -5410 -850 -5170
rect -610 -5410 -520 -5170
rect -280 -5410 -190 -5170
rect 50 -5410 230 -5170
rect -1320 -5500 230 -5410
rect -1320 -5740 -1180 -5500
rect -940 -5740 -850 -5500
rect -610 -5740 -520 -5500
rect -280 -5740 -190 -5500
rect 50 -5740 230 -5500
rect -1320 -5830 230 -5740
rect -1320 -6070 -1180 -5830
rect -940 -6070 -850 -5830
rect -610 -6070 -520 -5830
rect -280 -6070 -190 -5830
rect 50 -6070 230 -5830
rect -1320 -6210 230 -6070
rect 14550 -4840 16100 -4660
rect 14550 -5080 14730 -4840
rect 14970 -5080 15060 -4840
rect 15300 -5080 15390 -4840
rect 15630 -5080 15720 -4840
rect 15960 -5080 16100 -4840
rect 14550 -5170 16100 -5080
rect 14550 -5410 14730 -5170
rect 14970 -5410 15060 -5170
rect 15300 -5410 15390 -5170
rect 15630 -5410 15720 -5170
rect 15960 -5410 16100 -5170
rect 14550 -5500 16100 -5410
rect 14550 -5740 14730 -5500
rect 14970 -5740 15060 -5500
rect 15300 -5740 15390 -5500
rect 15630 -5740 15720 -5500
rect 15960 -5740 16100 -5500
rect 14550 -5830 16100 -5740
rect 14550 -6070 14730 -5830
rect 14970 -6070 15060 -5830
rect 15300 -6070 15390 -5830
rect 15630 -6070 15720 -5830
rect 15960 -6070 16100 -5830
rect 14550 -6210 16100 -6070
rect 31130 -4720 37830 -4630
rect 31130 -4960 31180 -4720
rect 31420 -4960 31510 -4720
rect 31750 -4960 31840 -4720
rect 32080 -4960 32170 -4720
rect 32410 -4960 32500 -4720
rect 32740 -4960 32830 -4720
rect 33070 -4960 33160 -4720
rect 33400 -4960 33490 -4720
rect 33730 -4960 33820 -4720
rect 34060 -4960 34150 -4720
rect 34390 -4960 34480 -4720
rect 34720 -4960 34810 -4720
rect 35050 -4960 35140 -4720
rect 35380 -4960 35470 -4720
rect 35710 -4960 35800 -4720
rect 36040 -4960 36130 -4720
rect 36370 -4960 36460 -4720
rect 36700 -4960 36790 -4720
rect 37030 -4960 37120 -4720
rect 37360 -4960 37450 -4720
rect 37690 -4960 37830 -4720
rect 31130 -5050 37830 -4960
rect 31130 -5290 31180 -5050
rect 31420 -5290 31510 -5050
rect 31750 -5290 31840 -5050
rect 32080 -5290 32170 -5050
rect 32410 -5290 32500 -5050
rect 32740 -5290 32830 -5050
rect 33070 -5290 33160 -5050
rect 33400 -5290 33490 -5050
rect 33730 -5290 33820 -5050
rect 34060 -5290 34150 -5050
rect 34390 -5290 34480 -5050
rect 34720 -5290 34810 -5050
rect 35050 -5290 35140 -5050
rect 35380 -5290 35470 -5050
rect 35710 -5290 35800 -5050
rect 36040 -5290 36130 -5050
rect 36370 -5290 36460 -5050
rect 36700 -5290 36790 -5050
rect 37030 -5290 37120 -5050
rect 37360 -5290 37450 -5050
rect 37690 -5290 37830 -5050
rect 31130 -5380 37830 -5290
rect 31130 -5620 31180 -5380
rect 31420 -5620 31510 -5380
rect 31750 -5620 31840 -5380
rect 32080 -5620 32170 -5380
rect 32410 -5620 32500 -5380
rect 32740 -5620 32830 -5380
rect 33070 -5620 33160 -5380
rect 33400 -5620 33490 -5380
rect 33730 -5620 33820 -5380
rect 34060 -5620 34150 -5380
rect 34390 -5620 34480 -5380
rect 34720 -5620 34810 -5380
rect 35050 -5620 35140 -5380
rect 35380 -5620 35470 -5380
rect 35710 -5620 35800 -5380
rect 36040 -5620 36130 -5380
rect 36370 -5620 36460 -5380
rect 36700 -5620 36790 -5380
rect 37030 -5620 37120 -5380
rect 37360 -5620 37450 -5380
rect 37690 -5620 37830 -5380
rect 31130 -5710 37830 -5620
rect 31130 -5950 31180 -5710
rect 31420 -5950 31510 -5710
rect 31750 -5950 31840 -5710
rect 32080 -5950 32170 -5710
rect 32410 -5950 32500 -5710
rect 32740 -5950 32830 -5710
rect 33070 -5950 33160 -5710
rect 33400 -5950 33490 -5710
rect 33730 -5950 33820 -5710
rect 34060 -5950 34150 -5710
rect 34390 -5950 34480 -5710
rect 34720 -5950 34810 -5710
rect 35050 -5950 35140 -5710
rect 35380 -5950 35470 -5710
rect 35710 -5950 35800 -5710
rect 36040 -5950 36130 -5710
rect 36370 -5950 36460 -5710
rect 36700 -5950 36790 -5710
rect 37030 -5950 37120 -5710
rect 37360 -5950 37450 -5710
rect 37690 -5950 37830 -5710
rect 31130 -6040 37830 -5950
rect 31130 -6280 31180 -6040
rect 31420 -6280 31510 -6040
rect 31750 -6280 31840 -6040
rect 32080 -6280 32170 -6040
rect 32410 -6280 32500 -6040
rect 32740 -6280 32830 -6040
rect 33070 -6280 33160 -6040
rect 33400 -6280 33490 -6040
rect 33730 -6280 33820 -6040
rect 34060 -6280 34150 -6040
rect 34390 -6280 34480 -6040
rect 34720 -6280 34810 -6040
rect 35050 -6280 35140 -6040
rect 35380 -6280 35470 -6040
rect 35710 -6280 35800 -6040
rect 36040 -6280 36130 -6040
rect 36370 -6280 36460 -6040
rect 36700 -6280 36790 -6040
rect 37030 -6280 37120 -6040
rect 37360 -6280 37450 -6040
rect 37690 -6280 37830 -6040
rect 31130 -6420 37830 -6280
<< mimcapcontact >>
rect -4670 20590 -4430 20830
rect -4340 20590 -4100 20830
rect -4010 20590 -3770 20830
rect -3680 20590 -3440 20830
rect -3350 20590 -3110 20830
rect -3020 20590 -2780 20830
rect -2690 20590 -2450 20830
rect -2360 20590 -2120 20830
rect -2030 20590 -1790 20830
rect -1700 20590 -1460 20830
rect -1370 20590 -1130 20830
rect -1040 20590 -800 20830
rect -710 20590 -470 20830
rect -380 20590 -140 20830
rect -50 20590 190 20830
rect 280 20590 520 20830
rect 610 20590 850 20830
rect 940 20590 1180 20830
rect 1270 20590 1510 20830
rect 1600 20590 1840 20830
rect 1930 20590 2170 20830
rect 2260 20590 2500 20830
rect 2590 20590 2830 20830
rect 2920 20590 3160 20830
rect 3250 20590 3490 20830
rect 3580 20590 3820 20830
rect 3910 20590 4150 20830
rect 4240 20590 4480 20830
rect 4570 20590 4810 20830
rect 4900 20590 5140 20830
rect 5230 20590 5470 20830
rect 5560 20590 5800 20830
rect 5890 20590 6130 20830
rect 6220 20590 6460 20830
rect 6550 20590 6790 20830
rect 6880 20590 7120 20830
rect -4670 20260 -4430 20500
rect -4340 20260 -4100 20500
rect -4010 20260 -3770 20500
rect -3680 20260 -3440 20500
rect -3350 20260 -3110 20500
rect -3020 20260 -2780 20500
rect -2690 20260 -2450 20500
rect -2360 20260 -2120 20500
rect -2030 20260 -1790 20500
rect -1700 20260 -1460 20500
rect -1370 20260 -1130 20500
rect -1040 20260 -800 20500
rect -710 20260 -470 20500
rect -380 20260 -140 20500
rect -50 20260 190 20500
rect 280 20260 520 20500
rect 610 20260 850 20500
rect 940 20260 1180 20500
rect 1270 20260 1510 20500
rect 1600 20260 1840 20500
rect 1930 20260 2170 20500
rect 2260 20260 2500 20500
rect 2590 20260 2830 20500
rect 2920 20260 3160 20500
rect 3250 20260 3490 20500
rect 3580 20260 3820 20500
rect 3910 20260 4150 20500
rect 4240 20260 4480 20500
rect 4570 20260 4810 20500
rect 4900 20260 5140 20500
rect 5230 20260 5470 20500
rect 5560 20260 5800 20500
rect 5890 20260 6130 20500
rect 6220 20260 6460 20500
rect 6550 20260 6790 20500
rect 6880 20260 7120 20500
rect -4670 19930 -4430 20170
rect -4340 19930 -4100 20170
rect -4010 19930 -3770 20170
rect -3680 19930 -3440 20170
rect -3350 19930 -3110 20170
rect -3020 19930 -2780 20170
rect -2690 19930 -2450 20170
rect -2360 19930 -2120 20170
rect -2030 19930 -1790 20170
rect -1700 19930 -1460 20170
rect -1370 19930 -1130 20170
rect -1040 19930 -800 20170
rect -710 19930 -470 20170
rect -380 19930 -140 20170
rect -50 19930 190 20170
rect 280 19930 520 20170
rect 610 19930 850 20170
rect 940 19930 1180 20170
rect 1270 19930 1510 20170
rect 1600 19930 1840 20170
rect 1930 19930 2170 20170
rect 2260 19930 2500 20170
rect 2590 19930 2830 20170
rect 2920 19930 3160 20170
rect 3250 19930 3490 20170
rect 3580 19930 3820 20170
rect 3910 19930 4150 20170
rect 4240 19930 4480 20170
rect 4570 19930 4810 20170
rect 4900 19930 5140 20170
rect 5230 19930 5470 20170
rect 5560 19930 5800 20170
rect 5890 19930 6130 20170
rect 6220 19930 6460 20170
rect 6550 19930 6790 20170
rect 6880 19930 7120 20170
rect -4670 19600 -4430 19840
rect -4340 19600 -4100 19840
rect -4010 19600 -3770 19840
rect -3680 19600 -3440 19840
rect -3350 19600 -3110 19840
rect -3020 19600 -2780 19840
rect -2690 19600 -2450 19840
rect -2360 19600 -2120 19840
rect -2030 19600 -1790 19840
rect -1700 19600 -1460 19840
rect -1370 19600 -1130 19840
rect -1040 19600 -800 19840
rect -710 19600 -470 19840
rect -380 19600 -140 19840
rect -50 19600 190 19840
rect 280 19600 520 19840
rect 610 19600 850 19840
rect 940 19600 1180 19840
rect 1270 19600 1510 19840
rect 1600 19600 1840 19840
rect 1930 19600 2170 19840
rect 2260 19600 2500 19840
rect 2590 19600 2830 19840
rect 2920 19600 3160 19840
rect 3250 19600 3490 19840
rect 3580 19600 3820 19840
rect 3910 19600 4150 19840
rect 4240 19600 4480 19840
rect 4570 19600 4810 19840
rect 4900 19600 5140 19840
rect 5230 19600 5470 19840
rect 5560 19600 5800 19840
rect 5890 19600 6130 19840
rect 6220 19600 6460 19840
rect 6550 19600 6790 19840
rect 6880 19600 7120 19840
rect -4670 19270 -4430 19510
rect -4340 19270 -4100 19510
rect -4010 19270 -3770 19510
rect -3680 19270 -3440 19510
rect -3350 19270 -3110 19510
rect -3020 19270 -2780 19510
rect -2690 19270 -2450 19510
rect -2360 19270 -2120 19510
rect -2030 19270 -1790 19510
rect -1700 19270 -1460 19510
rect -1370 19270 -1130 19510
rect -1040 19270 -800 19510
rect -710 19270 -470 19510
rect -380 19270 -140 19510
rect -50 19270 190 19510
rect 280 19270 520 19510
rect 610 19270 850 19510
rect 940 19270 1180 19510
rect 1270 19270 1510 19510
rect 1600 19270 1840 19510
rect 1930 19270 2170 19510
rect 2260 19270 2500 19510
rect 2590 19270 2830 19510
rect 2920 19270 3160 19510
rect 3250 19270 3490 19510
rect 3580 19270 3820 19510
rect 3910 19270 4150 19510
rect 4240 19270 4480 19510
rect 4570 19270 4810 19510
rect 4900 19270 5140 19510
rect 5230 19270 5470 19510
rect 5560 19270 5800 19510
rect 5890 19270 6130 19510
rect 6220 19270 6460 19510
rect 6550 19270 6790 19510
rect 6880 19270 7120 19510
rect -4670 18940 -4430 19180
rect -4340 18940 -4100 19180
rect -4010 18940 -3770 19180
rect -3680 18940 -3440 19180
rect -3350 18940 -3110 19180
rect -3020 18940 -2780 19180
rect -2690 18940 -2450 19180
rect -2360 18940 -2120 19180
rect -2030 18940 -1790 19180
rect -1700 18940 -1460 19180
rect -1370 18940 -1130 19180
rect -1040 18940 -800 19180
rect -710 18940 -470 19180
rect -380 18940 -140 19180
rect -50 18940 190 19180
rect 280 18940 520 19180
rect 610 18940 850 19180
rect 940 18940 1180 19180
rect 1270 18940 1510 19180
rect 1600 18940 1840 19180
rect 1930 18940 2170 19180
rect 2260 18940 2500 19180
rect 2590 18940 2830 19180
rect 2920 18940 3160 19180
rect 3250 18940 3490 19180
rect 3580 18940 3820 19180
rect 3910 18940 4150 19180
rect 4240 18940 4480 19180
rect 4570 18940 4810 19180
rect 4900 18940 5140 19180
rect 5230 18940 5470 19180
rect 5560 18940 5800 19180
rect 5890 18940 6130 19180
rect 6220 18940 6460 19180
rect 6550 18940 6790 19180
rect 6880 18940 7120 19180
rect -4670 18610 -4430 18850
rect -4340 18610 -4100 18850
rect -4010 18610 -3770 18850
rect -3680 18610 -3440 18850
rect -3350 18610 -3110 18850
rect -3020 18610 -2780 18850
rect -2690 18610 -2450 18850
rect -2360 18610 -2120 18850
rect -2030 18610 -1790 18850
rect -1700 18610 -1460 18850
rect -1370 18610 -1130 18850
rect -1040 18610 -800 18850
rect -710 18610 -470 18850
rect -380 18610 -140 18850
rect -50 18610 190 18850
rect 280 18610 520 18850
rect 610 18610 850 18850
rect 940 18610 1180 18850
rect 1270 18610 1510 18850
rect 1600 18610 1840 18850
rect 1930 18610 2170 18850
rect 2260 18610 2500 18850
rect 2590 18610 2830 18850
rect 2920 18610 3160 18850
rect 3250 18610 3490 18850
rect 3580 18610 3820 18850
rect 3910 18610 4150 18850
rect 4240 18610 4480 18850
rect 4570 18610 4810 18850
rect 4900 18610 5140 18850
rect 5230 18610 5470 18850
rect 5560 18610 5800 18850
rect 5890 18610 6130 18850
rect 6220 18610 6460 18850
rect 6550 18610 6790 18850
rect 6880 18610 7120 18850
rect -4670 18280 -4430 18520
rect -4340 18280 -4100 18520
rect -4010 18280 -3770 18520
rect -3680 18280 -3440 18520
rect -3350 18280 -3110 18520
rect -3020 18280 -2780 18520
rect -2690 18280 -2450 18520
rect -2360 18280 -2120 18520
rect -2030 18280 -1790 18520
rect -1700 18280 -1460 18520
rect -1370 18280 -1130 18520
rect -1040 18280 -800 18520
rect -710 18280 -470 18520
rect -380 18280 -140 18520
rect -50 18280 190 18520
rect 280 18280 520 18520
rect 610 18280 850 18520
rect 940 18280 1180 18520
rect 1270 18280 1510 18520
rect 1600 18280 1840 18520
rect 1930 18280 2170 18520
rect 2260 18280 2500 18520
rect 2590 18280 2830 18520
rect 2920 18280 3160 18520
rect 3250 18280 3490 18520
rect 3580 18280 3820 18520
rect 3910 18280 4150 18520
rect 4240 18280 4480 18520
rect 4570 18280 4810 18520
rect 4900 18280 5140 18520
rect 5230 18280 5470 18520
rect 5560 18280 5800 18520
rect 5890 18280 6130 18520
rect 6220 18280 6460 18520
rect 6550 18280 6790 18520
rect 6880 18280 7120 18520
rect -4670 17950 -4430 18190
rect -4340 17950 -4100 18190
rect -4010 17950 -3770 18190
rect -3680 17950 -3440 18190
rect -3350 17950 -3110 18190
rect -3020 17950 -2780 18190
rect -2690 17950 -2450 18190
rect -2360 17950 -2120 18190
rect -2030 17950 -1790 18190
rect -1700 17950 -1460 18190
rect -1370 17950 -1130 18190
rect -1040 17950 -800 18190
rect -710 17950 -470 18190
rect -380 17950 -140 18190
rect -50 17950 190 18190
rect 280 17950 520 18190
rect 610 17950 850 18190
rect 940 17950 1180 18190
rect 1270 17950 1510 18190
rect 1600 17950 1840 18190
rect 1930 17950 2170 18190
rect 2260 17950 2500 18190
rect 2590 17950 2830 18190
rect 2920 17950 3160 18190
rect 3250 17950 3490 18190
rect 3580 17950 3820 18190
rect 3910 17950 4150 18190
rect 4240 17950 4480 18190
rect 4570 17950 4810 18190
rect 4900 17950 5140 18190
rect 5230 17950 5470 18190
rect 5560 17950 5800 18190
rect 5890 17950 6130 18190
rect 6220 17950 6460 18190
rect 6550 17950 6790 18190
rect 6880 17950 7120 18190
rect -4670 17620 -4430 17860
rect -4340 17620 -4100 17860
rect -4010 17620 -3770 17860
rect -3680 17620 -3440 17860
rect -3350 17620 -3110 17860
rect -3020 17620 -2780 17860
rect -2690 17620 -2450 17860
rect -2360 17620 -2120 17860
rect -2030 17620 -1790 17860
rect -1700 17620 -1460 17860
rect -1370 17620 -1130 17860
rect -1040 17620 -800 17860
rect -710 17620 -470 17860
rect -380 17620 -140 17860
rect -50 17620 190 17860
rect 280 17620 520 17860
rect 610 17620 850 17860
rect 940 17620 1180 17860
rect 1270 17620 1510 17860
rect 1600 17620 1840 17860
rect 1930 17620 2170 17860
rect 2260 17620 2500 17860
rect 2590 17620 2830 17860
rect 2920 17620 3160 17860
rect 3250 17620 3490 17860
rect 3580 17620 3820 17860
rect 3910 17620 4150 17860
rect 4240 17620 4480 17860
rect 4570 17620 4810 17860
rect 4900 17620 5140 17860
rect 5230 17620 5470 17860
rect 5560 17620 5800 17860
rect 5890 17620 6130 17860
rect 6220 17620 6460 17860
rect 6550 17620 6790 17860
rect 6880 17620 7120 17860
rect -4670 17290 -4430 17530
rect -4340 17290 -4100 17530
rect -4010 17290 -3770 17530
rect -3680 17290 -3440 17530
rect -3350 17290 -3110 17530
rect -3020 17290 -2780 17530
rect -2690 17290 -2450 17530
rect -2360 17290 -2120 17530
rect -2030 17290 -1790 17530
rect -1700 17290 -1460 17530
rect -1370 17290 -1130 17530
rect -1040 17290 -800 17530
rect -710 17290 -470 17530
rect -380 17290 -140 17530
rect -50 17290 190 17530
rect 280 17290 520 17530
rect 610 17290 850 17530
rect 940 17290 1180 17530
rect 1270 17290 1510 17530
rect 1600 17290 1840 17530
rect 1930 17290 2170 17530
rect 2260 17290 2500 17530
rect 2590 17290 2830 17530
rect 2920 17290 3160 17530
rect 3250 17290 3490 17530
rect 3580 17290 3820 17530
rect 3910 17290 4150 17530
rect 4240 17290 4480 17530
rect 4570 17290 4810 17530
rect 4900 17290 5140 17530
rect 5230 17290 5470 17530
rect 5560 17290 5800 17530
rect 5890 17290 6130 17530
rect 6220 17290 6460 17530
rect 6550 17290 6790 17530
rect 6880 17290 7120 17530
rect -4670 16960 -4430 17200
rect -4340 16960 -4100 17200
rect -4010 16960 -3770 17200
rect -3680 16960 -3440 17200
rect -3350 16960 -3110 17200
rect -3020 16960 -2780 17200
rect -2690 16960 -2450 17200
rect -2360 16960 -2120 17200
rect -2030 16960 -1790 17200
rect -1700 16960 -1460 17200
rect -1370 16960 -1130 17200
rect -1040 16960 -800 17200
rect -710 16960 -470 17200
rect -380 16960 -140 17200
rect -50 16960 190 17200
rect 280 16960 520 17200
rect 610 16960 850 17200
rect 940 16960 1180 17200
rect 1270 16960 1510 17200
rect 1600 16960 1840 17200
rect 1930 16960 2170 17200
rect 2260 16960 2500 17200
rect 2590 16960 2830 17200
rect 2920 16960 3160 17200
rect 3250 16960 3490 17200
rect 3580 16960 3820 17200
rect 3910 16960 4150 17200
rect 4240 16960 4480 17200
rect 4570 16960 4810 17200
rect 4900 16960 5140 17200
rect 5230 16960 5470 17200
rect 5560 16960 5800 17200
rect 5890 16960 6130 17200
rect 6220 16960 6460 17200
rect 6550 16960 6790 17200
rect 6880 16960 7120 17200
rect -4670 16630 -4430 16870
rect -4340 16630 -4100 16870
rect -4010 16630 -3770 16870
rect -3680 16630 -3440 16870
rect -3350 16630 -3110 16870
rect -3020 16630 -2780 16870
rect -2690 16630 -2450 16870
rect -2360 16630 -2120 16870
rect -2030 16630 -1790 16870
rect -1700 16630 -1460 16870
rect -1370 16630 -1130 16870
rect -1040 16630 -800 16870
rect -710 16630 -470 16870
rect -380 16630 -140 16870
rect -50 16630 190 16870
rect 280 16630 520 16870
rect 610 16630 850 16870
rect 940 16630 1180 16870
rect 1270 16630 1510 16870
rect 1600 16630 1840 16870
rect 1930 16630 2170 16870
rect 2260 16630 2500 16870
rect 2590 16630 2830 16870
rect 2920 16630 3160 16870
rect 3250 16630 3490 16870
rect 3580 16630 3820 16870
rect 3910 16630 4150 16870
rect 4240 16630 4480 16870
rect 4570 16630 4810 16870
rect 4900 16630 5140 16870
rect 5230 16630 5470 16870
rect 5560 16630 5800 16870
rect 5890 16630 6130 16870
rect 6220 16630 6460 16870
rect 6550 16630 6790 16870
rect 6880 16630 7120 16870
rect -4670 16300 -4430 16540
rect -4340 16300 -4100 16540
rect -4010 16300 -3770 16540
rect -3680 16300 -3440 16540
rect -3350 16300 -3110 16540
rect -3020 16300 -2780 16540
rect -2690 16300 -2450 16540
rect -2360 16300 -2120 16540
rect -2030 16300 -1790 16540
rect -1700 16300 -1460 16540
rect -1370 16300 -1130 16540
rect -1040 16300 -800 16540
rect -710 16300 -470 16540
rect -380 16300 -140 16540
rect -50 16300 190 16540
rect 280 16300 520 16540
rect 610 16300 850 16540
rect 940 16300 1180 16540
rect 1270 16300 1510 16540
rect 1600 16300 1840 16540
rect 1930 16300 2170 16540
rect 2260 16300 2500 16540
rect 2590 16300 2830 16540
rect 2920 16300 3160 16540
rect 3250 16300 3490 16540
rect 3580 16300 3820 16540
rect 3910 16300 4150 16540
rect 4240 16300 4480 16540
rect 4570 16300 4810 16540
rect 4900 16300 5140 16540
rect 5230 16300 5470 16540
rect 5560 16300 5800 16540
rect 5890 16300 6130 16540
rect 6220 16300 6460 16540
rect 6550 16300 6790 16540
rect 6880 16300 7120 16540
rect -4670 15970 -4430 16210
rect -4340 15970 -4100 16210
rect -4010 15970 -3770 16210
rect -3680 15970 -3440 16210
rect -3350 15970 -3110 16210
rect -3020 15970 -2780 16210
rect -2690 15970 -2450 16210
rect -2360 15970 -2120 16210
rect -2030 15970 -1790 16210
rect -1700 15970 -1460 16210
rect -1370 15970 -1130 16210
rect -1040 15970 -800 16210
rect -710 15970 -470 16210
rect -380 15970 -140 16210
rect -50 15970 190 16210
rect 280 15970 520 16210
rect 610 15970 850 16210
rect 940 15970 1180 16210
rect 1270 15970 1510 16210
rect 1600 15970 1840 16210
rect 1930 15970 2170 16210
rect 2260 15970 2500 16210
rect 2590 15970 2830 16210
rect 2920 15970 3160 16210
rect 3250 15970 3490 16210
rect 3580 15970 3820 16210
rect 3910 15970 4150 16210
rect 4240 15970 4480 16210
rect 4570 15970 4810 16210
rect 4900 15970 5140 16210
rect 5230 15970 5470 16210
rect 5560 15970 5800 16210
rect 5890 15970 6130 16210
rect 6220 15970 6460 16210
rect 6550 15970 6790 16210
rect 6880 15970 7120 16210
rect -4670 15640 -4430 15880
rect -4340 15640 -4100 15880
rect -4010 15640 -3770 15880
rect -3680 15640 -3440 15880
rect -3350 15640 -3110 15880
rect -3020 15640 -2780 15880
rect -2690 15640 -2450 15880
rect -2360 15640 -2120 15880
rect -2030 15640 -1790 15880
rect -1700 15640 -1460 15880
rect -1370 15640 -1130 15880
rect -1040 15640 -800 15880
rect -710 15640 -470 15880
rect -380 15640 -140 15880
rect -50 15640 190 15880
rect 280 15640 520 15880
rect 610 15640 850 15880
rect 940 15640 1180 15880
rect 1270 15640 1510 15880
rect 1600 15640 1840 15880
rect 1930 15640 2170 15880
rect 2260 15640 2500 15880
rect 2590 15640 2830 15880
rect 2920 15640 3160 15880
rect 3250 15640 3490 15880
rect 3580 15640 3820 15880
rect 3910 15640 4150 15880
rect 4240 15640 4480 15880
rect 4570 15640 4810 15880
rect 4900 15640 5140 15880
rect 5230 15640 5470 15880
rect 5560 15640 5800 15880
rect 5890 15640 6130 15880
rect 6220 15640 6460 15880
rect 6550 15640 6790 15880
rect 6880 15640 7120 15880
rect -4670 15310 -4430 15550
rect -4340 15310 -4100 15550
rect -4010 15310 -3770 15550
rect -3680 15310 -3440 15550
rect -3350 15310 -3110 15550
rect -3020 15310 -2780 15550
rect -2690 15310 -2450 15550
rect -2360 15310 -2120 15550
rect -2030 15310 -1790 15550
rect -1700 15310 -1460 15550
rect -1370 15310 -1130 15550
rect -1040 15310 -800 15550
rect -710 15310 -470 15550
rect -380 15310 -140 15550
rect -50 15310 190 15550
rect 280 15310 520 15550
rect 610 15310 850 15550
rect 940 15310 1180 15550
rect 1270 15310 1510 15550
rect 1600 15310 1840 15550
rect 1930 15310 2170 15550
rect 2260 15310 2500 15550
rect 2590 15310 2830 15550
rect 2920 15310 3160 15550
rect 3250 15310 3490 15550
rect 3580 15310 3820 15550
rect 3910 15310 4150 15550
rect 4240 15310 4480 15550
rect 4570 15310 4810 15550
rect 4900 15310 5140 15550
rect 5230 15310 5470 15550
rect 5560 15310 5800 15550
rect 5890 15310 6130 15550
rect 6220 15310 6460 15550
rect 6550 15310 6790 15550
rect 6880 15310 7120 15550
rect -4670 14980 -4430 15220
rect -4340 14980 -4100 15220
rect -4010 14980 -3770 15220
rect -3680 14980 -3440 15220
rect -3350 14980 -3110 15220
rect -3020 14980 -2780 15220
rect -2690 14980 -2450 15220
rect -2360 14980 -2120 15220
rect -2030 14980 -1790 15220
rect -1700 14980 -1460 15220
rect -1370 14980 -1130 15220
rect -1040 14980 -800 15220
rect -710 14980 -470 15220
rect -380 14980 -140 15220
rect -50 14980 190 15220
rect 280 14980 520 15220
rect 610 14980 850 15220
rect 940 14980 1180 15220
rect 1270 14980 1510 15220
rect 1600 14980 1840 15220
rect 1930 14980 2170 15220
rect 2260 14980 2500 15220
rect 2590 14980 2830 15220
rect 2920 14980 3160 15220
rect 3250 14980 3490 15220
rect 3580 14980 3820 15220
rect 3910 14980 4150 15220
rect 4240 14980 4480 15220
rect 4570 14980 4810 15220
rect 4900 14980 5140 15220
rect 5230 14980 5470 15220
rect 5560 14980 5800 15220
rect 5890 14980 6130 15220
rect 6220 14980 6460 15220
rect 6550 14980 6790 15220
rect 6880 14980 7120 15220
rect -4670 14650 -4430 14890
rect -4340 14650 -4100 14890
rect -4010 14650 -3770 14890
rect -3680 14650 -3440 14890
rect -3350 14650 -3110 14890
rect -3020 14650 -2780 14890
rect -2690 14650 -2450 14890
rect -2360 14650 -2120 14890
rect -2030 14650 -1790 14890
rect -1700 14650 -1460 14890
rect -1370 14650 -1130 14890
rect -1040 14650 -800 14890
rect -710 14650 -470 14890
rect -380 14650 -140 14890
rect -50 14650 190 14890
rect 280 14650 520 14890
rect 610 14650 850 14890
rect 940 14650 1180 14890
rect 1270 14650 1510 14890
rect 1600 14650 1840 14890
rect 1930 14650 2170 14890
rect 2260 14650 2500 14890
rect 2590 14650 2830 14890
rect 2920 14650 3160 14890
rect 3250 14650 3490 14890
rect 3580 14650 3820 14890
rect 3910 14650 4150 14890
rect 4240 14650 4480 14890
rect 4570 14650 4810 14890
rect 4900 14650 5140 14890
rect 5230 14650 5470 14890
rect 5560 14650 5800 14890
rect 5890 14650 6130 14890
rect 6220 14650 6460 14890
rect 6550 14650 6790 14890
rect 6880 14650 7120 14890
rect -4670 14320 -4430 14560
rect -4340 14320 -4100 14560
rect -4010 14320 -3770 14560
rect -3680 14320 -3440 14560
rect -3350 14320 -3110 14560
rect -3020 14320 -2780 14560
rect -2690 14320 -2450 14560
rect -2360 14320 -2120 14560
rect -2030 14320 -1790 14560
rect -1700 14320 -1460 14560
rect -1370 14320 -1130 14560
rect -1040 14320 -800 14560
rect -710 14320 -470 14560
rect -380 14320 -140 14560
rect -50 14320 190 14560
rect 280 14320 520 14560
rect 610 14320 850 14560
rect 940 14320 1180 14560
rect 1270 14320 1510 14560
rect 1600 14320 1840 14560
rect 1930 14320 2170 14560
rect 2260 14320 2500 14560
rect 2590 14320 2830 14560
rect 2920 14320 3160 14560
rect 3250 14320 3490 14560
rect 3580 14320 3820 14560
rect 3910 14320 4150 14560
rect 4240 14320 4480 14560
rect 4570 14320 4810 14560
rect 4900 14320 5140 14560
rect 5230 14320 5470 14560
rect 5560 14320 5800 14560
rect 5890 14320 6130 14560
rect 6220 14320 6460 14560
rect 6550 14320 6790 14560
rect 6880 14320 7120 14560
rect -4670 13990 -4430 14230
rect -4340 13990 -4100 14230
rect -4010 13990 -3770 14230
rect -3680 13990 -3440 14230
rect -3350 13990 -3110 14230
rect -3020 13990 -2780 14230
rect -2690 13990 -2450 14230
rect -2360 13990 -2120 14230
rect -2030 13990 -1790 14230
rect -1700 13990 -1460 14230
rect -1370 13990 -1130 14230
rect -1040 13990 -800 14230
rect -710 13990 -470 14230
rect -380 13990 -140 14230
rect -50 13990 190 14230
rect 280 13990 520 14230
rect 610 13990 850 14230
rect 940 13990 1180 14230
rect 1270 13990 1510 14230
rect 1600 13990 1840 14230
rect 1930 13990 2170 14230
rect 2260 13990 2500 14230
rect 2590 13990 2830 14230
rect 2920 13990 3160 14230
rect 3250 13990 3490 14230
rect 3580 13990 3820 14230
rect 3910 13990 4150 14230
rect 4240 13990 4480 14230
rect 4570 13990 4810 14230
rect 4900 13990 5140 14230
rect 5230 13990 5470 14230
rect 5560 13990 5800 14230
rect 5890 13990 6130 14230
rect 6220 13990 6460 14230
rect 6550 13990 6790 14230
rect 6880 13990 7120 14230
rect -4670 13660 -4430 13900
rect -4340 13660 -4100 13900
rect -4010 13660 -3770 13900
rect -3680 13660 -3440 13900
rect -3350 13660 -3110 13900
rect -3020 13660 -2780 13900
rect -2690 13660 -2450 13900
rect -2360 13660 -2120 13900
rect -2030 13660 -1790 13900
rect -1700 13660 -1460 13900
rect -1370 13660 -1130 13900
rect -1040 13660 -800 13900
rect -710 13660 -470 13900
rect -380 13660 -140 13900
rect -50 13660 190 13900
rect 280 13660 520 13900
rect 610 13660 850 13900
rect 940 13660 1180 13900
rect 1270 13660 1510 13900
rect 1600 13660 1840 13900
rect 1930 13660 2170 13900
rect 2260 13660 2500 13900
rect 2590 13660 2830 13900
rect 2920 13660 3160 13900
rect 3250 13660 3490 13900
rect 3580 13660 3820 13900
rect 3910 13660 4150 13900
rect 4240 13660 4480 13900
rect 4570 13660 4810 13900
rect 4900 13660 5140 13900
rect 5230 13660 5470 13900
rect 5560 13660 5800 13900
rect 5890 13660 6130 13900
rect 6220 13660 6460 13900
rect 6550 13660 6790 13900
rect 6880 13660 7120 13900
rect -4670 13330 -4430 13570
rect -4340 13330 -4100 13570
rect -4010 13330 -3770 13570
rect -3680 13330 -3440 13570
rect -3350 13330 -3110 13570
rect -3020 13330 -2780 13570
rect -2690 13330 -2450 13570
rect -2360 13330 -2120 13570
rect -2030 13330 -1790 13570
rect -1700 13330 -1460 13570
rect -1370 13330 -1130 13570
rect -1040 13330 -800 13570
rect -710 13330 -470 13570
rect -380 13330 -140 13570
rect -50 13330 190 13570
rect 280 13330 520 13570
rect 610 13330 850 13570
rect 940 13330 1180 13570
rect 1270 13330 1510 13570
rect 1600 13330 1840 13570
rect 1930 13330 2170 13570
rect 2260 13330 2500 13570
rect 2590 13330 2830 13570
rect 2920 13330 3160 13570
rect 3250 13330 3490 13570
rect 3580 13330 3820 13570
rect 3910 13330 4150 13570
rect 4240 13330 4480 13570
rect 4570 13330 4810 13570
rect 4900 13330 5140 13570
rect 5230 13330 5470 13570
rect 5560 13330 5800 13570
rect 5890 13330 6130 13570
rect 6220 13330 6460 13570
rect 6550 13330 6790 13570
rect 6880 13330 7120 13570
rect -4670 13000 -4430 13240
rect -4340 13000 -4100 13240
rect -4010 13000 -3770 13240
rect -3680 13000 -3440 13240
rect -3350 13000 -3110 13240
rect -3020 13000 -2780 13240
rect -2690 13000 -2450 13240
rect -2360 13000 -2120 13240
rect -2030 13000 -1790 13240
rect -1700 13000 -1460 13240
rect -1370 13000 -1130 13240
rect -1040 13000 -800 13240
rect -710 13000 -470 13240
rect -380 13000 -140 13240
rect -50 13000 190 13240
rect 280 13000 520 13240
rect 610 13000 850 13240
rect 940 13000 1180 13240
rect 1270 13000 1510 13240
rect 1600 13000 1840 13240
rect 1930 13000 2170 13240
rect 2260 13000 2500 13240
rect 2590 13000 2830 13240
rect 2920 13000 3160 13240
rect 3250 13000 3490 13240
rect 3580 13000 3820 13240
rect 3910 13000 4150 13240
rect 4240 13000 4480 13240
rect 4570 13000 4810 13240
rect 4900 13000 5140 13240
rect 5230 13000 5470 13240
rect 5560 13000 5800 13240
rect 5890 13000 6130 13240
rect 6220 13000 6460 13240
rect 6550 13000 6790 13240
rect 6880 13000 7120 13240
rect -4670 12670 -4430 12910
rect -4340 12670 -4100 12910
rect -4010 12670 -3770 12910
rect -3680 12670 -3440 12910
rect -3350 12670 -3110 12910
rect -3020 12670 -2780 12910
rect -2690 12670 -2450 12910
rect -2360 12670 -2120 12910
rect -2030 12670 -1790 12910
rect -1700 12670 -1460 12910
rect -1370 12670 -1130 12910
rect -1040 12670 -800 12910
rect -710 12670 -470 12910
rect -380 12670 -140 12910
rect -50 12670 190 12910
rect 280 12670 520 12910
rect 610 12670 850 12910
rect 940 12670 1180 12910
rect 1270 12670 1510 12910
rect 1600 12670 1840 12910
rect 1930 12670 2170 12910
rect 2260 12670 2500 12910
rect 2590 12670 2830 12910
rect 2920 12670 3160 12910
rect 3250 12670 3490 12910
rect 3580 12670 3820 12910
rect 3910 12670 4150 12910
rect 4240 12670 4480 12910
rect 4570 12670 4810 12910
rect 4900 12670 5140 12910
rect 5230 12670 5470 12910
rect 5560 12670 5800 12910
rect 5890 12670 6130 12910
rect 6220 12670 6460 12910
rect 6550 12670 6790 12910
rect 6880 12670 7120 12910
rect -4670 12340 -4430 12580
rect -4340 12340 -4100 12580
rect -4010 12340 -3770 12580
rect -3680 12340 -3440 12580
rect -3350 12340 -3110 12580
rect -3020 12340 -2780 12580
rect -2690 12340 -2450 12580
rect -2360 12340 -2120 12580
rect -2030 12340 -1790 12580
rect -1700 12340 -1460 12580
rect -1370 12340 -1130 12580
rect -1040 12340 -800 12580
rect -710 12340 -470 12580
rect -380 12340 -140 12580
rect -50 12340 190 12580
rect 280 12340 520 12580
rect 610 12340 850 12580
rect 940 12340 1180 12580
rect 1270 12340 1510 12580
rect 1600 12340 1840 12580
rect 1930 12340 2170 12580
rect 2260 12340 2500 12580
rect 2590 12340 2830 12580
rect 2920 12340 3160 12580
rect 3250 12340 3490 12580
rect 3580 12340 3820 12580
rect 3910 12340 4150 12580
rect 4240 12340 4480 12580
rect 4570 12340 4810 12580
rect 4900 12340 5140 12580
rect 5230 12340 5470 12580
rect 5560 12340 5800 12580
rect 5890 12340 6130 12580
rect 6220 12340 6460 12580
rect 6550 12340 6790 12580
rect 6880 12340 7120 12580
rect -4670 12010 -4430 12250
rect -4340 12010 -4100 12250
rect -4010 12010 -3770 12250
rect -3680 12010 -3440 12250
rect -3350 12010 -3110 12250
rect -3020 12010 -2780 12250
rect -2690 12010 -2450 12250
rect -2360 12010 -2120 12250
rect -2030 12010 -1790 12250
rect -1700 12010 -1460 12250
rect -1370 12010 -1130 12250
rect -1040 12010 -800 12250
rect -710 12010 -470 12250
rect -380 12010 -140 12250
rect -50 12010 190 12250
rect 280 12010 520 12250
rect 610 12010 850 12250
rect 940 12010 1180 12250
rect 1270 12010 1510 12250
rect 1600 12010 1840 12250
rect 1930 12010 2170 12250
rect 2260 12010 2500 12250
rect 2590 12010 2830 12250
rect 2920 12010 3160 12250
rect 3250 12010 3490 12250
rect 3580 12010 3820 12250
rect 3910 12010 4150 12250
rect 4240 12010 4480 12250
rect 4570 12010 4810 12250
rect 4900 12010 5140 12250
rect 5230 12010 5470 12250
rect 5560 12010 5800 12250
rect 5890 12010 6130 12250
rect 6220 12010 6460 12250
rect 6550 12010 6790 12250
rect 6880 12010 7120 12250
rect -4670 11680 -4430 11920
rect -4340 11680 -4100 11920
rect -4010 11680 -3770 11920
rect -3680 11680 -3440 11920
rect -3350 11680 -3110 11920
rect -3020 11680 -2780 11920
rect -2690 11680 -2450 11920
rect -2360 11680 -2120 11920
rect -2030 11680 -1790 11920
rect -1700 11680 -1460 11920
rect -1370 11680 -1130 11920
rect -1040 11680 -800 11920
rect -710 11680 -470 11920
rect -380 11680 -140 11920
rect -50 11680 190 11920
rect 280 11680 520 11920
rect 610 11680 850 11920
rect 940 11680 1180 11920
rect 1270 11680 1510 11920
rect 1600 11680 1840 11920
rect 1930 11680 2170 11920
rect 2260 11680 2500 11920
rect 2590 11680 2830 11920
rect 2920 11680 3160 11920
rect 3250 11680 3490 11920
rect 3580 11680 3820 11920
rect 3910 11680 4150 11920
rect 4240 11680 4480 11920
rect 4570 11680 4810 11920
rect 4900 11680 5140 11920
rect 5230 11680 5470 11920
rect 5560 11680 5800 11920
rect 5890 11680 6130 11920
rect 6220 11680 6460 11920
rect 6550 11680 6790 11920
rect 6880 11680 7120 11920
rect -4670 11350 -4430 11590
rect -4340 11350 -4100 11590
rect -4010 11350 -3770 11590
rect -3680 11350 -3440 11590
rect -3350 11350 -3110 11590
rect -3020 11350 -2780 11590
rect -2690 11350 -2450 11590
rect -2360 11350 -2120 11590
rect -2030 11350 -1790 11590
rect -1700 11350 -1460 11590
rect -1370 11350 -1130 11590
rect -1040 11350 -800 11590
rect -710 11350 -470 11590
rect -380 11350 -140 11590
rect -50 11350 190 11590
rect 280 11350 520 11590
rect 610 11350 850 11590
rect 940 11350 1180 11590
rect 1270 11350 1510 11590
rect 1600 11350 1840 11590
rect 1930 11350 2170 11590
rect 2260 11350 2500 11590
rect 2590 11350 2830 11590
rect 2920 11350 3160 11590
rect 3250 11350 3490 11590
rect 3580 11350 3820 11590
rect 3910 11350 4150 11590
rect 4240 11350 4480 11590
rect 4570 11350 4810 11590
rect 4900 11350 5140 11590
rect 5230 11350 5470 11590
rect 5560 11350 5800 11590
rect 5890 11350 6130 11590
rect 6220 11350 6460 11590
rect 6550 11350 6790 11590
rect 6880 11350 7120 11590
rect -4670 11020 -4430 11260
rect -4340 11020 -4100 11260
rect -4010 11020 -3770 11260
rect -3680 11020 -3440 11260
rect -3350 11020 -3110 11260
rect -3020 11020 -2780 11260
rect -2690 11020 -2450 11260
rect -2360 11020 -2120 11260
rect -2030 11020 -1790 11260
rect -1700 11020 -1460 11260
rect -1370 11020 -1130 11260
rect -1040 11020 -800 11260
rect -710 11020 -470 11260
rect -380 11020 -140 11260
rect -50 11020 190 11260
rect 280 11020 520 11260
rect 610 11020 850 11260
rect 940 11020 1180 11260
rect 1270 11020 1510 11260
rect 1600 11020 1840 11260
rect 1930 11020 2170 11260
rect 2260 11020 2500 11260
rect 2590 11020 2830 11260
rect 2920 11020 3160 11260
rect 3250 11020 3490 11260
rect 3580 11020 3820 11260
rect 3910 11020 4150 11260
rect 4240 11020 4480 11260
rect 4570 11020 4810 11260
rect 4900 11020 5140 11260
rect 5230 11020 5470 11260
rect 5560 11020 5800 11260
rect 5890 11020 6130 11260
rect 6220 11020 6460 11260
rect 6550 11020 6790 11260
rect 6880 11020 7120 11260
rect -4670 10690 -4430 10930
rect -4340 10690 -4100 10930
rect -4010 10690 -3770 10930
rect -3680 10690 -3440 10930
rect -3350 10690 -3110 10930
rect -3020 10690 -2780 10930
rect -2690 10690 -2450 10930
rect -2360 10690 -2120 10930
rect -2030 10690 -1790 10930
rect -1700 10690 -1460 10930
rect -1370 10690 -1130 10930
rect -1040 10690 -800 10930
rect -710 10690 -470 10930
rect -380 10690 -140 10930
rect -50 10690 190 10930
rect 280 10690 520 10930
rect 610 10690 850 10930
rect 940 10690 1180 10930
rect 1270 10690 1510 10930
rect 1600 10690 1840 10930
rect 1930 10690 2170 10930
rect 2260 10690 2500 10930
rect 2590 10690 2830 10930
rect 2920 10690 3160 10930
rect 3250 10690 3490 10930
rect 3580 10690 3820 10930
rect 3910 10690 4150 10930
rect 4240 10690 4480 10930
rect 4570 10690 4810 10930
rect 4900 10690 5140 10930
rect 5230 10690 5470 10930
rect 5560 10690 5800 10930
rect 5890 10690 6130 10930
rect 6220 10690 6460 10930
rect 6550 10690 6790 10930
rect 6880 10690 7120 10930
rect -4670 10360 -4430 10600
rect -4340 10360 -4100 10600
rect -4010 10360 -3770 10600
rect -3680 10360 -3440 10600
rect -3350 10360 -3110 10600
rect -3020 10360 -2780 10600
rect -2690 10360 -2450 10600
rect -2360 10360 -2120 10600
rect -2030 10360 -1790 10600
rect -1700 10360 -1460 10600
rect -1370 10360 -1130 10600
rect -1040 10360 -800 10600
rect -710 10360 -470 10600
rect -380 10360 -140 10600
rect -50 10360 190 10600
rect 280 10360 520 10600
rect 610 10360 850 10600
rect 940 10360 1180 10600
rect 1270 10360 1510 10600
rect 1600 10360 1840 10600
rect 1930 10360 2170 10600
rect 2260 10360 2500 10600
rect 2590 10360 2830 10600
rect 2920 10360 3160 10600
rect 3250 10360 3490 10600
rect 3580 10360 3820 10600
rect 3910 10360 4150 10600
rect 4240 10360 4480 10600
rect 4570 10360 4810 10600
rect 4900 10360 5140 10600
rect 5230 10360 5470 10600
rect 5560 10360 5800 10600
rect 5890 10360 6130 10600
rect 6220 10360 6460 10600
rect 6550 10360 6790 10600
rect 6880 10360 7120 10600
rect -4670 10030 -4430 10270
rect -4340 10030 -4100 10270
rect -4010 10030 -3770 10270
rect -3680 10030 -3440 10270
rect -3350 10030 -3110 10270
rect -3020 10030 -2780 10270
rect -2690 10030 -2450 10270
rect -2360 10030 -2120 10270
rect -2030 10030 -1790 10270
rect -1700 10030 -1460 10270
rect -1370 10030 -1130 10270
rect -1040 10030 -800 10270
rect -710 10030 -470 10270
rect -380 10030 -140 10270
rect -50 10030 190 10270
rect 280 10030 520 10270
rect 610 10030 850 10270
rect 940 10030 1180 10270
rect 1270 10030 1510 10270
rect 1600 10030 1840 10270
rect 1930 10030 2170 10270
rect 2260 10030 2500 10270
rect 2590 10030 2830 10270
rect 2920 10030 3160 10270
rect 3250 10030 3490 10270
rect 3580 10030 3820 10270
rect 3910 10030 4150 10270
rect 4240 10030 4480 10270
rect 4570 10030 4810 10270
rect 4900 10030 5140 10270
rect 5230 10030 5470 10270
rect 5560 10030 5800 10270
rect 5890 10030 6130 10270
rect 6220 10030 6460 10270
rect 6550 10030 6790 10270
rect 6880 10030 7120 10270
rect -4670 9700 -4430 9940
rect -4340 9700 -4100 9940
rect -4010 9700 -3770 9940
rect -3680 9700 -3440 9940
rect -3350 9700 -3110 9940
rect -3020 9700 -2780 9940
rect -2690 9700 -2450 9940
rect -2360 9700 -2120 9940
rect -2030 9700 -1790 9940
rect -1700 9700 -1460 9940
rect -1370 9700 -1130 9940
rect -1040 9700 -800 9940
rect -710 9700 -470 9940
rect -380 9700 -140 9940
rect -50 9700 190 9940
rect 280 9700 520 9940
rect 610 9700 850 9940
rect 940 9700 1180 9940
rect 1270 9700 1510 9940
rect 1600 9700 1840 9940
rect 1930 9700 2170 9940
rect 2260 9700 2500 9940
rect 2590 9700 2830 9940
rect 2920 9700 3160 9940
rect 3250 9700 3490 9940
rect 3580 9700 3820 9940
rect 3910 9700 4150 9940
rect 4240 9700 4480 9940
rect 4570 9700 4810 9940
rect 4900 9700 5140 9940
rect 5230 9700 5470 9940
rect 5560 9700 5800 9940
rect 5890 9700 6130 9940
rect 6220 9700 6460 9940
rect 6550 9700 6790 9940
rect 6880 9700 7120 9940
rect -4670 9370 -4430 9610
rect -4340 9370 -4100 9610
rect -4010 9370 -3770 9610
rect -3680 9370 -3440 9610
rect -3350 9370 -3110 9610
rect -3020 9370 -2780 9610
rect -2690 9370 -2450 9610
rect -2360 9370 -2120 9610
rect -2030 9370 -1790 9610
rect -1700 9370 -1460 9610
rect -1370 9370 -1130 9610
rect -1040 9370 -800 9610
rect -710 9370 -470 9610
rect -380 9370 -140 9610
rect -50 9370 190 9610
rect 280 9370 520 9610
rect 610 9370 850 9610
rect 940 9370 1180 9610
rect 1270 9370 1510 9610
rect 1600 9370 1840 9610
rect 1930 9370 2170 9610
rect 2260 9370 2500 9610
rect 2590 9370 2830 9610
rect 2920 9370 3160 9610
rect 3250 9370 3490 9610
rect 3580 9370 3820 9610
rect 3910 9370 4150 9610
rect 4240 9370 4480 9610
rect 4570 9370 4810 9610
rect 4900 9370 5140 9610
rect 5230 9370 5470 9610
rect 5560 9370 5800 9610
rect 5890 9370 6130 9610
rect 6220 9370 6460 9610
rect 6550 9370 6790 9610
rect 6880 9370 7120 9610
rect -4670 9040 -4430 9280
rect -4340 9040 -4100 9280
rect -4010 9040 -3770 9280
rect -3680 9040 -3440 9280
rect -3350 9040 -3110 9280
rect -3020 9040 -2780 9280
rect -2690 9040 -2450 9280
rect -2360 9040 -2120 9280
rect -2030 9040 -1790 9280
rect -1700 9040 -1460 9280
rect -1370 9040 -1130 9280
rect -1040 9040 -800 9280
rect -710 9040 -470 9280
rect -380 9040 -140 9280
rect -50 9040 190 9280
rect 280 9040 520 9280
rect 610 9040 850 9280
rect 940 9040 1180 9280
rect 1270 9040 1510 9280
rect 1600 9040 1840 9280
rect 1930 9040 2170 9280
rect 2260 9040 2500 9280
rect 2590 9040 2830 9280
rect 2920 9040 3160 9280
rect 3250 9040 3490 9280
rect 3580 9040 3820 9280
rect 3910 9040 4150 9280
rect 4240 9040 4480 9280
rect 4570 9040 4810 9280
rect 4900 9040 5140 9280
rect 5230 9040 5470 9280
rect 5560 9040 5800 9280
rect 5890 9040 6130 9280
rect 6220 9040 6460 9280
rect 6550 9040 6790 9280
rect 6880 9040 7120 9280
rect 7780 20590 8020 20830
rect 8110 20590 8350 20830
rect 8440 20590 8680 20830
rect 8770 20590 9010 20830
rect 9100 20590 9340 20830
rect 9430 20590 9670 20830
rect 9760 20590 10000 20830
rect 10090 20590 10330 20830
rect 10420 20590 10660 20830
rect 10750 20590 10990 20830
rect 11080 20590 11320 20830
rect 11410 20590 11650 20830
rect 11740 20590 11980 20830
rect 12070 20590 12310 20830
rect 12400 20590 12640 20830
rect 12730 20590 12970 20830
rect 13060 20590 13300 20830
rect 13390 20590 13630 20830
rect 13720 20590 13960 20830
rect 14050 20590 14290 20830
rect 14380 20590 14620 20830
rect 14710 20590 14950 20830
rect 15040 20590 15280 20830
rect 15370 20590 15610 20830
rect 15700 20590 15940 20830
rect 16030 20590 16270 20830
rect 16360 20590 16600 20830
rect 16690 20590 16930 20830
rect 17020 20590 17260 20830
rect 17350 20590 17590 20830
rect 17680 20590 17920 20830
rect 18010 20590 18250 20830
rect 18340 20590 18580 20830
rect 18670 20590 18910 20830
rect 19000 20590 19240 20830
rect 19330 20590 19570 20830
rect 7780 20260 8020 20500
rect 8110 20260 8350 20500
rect 8440 20260 8680 20500
rect 8770 20260 9010 20500
rect 9100 20260 9340 20500
rect 9430 20260 9670 20500
rect 9760 20260 10000 20500
rect 10090 20260 10330 20500
rect 10420 20260 10660 20500
rect 10750 20260 10990 20500
rect 11080 20260 11320 20500
rect 11410 20260 11650 20500
rect 11740 20260 11980 20500
rect 12070 20260 12310 20500
rect 12400 20260 12640 20500
rect 12730 20260 12970 20500
rect 13060 20260 13300 20500
rect 13390 20260 13630 20500
rect 13720 20260 13960 20500
rect 14050 20260 14290 20500
rect 14380 20260 14620 20500
rect 14710 20260 14950 20500
rect 15040 20260 15280 20500
rect 15370 20260 15610 20500
rect 15700 20260 15940 20500
rect 16030 20260 16270 20500
rect 16360 20260 16600 20500
rect 16690 20260 16930 20500
rect 17020 20260 17260 20500
rect 17350 20260 17590 20500
rect 17680 20260 17920 20500
rect 18010 20260 18250 20500
rect 18340 20260 18580 20500
rect 18670 20260 18910 20500
rect 19000 20260 19240 20500
rect 19330 20260 19570 20500
rect 7780 19930 8020 20170
rect 8110 19930 8350 20170
rect 8440 19930 8680 20170
rect 8770 19930 9010 20170
rect 9100 19930 9340 20170
rect 9430 19930 9670 20170
rect 9760 19930 10000 20170
rect 10090 19930 10330 20170
rect 10420 19930 10660 20170
rect 10750 19930 10990 20170
rect 11080 19930 11320 20170
rect 11410 19930 11650 20170
rect 11740 19930 11980 20170
rect 12070 19930 12310 20170
rect 12400 19930 12640 20170
rect 12730 19930 12970 20170
rect 13060 19930 13300 20170
rect 13390 19930 13630 20170
rect 13720 19930 13960 20170
rect 14050 19930 14290 20170
rect 14380 19930 14620 20170
rect 14710 19930 14950 20170
rect 15040 19930 15280 20170
rect 15370 19930 15610 20170
rect 15700 19930 15940 20170
rect 16030 19930 16270 20170
rect 16360 19930 16600 20170
rect 16690 19930 16930 20170
rect 17020 19930 17260 20170
rect 17350 19930 17590 20170
rect 17680 19930 17920 20170
rect 18010 19930 18250 20170
rect 18340 19930 18580 20170
rect 18670 19930 18910 20170
rect 19000 19930 19240 20170
rect 19330 19930 19570 20170
rect 7780 19600 8020 19840
rect 8110 19600 8350 19840
rect 8440 19600 8680 19840
rect 8770 19600 9010 19840
rect 9100 19600 9340 19840
rect 9430 19600 9670 19840
rect 9760 19600 10000 19840
rect 10090 19600 10330 19840
rect 10420 19600 10660 19840
rect 10750 19600 10990 19840
rect 11080 19600 11320 19840
rect 11410 19600 11650 19840
rect 11740 19600 11980 19840
rect 12070 19600 12310 19840
rect 12400 19600 12640 19840
rect 12730 19600 12970 19840
rect 13060 19600 13300 19840
rect 13390 19600 13630 19840
rect 13720 19600 13960 19840
rect 14050 19600 14290 19840
rect 14380 19600 14620 19840
rect 14710 19600 14950 19840
rect 15040 19600 15280 19840
rect 15370 19600 15610 19840
rect 15700 19600 15940 19840
rect 16030 19600 16270 19840
rect 16360 19600 16600 19840
rect 16690 19600 16930 19840
rect 17020 19600 17260 19840
rect 17350 19600 17590 19840
rect 17680 19600 17920 19840
rect 18010 19600 18250 19840
rect 18340 19600 18580 19840
rect 18670 19600 18910 19840
rect 19000 19600 19240 19840
rect 19330 19600 19570 19840
rect 7780 19270 8020 19510
rect 8110 19270 8350 19510
rect 8440 19270 8680 19510
rect 8770 19270 9010 19510
rect 9100 19270 9340 19510
rect 9430 19270 9670 19510
rect 9760 19270 10000 19510
rect 10090 19270 10330 19510
rect 10420 19270 10660 19510
rect 10750 19270 10990 19510
rect 11080 19270 11320 19510
rect 11410 19270 11650 19510
rect 11740 19270 11980 19510
rect 12070 19270 12310 19510
rect 12400 19270 12640 19510
rect 12730 19270 12970 19510
rect 13060 19270 13300 19510
rect 13390 19270 13630 19510
rect 13720 19270 13960 19510
rect 14050 19270 14290 19510
rect 14380 19270 14620 19510
rect 14710 19270 14950 19510
rect 15040 19270 15280 19510
rect 15370 19270 15610 19510
rect 15700 19270 15940 19510
rect 16030 19270 16270 19510
rect 16360 19270 16600 19510
rect 16690 19270 16930 19510
rect 17020 19270 17260 19510
rect 17350 19270 17590 19510
rect 17680 19270 17920 19510
rect 18010 19270 18250 19510
rect 18340 19270 18580 19510
rect 18670 19270 18910 19510
rect 19000 19270 19240 19510
rect 19330 19270 19570 19510
rect 7780 18940 8020 19180
rect 8110 18940 8350 19180
rect 8440 18940 8680 19180
rect 8770 18940 9010 19180
rect 9100 18940 9340 19180
rect 9430 18940 9670 19180
rect 9760 18940 10000 19180
rect 10090 18940 10330 19180
rect 10420 18940 10660 19180
rect 10750 18940 10990 19180
rect 11080 18940 11320 19180
rect 11410 18940 11650 19180
rect 11740 18940 11980 19180
rect 12070 18940 12310 19180
rect 12400 18940 12640 19180
rect 12730 18940 12970 19180
rect 13060 18940 13300 19180
rect 13390 18940 13630 19180
rect 13720 18940 13960 19180
rect 14050 18940 14290 19180
rect 14380 18940 14620 19180
rect 14710 18940 14950 19180
rect 15040 18940 15280 19180
rect 15370 18940 15610 19180
rect 15700 18940 15940 19180
rect 16030 18940 16270 19180
rect 16360 18940 16600 19180
rect 16690 18940 16930 19180
rect 17020 18940 17260 19180
rect 17350 18940 17590 19180
rect 17680 18940 17920 19180
rect 18010 18940 18250 19180
rect 18340 18940 18580 19180
rect 18670 18940 18910 19180
rect 19000 18940 19240 19180
rect 19330 18940 19570 19180
rect 7780 18610 8020 18850
rect 8110 18610 8350 18850
rect 8440 18610 8680 18850
rect 8770 18610 9010 18850
rect 9100 18610 9340 18850
rect 9430 18610 9670 18850
rect 9760 18610 10000 18850
rect 10090 18610 10330 18850
rect 10420 18610 10660 18850
rect 10750 18610 10990 18850
rect 11080 18610 11320 18850
rect 11410 18610 11650 18850
rect 11740 18610 11980 18850
rect 12070 18610 12310 18850
rect 12400 18610 12640 18850
rect 12730 18610 12970 18850
rect 13060 18610 13300 18850
rect 13390 18610 13630 18850
rect 13720 18610 13960 18850
rect 14050 18610 14290 18850
rect 14380 18610 14620 18850
rect 14710 18610 14950 18850
rect 15040 18610 15280 18850
rect 15370 18610 15610 18850
rect 15700 18610 15940 18850
rect 16030 18610 16270 18850
rect 16360 18610 16600 18850
rect 16690 18610 16930 18850
rect 17020 18610 17260 18850
rect 17350 18610 17590 18850
rect 17680 18610 17920 18850
rect 18010 18610 18250 18850
rect 18340 18610 18580 18850
rect 18670 18610 18910 18850
rect 19000 18610 19240 18850
rect 19330 18610 19570 18850
rect 7780 18280 8020 18520
rect 8110 18280 8350 18520
rect 8440 18280 8680 18520
rect 8770 18280 9010 18520
rect 9100 18280 9340 18520
rect 9430 18280 9670 18520
rect 9760 18280 10000 18520
rect 10090 18280 10330 18520
rect 10420 18280 10660 18520
rect 10750 18280 10990 18520
rect 11080 18280 11320 18520
rect 11410 18280 11650 18520
rect 11740 18280 11980 18520
rect 12070 18280 12310 18520
rect 12400 18280 12640 18520
rect 12730 18280 12970 18520
rect 13060 18280 13300 18520
rect 13390 18280 13630 18520
rect 13720 18280 13960 18520
rect 14050 18280 14290 18520
rect 14380 18280 14620 18520
rect 14710 18280 14950 18520
rect 15040 18280 15280 18520
rect 15370 18280 15610 18520
rect 15700 18280 15940 18520
rect 16030 18280 16270 18520
rect 16360 18280 16600 18520
rect 16690 18280 16930 18520
rect 17020 18280 17260 18520
rect 17350 18280 17590 18520
rect 17680 18280 17920 18520
rect 18010 18280 18250 18520
rect 18340 18280 18580 18520
rect 18670 18280 18910 18520
rect 19000 18280 19240 18520
rect 19330 18280 19570 18520
rect 7780 17950 8020 18190
rect 8110 17950 8350 18190
rect 8440 17950 8680 18190
rect 8770 17950 9010 18190
rect 9100 17950 9340 18190
rect 9430 17950 9670 18190
rect 9760 17950 10000 18190
rect 10090 17950 10330 18190
rect 10420 17950 10660 18190
rect 10750 17950 10990 18190
rect 11080 17950 11320 18190
rect 11410 17950 11650 18190
rect 11740 17950 11980 18190
rect 12070 17950 12310 18190
rect 12400 17950 12640 18190
rect 12730 17950 12970 18190
rect 13060 17950 13300 18190
rect 13390 17950 13630 18190
rect 13720 17950 13960 18190
rect 14050 17950 14290 18190
rect 14380 17950 14620 18190
rect 14710 17950 14950 18190
rect 15040 17950 15280 18190
rect 15370 17950 15610 18190
rect 15700 17950 15940 18190
rect 16030 17950 16270 18190
rect 16360 17950 16600 18190
rect 16690 17950 16930 18190
rect 17020 17950 17260 18190
rect 17350 17950 17590 18190
rect 17680 17950 17920 18190
rect 18010 17950 18250 18190
rect 18340 17950 18580 18190
rect 18670 17950 18910 18190
rect 19000 17950 19240 18190
rect 19330 17950 19570 18190
rect 7780 17620 8020 17860
rect 8110 17620 8350 17860
rect 8440 17620 8680 17860
rect 8770 17620 9010 17860
rect 9100 17620 9340 17860
rect 9430 17620 9670 17860
rect 9760 17620 10000 17860
rect 10090 17620 10330 17860
rect 10420 17620 10660 17860
rect 10750 17620 10990 17860
rect 11080 17620 11320 17860
rect 11410 17620 11650 17860
rect 11740 17620 11980 17860
rect 12070 17620 12310 17860
rect 12400 17620 12640 17860
rect 12730 17620 12970 17860
rect 13060 17620 13300 17860
rect 13390 17620 13630 17860
rect 13720 17620 13960 17860
rect 14050 17620 14290 17860
rect 14380 17620 14620 17860
rect 14710 17620 14950 17860
rect 15040 17620 15280 17860
rect 15370 17620 15610 17860
rect 15700 17620 15940 17860
rect 16030 17620 16270 17860
rect 16360 17620 16600 17860
rect 16690 17620 16930 17860
rect 17020 17620 17260 17860
rect 17350 17620 17590 17860
rect 17680 17620 17920 17860
rect 18010 17620 18250 17860
rect 18340 17620 18580 17860
rect 18670 17620 18910 17860
rect 19000 17620 19240 17860
rect 19330 17620 19570 17860
rect 7780 17290 8020 17530
rect 8110 17290 8350 17530
rect 8440 17290 8680 17530
rect 8770 17290 9010 17530
rect 9100 17290 9340 17530
rect 9430 17290 9670 17530
rect 9760 17290 10000 17530
rect 10090 17290 10330 17530
rect 10420 17290 10660 17530
rect 10750 17290 10990 17530
rect 11080 17290 11320 17530
rect 11410 17290 11650 17530
rect 11740 17290 11980 17530
rect 12070 17290 12310 17530
rect 12400 17290 12640 17530
rect 12730 17290 12970 17530
rect 13060 17290 13300 17530
rect 13390 17290 13630 17530
rect 13720 17290 13960 17530
rect 14050 17290 14290 17530
rect 14380 17290 14620 17530
rect 14710 17290 14950 17530
rect 15040 17290 15280 17530
rect 15370 17290 15610 17530
rect 15700 17290 15940 17530
rect 16030 17290 16270 17530
rect 16360 17290 16600 17530
rect 16690 17290 16930 17530
rect 17020 17290 17260 17530
rect 17350 17290 17590 17530
rect 17680 17290 17920 17530
rect 18010 17290 18250 17530
rect 18340 17290 18580 17530
rect 18670 17290 18910 17530
rect 19000 17290 19240 17530
rect 19330 17290 19570 17530
rect 7780 16960 8020 17200
rect 8110 16960 8350 17200
rect 8440 16960 8680 17200
rect 8770 16960 9010 17200
rect 9100 16960 9340 17200
rect 9430 16960 9670 17200
rect 9760 16960 10000 17200
rect 10090 16960 10330 17200
rect 10420 16960 10660 17200
rect 10750 16960 10990 17200
rect 11080 16960 11320 17200
rect 11410 16960 11650 17200
rect 11740 16960 11980 17200
rect 12070 16960 12310 17200
rect 12400 16960 12640 17200
rect 12730 16960 12970 17200
rect 13060 16960 13300 17200
rect 13390 16960 13630 17200
rect 13720 16960 13960 17200
rect 14050 16960 14290 17200
rect 14380 16960 14620 17200
rect 14710 16960 14950 17200
rect 15040 16960 15280 17200
rect 15370 16960 15610 17200
rect 15700 16960 15940 17200
rect 16030 16960 16270 17200
rect 16360 16960 16600 17200
rect 16690 16960 16930 17200
rect 17020 16960 17260 17200
rect 17350 16960 17590 17200
rect 17680 16960 17920 17200
rect 18010 16960 18250 17200
rect 18340 16960 18580 17200
rect 18670 16960 18910 17200
rect 19000 16960 19240 17200
rect 19330 16960 19570 17200
rect 7780 16630 8020 16870
rect 8110 16630 8350 16870
rect 8440 16630 8680 16870
rect 8770 16630 9010 16870
rect 9100 16630 9340 16870
rect 9430 16630 9670 16870
rect 9760 16630 10000 16870
rect 10090 16630 10330 16870
rect 10420 16630 10660 16870
rect 10750 16630 10990 16870
rect 11080 16630 11320 16870
rect 11410 16630 11650 16870
rect 11740 16630 11980 16870
rect 12070 16630 12310 16870
rect 12400 16630 12640 16870
rect 12730 16630 12970 16870
rect 13060 16630 13300 16870
rect 13390 16630 13630 16870
rect 13720 16630 13960 16870
rect 14050 16630 14290 16870
rect 14380 16630 14620 16870
rect 14710 16630 14950 16870
rect 15040 16630 15280 16870
rect 15370 16630 15610 16870
rect 15700 16630 15940 16870
rect 16030 16630 16270 16870
rect 16360 16630 16600 16870
rect 16690 16630 16930 16870
rect 17020 16630 17260 16870
rect 17350 16630 17590 16870
rect 17680 16630 17920 16870
rect 18010 16630 18250 16870
rect 18340 16630 18580 16870
rect 18670 16630 18910 16870
rect 19000 16630 19240 16870
rect 19330 16630 19570 16870
rect 7780 16300 8020 16540
rect 8110 16300 8350 16540
rect 8440 16300 8680 16540
rect 8770 16300 9010 16540
rect 9100 16300 9340 16540
rect 9430 16300 9670 16540
rect 9760 16300 10000 16540
rect 10090 16300 10330 16540
rect 10420 16300 10660 16540
rect 10750 16300 10990 16540
rect 11080 16300 11320 16540
rect 11410 16300 11650 16540
rect 11740 16300 11980 16540
rect 12070 16300 12310 16540
rect 12400 16300 12640 16540
rect 12730 16300 12970 16540
rect 13060 16300 13300 16540
rect 13390 16300 13630 16540
rect 13720 16300 13960 16540
rect 14050 16300 14290 16540
rect 14380 16300 14620 16540
rect 14710 16300 14950 16540
rect 15040 16300 15280 16540
rect 15370 16300 15610 16540
rect 15700 16300 15940 16540
rect 16030 16300 16270 16540
rect 16360 16300 16600 16540
rect 16690 16300 16930 16540
rect 17020 16300 17260 16540
rect 17350 16300 17590 16540
rect 17680 16300 17920 16540
rect 18010 16300 18250 16540
rect 18340 16300 18580 16540
rect 18670 16300 18910 16540
rect 19000 16300 19240 16540
rect 19330 16300 19570 16540
rect 7780 15970 8020 16210
rect 8110 15970 8350 16210
rect 8440 15970 8680 16210
rect 8770 15970 9010 16210
rect 9100 15970 9340 16210
rect 9430 15970 9670 16210
rect 9760 15970 10000 16210
rect 10090 15970 10330 16210
rect 10420 15970 10660 16210
rect 10750 15970 10990 16210
rect 11080 15970 11320 16210
rect 11410 15970 11650 16210
rect 11740 15970 11980 16210
rect 12070 15970 12310 16210
rect 12400 15970 12640 16210
rect 12730 15970 12970 16210
rect 13060 15970 13300 16210
rect 13390 15970 13630 16210
rect 13720 15970 13960 16210
rect 14050 15970 14290 16210
rect 14380 15970 14620 16210
rect 14710 15970 14950 16210
rect 15040 15970 15280 16210
rect 15370 15970 15610 16210
rect 15700 15970 15940 16210
rect 16030 15970 16270 16210
rect 16360 15970 16600 16210
rect 16690 15970 16930 16210
rect 17020 15970 17260 16210
rect 17350 15970 17590 16210
rect 17680 15970 17920 16210
rect 18010 15970 18250 16210
rect 18340 15970 18580 16210
rect 18670 15970 18910 16210
rect 19000 15970 19240 16210
rect 19330 15970 19570 16210
rect 7780 15640 8020 15880
rect 8110 15640 8350 15880
rect 8440 15640 8680 15880
rect 8770 15640 9010 15880
rect 9100 15640 9340 15880
rect 9430 15640 9670 15880
rect 9760 15640 10000 15880
rect 10090 15640 10330 15880
rect 10420 15640 10660 15880
rect 10750 15640 10990 15880
rect 11080 15640 11320 15880
rect 11410 15640 11650 15880
rect 11740 15640 11980 15880
rect 12070 15640 12310 15880
rect 12400 15640 12640 15880
rect 12730 15640 12970 15880
rect 13060 15640 13300 15880
rect 13390 15640 13630 15880
rect 13720 15640 13960 15880
rect 14050 15640 14290 15880
rect 14380 15640 14620 15880
rect 14710 15640 14950 15880
rect 15040 15640 15280 15880
rect 15370 15640 15610 15880
rect 15700 15640 15940 15880
rect 16030 15640 16270 15880
rect 16360 15640 16600 15880
rect 16690 15640 16930 15880
rect 17020 15640 17260 15880
rect 17350 15640 17590 15880
rect 17680 15640 17920 15880
rect 18010 15640 18250 15880
rect 18340 15640 18580 15880
rect 18670 15640 18910 15880
rect 19000 15640 19240 15880
rect 19330 15640 19570 15880
rect 7780 15310 8020 15550
rect 8110 15310 8350 15550
rect 8440 15310 8680 15550
rect 8770 15310 9010 15550
rect 9100 15310 9340 15550
rect 9430 15310 9670 15550
rect 9760 15310 10000 15550
rect 10090 15310 10330 15550
rect 10420 15310 10660 15550
rect 10750 15310 10990 15550
rect 11080 15310 11320 15550
rect 11410 15310 11650 15550
rect 11740 15310 11980 15550
rect 12070 15310 12310 15550
rect 12400 15310 12640 15550
rect 12730 15310 12970 15550
rect 13060 15310 13300 15550
rect 13390 15310 13630 15550
rect 13720 15310 13960 15550
rect 14050 15310 14290 15550
rect 14380 15310 14620 15550
rect 14710 15310 14950 15550
rect 15040 15310 15280 15550
rect 15370 15310 15610 15550
rect 15700 15310 15940 15550
rect 16030 15310 16270 15550
rect 16360 15310 16600 15550
rect 16690 15310 16930 15550
rect 17020 15310 17260 15550
rect 17350 15310 17590 15550
rect 17680 15310 17920 15550
rect 18010 15310 18250 15550
rect 18340 15310 18580 15550
rect 18670 15310 18910 15550
rect 19000 15310 19240 15550
rect 19330 15310 19570 15550
rect 7780 14980 8020 15220
rect 8110 14980 8350 15220
rect 8440 14980 8680 15220
rect 8770 14980 9010 15220
rect 9100 14980 9340 15220
rect 9430 14980 9670 15220
rect 9760 14980 10000 15220
rect 10090 14980 10330 15220
rect 10420 14980 10660 15220
rect 10750 14980 10990 15220
rect 11080 14980 11320 15220
rect 11410 14980 11650 15220
rect 11740 14980 11980 15220
rect 12070 14980 12310 15220
rect 12400 14980 12640 15220
rect 12730 14980 12970 15220
rect 13060 14980 13300 15220
rect 13390 14980 13630 15220
rect 13720 14980 13960 15220
rect 14050 14980 14290 15220
rect 14380 14980 14620 15220
rect 14710 14980 14950 15220
rect 15040 14980 15280 15220
rect 15370 14980 15610 15220
rect 15700 14980 15940 15220
rect 16030 14980 16270 15220
rect 16360 14980 16600 15220
rect 16690 14980 16930 15220
rect 17020 14980 17260 15220
rect 17350 14980 17590 15220
rect 17680 14980 17920 15220
rect 18010 14980 18250 15220
rect 18340 14980 18580 15220
rect 18670 14980 18910 15220
rect 19000 14980 19240 15220
rect 19330 14980 19570 15220
rect 7780 14650 8020 14890
rect 8110 14650 8350 14890
rect 8440 14650 8680 14890
rect 8770 14650 9010 14890
rect 9100 14650 9340 14890
rect 9430 14650 9670 14890
rect 9760 14650 10000 14890
rect 10090 14650 10330 14890
rect 10420 14650 10660 14890
rect 10750 14650 10990 14890
rect 11080 14650 11320 14890
rect 11410 14650 11650 14890
rect 11740 14650 11980 14890
rect 12070 14650 12310 14890
rect 12400 14650 12640 14890
rect 12730 14650 12970 14890
rect 13060 14650 13300 14890
rect 13390 14650 13630 14890
rect 13720 14650 13960 14890
rect 14050 14650 14290 14890
rect 14380 14650 14620 14890
rect 14710 14650 14950 14890
rect 15040 14650 15280 14890
rect 15370 14650 15610 14890
rect 15700 14650 15940 14890
rect 16030 14650 16270 14890
rect 16360 14650 16600 14890
rect 16690 14650 16930 14890
rect 17020 14650 17260 14890
rect 17350 14650 17590 14890
rect 17680 14650 17920 14890
rect 18010 14650 18250 14890
rect 18340 14650 18580 14890
rect 18670 14650 18910 14890
rect 19000 14650 19240 14890
rect 19330 14650 19570 14890
rect 7780 14320 8020 14560
rect 8110 14320 8350 14560
rect 8440 14320 8680 14560
rect 8770 14320 9010 14560
rect 9100 14320 9340 14560
rect 9430 14320 9670 14560
rect 9760 14320 10000 14560
rect 10090 14320 10330 14560
rect 10420 14320 10660 14560
rect 10750 14320 10990 14560
rect 11080 14320 11320 14560
rect 11410 14320 11650 14560
rect 11740 14320 11980 14560
rect 12070 14320 12310 14560
rect 12400 14320 12640 14560
rect 12730 14320 12970 14560
rect 13060 14320 13300 14560
rect 13390 14320 13630 14560
rect 13720 14320 13960 14560
rect 14050 14320 14290 14560
rect 14380 14320 14620 14560
rect 14710 14320 14950 14560
rect 15040 14320 15280 14560
rect 15370 14320 15610 14560
rect 15700 14320 15940 14560
rect 16030 14320 16270 14560
rect 16360 14320 16600 14560
rect 16690 14320 16930 14560
rect 17020 14320 17260 14560
rect 17350 14320 17590 14560
rect 17680 14320 17920 14560
rect 18010 14320 18250 14560
rect 18340 14320 18580 14560
rect 18670 14320 18910 14560
rect 19000 14320 19240 14560
rect 19330 14320 19570 14560
rect 7780 13990 8020 14230
rect 8110 13990 8350 14230
rect 8440 13990 8680 14230
rect 8770 13990 9010 14230
rect 9100 13990 9340 14230
rect 9430 13990 9670 14230
rect 9760 13990 10000 14230
rect 10090 13990 10330 14230
rect 10420 13990 10660 14230
rect 10750 13990 10990 14230
rect 11080 13990 11320 14230
rect 11410 13990 11650 14230
rect 11740 13990 11980 14230
rect 12070 13990 12310 14230
rect 12400 13990 12640 14230
rect 12730 13990 12970 14230
rect 13060 13990 13300 14230
rect 13390 13990 13630 14230
rect 13720 13990 13960 14230
rect 14050 13990 14290 14230
rect 14380 13990 14620 14230
rect 14710 13990 14950 14230
rect 15040 13990 15280 14230
rect 15370 13990 15610 14230
rect 15700 13990 15940 14230
rect 16030 13990 16270 14230
rect 16360 13990 16600 14230
rect 16690 13990 16930 14230
rect 17020 13990 17260 14230
rect 17350 13990 17590 14230
rect 17680 13990 17920 14230
rect 18010 13990 18250 14230
rect 18340 13990 18580 14230
rect 18670 13990 18910 14230
rect 19000 13990 19240 14230
rect 19330 13990 19570 14230
rect 7780 13660 8020 13900
rect 8110 13660 8350 13900
rect 8440 13660 8680 13900
rect 8770 13660 9010 13900
rect 9100 13660 9340 13900
rect 9430 13660 9670 13900
rect 9760 13660 10000 13900
rect 10090 13660 10330 13900
rect 10420 13660 10660 13900
rect 10750 13660 10990 13900
rect 11080 13660 11320 13900
rect 11410 13660 11650 13900
rect 11740 13660 11980 13900
rect 12070 13660 12310 13900
rect 12400 13660 12640 13900
rect 12730 13660 12970 13900
rect 13060 13660 13300 13900
rect 13390 13660 13630 13900
rect 13720 13660 13960 13900
rect 14050 13660 14290 13900
rect 14380 13660 14620 13900
rect 14710 13660 14950 13900
rect 15040 13660 15280 13900
rect 15370 13660 15610 13900
rect 15700 13660 15940 13900
rect 16030 13660 16270 13900
rect 16360 13660 16600 13900
rect 16690 13660 16930 13900
rect 17020 13660 17260 13900
rect 17350 13660 17590 13900
rect 17680 13660 17920 13900
rect 18010 13660 18250 13900
rect 18340 13660 18580 13900
rect 18670 13660 18910 13900
rect 19000 13660 19240 13900
rect 19330 13660 19570 13900
rect 7780 13330 8020 13570
rect 8110 13330 8350 13570
rect 8440 13330 8680 13570
rect 8770 13330 9010 13570
rect 9100 13330 9340 13570
rect 9430 13330 9670 13570
rect 9760 13330 10000 13570
rect 10090 13330 10330 13570
rect 10420 13330 10660 13570
rect 10750 13330 10990 13570
rect 11080 13330 11320 13570
rect 11410 13330 11650 13570
rect 11740 13330 11980 13570
rect 12070 13330 12310 13570
rect 12400 13330 12640 13570
rect 12730 13330 12970 13570
rect 13060 13330 13300 13570
rect 13390 13330 13630 13570
rect 13720 13330 13960 13570
rect 14050 13330 14290 13570
rect 14380 13330 14620 13570
rect 14710 13330 14950 13570
rect 15040 13330 15280 13570
rect 15370 13330 15610 13570
rect 15700 13330 15940 13570
rect 16030 13330 16270 13570
rect 16360 13330 16600 13570
rect 16690 13330 16930 13570
rect 17020 13330 17260 13570
rect 17350 13330 17590 13570
rect 17680 13330 17920 13570
rect 18010 13330 18250 13570
rect 18340 13330 18580 13570
rect 18670 13330 18910 13570
rect 19000 13330 19240 13570
rect 19330 13330 19570 13570
rect 7780 13000 8020 13240
rect 8110 13000 8350 13240
rect 8440 13000 8680 13240
rect 8770 13000 9010 13240
rect 9100 13000 9340 13240
rect 9430 13000 9670 13240
rect 9760 13000 10000 13240
rect 10090 13000 10330 13240
rect 10420 13000 10660 13240
rect 10750 13000 10990 13240
rect 11080 13000 11320 13240
rect 11410 13000 11650 13240
rect 11740 13000 11980 13240
rect 12070 13000 12310 13240
rect 12400 13000 12640 13240
rect 12730 13000 12970 13240
rect 13060 13000 13300 13240
rect 13390 13000 13630 13240
rect 13720 13000 13960 13240
rect 14050 13000 14290 13240
rect 14380 13000 14620 13240
rect 14710 13000 14950 13240
rect 15040 13000 15280 13240
rect 15370 13000 15610 13240
rect 15700 13000 15940 13240
rect 16030 13000 16270 13240
rect 16360 13000 16600 13240
rect 16690 13000 16930 13240
rect 17020 13000 17260 13240
rect 17350 13000 17590 13240
rect 17680 13000 17920 13240
rect 18010 13000 18250 13240
rect 18340 13000 18580 13240
rect 18670 13000 18910 13240
rect 19000 13000 19240 13240
rect 19330 13000 19570 13240
rect 7780 12670 8020 12910
rect 8110 12670 8350 12910
rect 8440 12670 8680 12910
rect 8770 12670 9010 12910
rect 9100 12670 9340 12910
rect 9430 12670 9670 12910
rect 9760 12670 10000 12910
rect 10090 12670 10330 12910
rect 10420 12670 10660 12910
rect 10750 12670 10990 12910
rect 11080 12670 11320 12910
rect 11410 12670 11650 12910
rect 11740 12670 11980 12910
rect 12070 12670 12310 12910
rect 12400 12670 12640 12910
rect 12730 12670 12970 12910
rect 13060 12670 13300 12910
rect 13390 12670 13630 12910
rect 13720 12670 13960 12910
rect 14050 12670 14290 12910
rect 14380 12670 14620 12910
rect 14710 12670 14950 12910
rect 15040 12670 15280 12910
rect 15370 12670 15610 12910
rect 15700 12670 15940 12910
rect 16030 12670 16270 12910
rect 16360 12670 16600 12910
rect 16690 12670 16930 12910
rect 17020 12670 17260 12910
rect 17350 12670 17590 12910
rect 17680 12670 17920 12910
rect 18010 12670 18250 12910
rect 18340 12670 18580 12910
rect 18670 12670 18910 12910
rect 19000 12670 19240 12910
rect 19330 12670 19570 12910
rect 7780 12340 8020 12580
rect 8110 12340 8350 12580
rect 8440 12340 8680 12580
rect 8770 12340 9010 12580
rect 9100 12340 9340 12580
rect 9430 12340 9670 12580
rect 9760 12340 10000 12580
rect 10090 12340 10330 12580
rect 10420 12340 10660 12580
rect 10750 12340 10990 12580
rect 11080 12340 11320 12580
rect 11410 12340 11650 12580
rect 11740 12340 11980 12580
rect 12070 12340 12310 12580
rect 12400 12340 12640 12580
rect 12730 12340 12970 12580
rect 13060 12340 13300 12580
rect 13390 12340 13630 12580
rect 13720 12340 13960 12580
rect 14050 12340 14290 12580
rect 14380 12340 14620 12580
rect 14710 12340 14950 12580
rect 15040 12340 15280 12580
rect 15370 12340 15610 12580
rect 15700 12340 15940 12580
rect 16030 12340 16270 12580
rect 16360 12340 16600 12580
rect 16690 12340 16930 12580
rect 17020 12340 17260 12580
rect 17350 12340 17590 12580
rect 17680 12340 17920 12580
rect 18010 12340 18250 12580
rect 18340 12340 18580 12580
rect 18670 12340 18910 12580
rect 19000 12340 19240 12580
rect 19330 12340 19570 12580
rect 7780 12010 8020 12250
rect 8110 12010 8350 12250
rect 8440 12010 8680 12250
rect 8770 12010 9010 12250
rect 9100 12010 9340 12250
rect 9430 12010 9670 12250
rect 9760 12010 10000 12250
rect 10090 12010 10330 12250
rect 10420 12010 10660 12250
rect 10750 12010 10990 12250
rect 11080 12010 11320 12250
rect 11410 12010 11650 12250
rect 11740 12010 11980 12250
rect 12070 12010 12310 12250
rect 12400 12010 12640 12250
rect 12730 12010 12970 12250
rect 13060 12010 13300 12250
rect 13390 12010 13630 12250
rect 13720 12010 13960 12250
rect 14050 12010 14290 12250
rect 14380 12010 14620 12250
rect 14710 12010 14950 12250
rect 15040 12010 15280 12250
rect 15370 12010 15610 12250
rect 15700 12010 15940 12250
rect 16030 12010 16270 12250
rect 16360 12010 16600 12250
rect 16690 12010 16930 12250
rect 17020 12010 17260 12250
rect 17350 12010 17590 12250
rect 17680 12010 17920 12250
rect 18010 12010 18250 12250
rect 18340 12010 18580 12250
rect 18670 12010 18910 12250
rect 19000 12010 19240 12250
rect 19330 12010 19570 12250
rect 7780 11680 8020 11920
rect 8110 11680 8350 11920
rect 8440 11680 8680 11920
rect 8770 11680 9010 11920
rect 9100 11680 9340 11920
rect 9430 11680 9670 11920
rect 9760 11680 10000 11920
rect 10090 11680 10330 11920
rect 10420 11680 10660 11920
rect 10750 11680 10990 11920
rect 11080 11680 11320 11920
rect 11410 11680 11650 11920
rect 11740 11680 11980 11920
rect 12070 11680 12310 11920
rect 12400 11680 12640 11920
rect 12730 11680 12970 11920
rect 13060 11680 13300 11920
rect 13390 11680 13630 11920
rect 13720 11680 13960 11920
rect 14050 11680 14290 11920
rect 14380 11680 14620 11920
rect 14710 11680 14950 11920
rect 15040 11680 15280 11920
rect 15370 11680 15610 11920
rect 15700 11680 15940 11920
rect 16030 11680 16270 11920
rect 16360 11680 16600 11920
rect 16690 11680 16930 11920
rect 17020 11680 17260 11920
rect 17350 11680 17590 11920
rect 17680 11680 17920 11920
rect 18010 11680 18250 11920
rect 18340 11680 18580 11920
rect 18670 11680 18910 11920
rect 19000 11680 19240 11920
rect 19330 11680 19570 11920
rect 7780 11350 8020 11590
rect 8110 11350 8350 11590
rect 8440 11350 8680 11590
rect 8770 11350 9010 11590
rect 9100 11350 9340 11590
rect 9430 11350 9670 11590
rect 9760 11350 10000 11590
rect 10090 11350 10330 11590
rect 10420 11350 10660 11590
rect 10750 11350 10990 11590
rect 11080 11350 11320 11590
rect 11410 11350 11650 11590
rect 11740 11350 11980 11590
rect 12070 11350 12310 11590
rect 12400 11350 12640 11590
rect 12730 11350 12970 11590
rect 13060 11350 13300 11590
rect 13390 11350 13630 11590
rect 13720 11350 13960 11590
rect 14050 11350 14290 11590
rect 14380 11350 14620 11590
rect 14710 11350 14950 11590
rect 15040 11350 15280 11590
rect 15370 11350 15610 11590
rect 15700 11350 15940 11590
rect 16030 11350 16270 11590
rect 16360 11350 16600 11590
rect 16690 11350 16930 11590
rect 17020 11350 17260 11590
rect 17350 11350 17590 11590
rect 17680 11350 17920 11590
rect 18010 11350 18250 11590
rect 18340 11350 18580 11590
rect 18670 11350 18910 11590
rect 19000 11350 19240 11590
rect 19330 11350 19570 11590
rect 7780 11020 8020 11260
rect 8110 11020 8350 11260
rect 8440 11020 8680 11260
rect 8770 11020 9010 11260
rect 9100 11020 9340 11260
rect 9430 11020 9670 11260
rect 9760 11020 10000 11260
rect 10090 11020 10330 11260
rect 10420 11020 10660 11260
rect 10750 11020 10990 11260
rect 11080 11020 11320 11260
rect 11410 11020 11650 11260
rect 11740 11020 11980 11260
rect 12070 11020 12310 11260
rect 12400 11020 12640 11260
rect 12730 11020 12970 11260
rect 13060 11020 13300 11260
rect 13390 11020 13630 11260
rect 13720 11020 13960 11260
rect 14050 11020 14290 11260
rect 14380 11020 14620 11260
rect 14710 11020 14950 11260
rect 15040 11020 15280 11260
rect 15370 11020 15610 11260
rect 15700 11020 15940 11260
rect 16030 11020 16270 11260
rect 16360 11020 16600 11260
rect 16690 11020 16930 11260
rect 17020 11020 17260 11260
rect 17350 11020 17590 11260
rect 17680 11020 17920 11260
rect 18010 11020 18250 11260
rect 18340 11020 18580 11260
rect 18670 11020 18910 11260
rect 19000 11020 19240 11260
rect 19330 11020 19570 11260
rect 7780 10690 8020 10930
rect 8110 10690 8350 10930
rect 8440 10690 8680 10930
rect 8770 10690 9010 10930
rect 9100 10690 9340 10930
rect 9430 10690 9670 10930
rect 9760 10690 10000 10930
rect 10090 10690 10330 10930
rect 10420 10690 10660 10930
rect 10750 10690 10990 10930
rect 11080 10690 11320 10930
rect 11410 10690 11650 10930
rect 11740 10690 11980 10930
rect 12070 10690 12310 10930
rect 12400 10690 12640 10930
rect 12730 10690 12970 10930
rect 13060 10690 13300 10930
rect 13390 10690 13630 10930
rect 13720 10690 13960 10930
rect 14050 10690 14290 10930
rect 14380 10690 14620 10930
rect 14710 10690 14950 10930
rect 15040 10690 15280 10930
rect 15370 10690 15610 10930
rect 15700 10690 15940 10930
rect 16030 10690 16270 10930
rect 16360 10690 16600 10930
rect 16690 10690 16930 10930
rect 17020 10690 17260 10930
rect 17350 10690 17590 10930
rect 17680 10690 17920 10930
rect 18010 10690 18250 10930
rect 18340 10690 18580 10930
rect 18670 10690 18910 10930
rect 19000 10690 19240 10930
rect 19330 10690 19570 10930
rect 7780 10360 8020 10600
rect 8110 10360 8350 10600
rect 8440 10360 8680 10600
rect 8770 10360 9010 10600
rect 9100 10360 9340 10600
rect 9430 10360 9670 10600
rect 9760 10360 10000 10600
rect 10090 10360 10330 10600
rect 10420 10360 10660 10600
rect 10750 10360 10990 10600
rect 11080 10360 11320 10600
rect 11410 10360 11650 10600
rect 11740 10360 11980 10600
rect 12070 10360 12310 10600
rect 12400 10360 12640 10600
rect 12730 10360 12970 10600
rect 13060 10360 13300 10600
rect 13390 10360 13630 10600
rect 13720 10360 13960 10600
rect 14050 10360 14290 10600
rect 14380 10360 14620 10600
rect 14710 10360 14950 10600
rect 15040 10360 15280 10600
rect 15370 10360 15610 10600
rect 15700 10360 15940 10600
rect 16030 10360 16270 10600
rect 16360 10360 16600 10600
rect 16690 10360 16930 10600
rect 17020 10360 17260 10600
rect 17350 10360 17590 10600
rect 17680 10360 17920 10600
rect 18010 10360 18250 10600
rect 18340 10360 18580 10600
rect 18670 10360 18910 10600
rect 19000 10360 19240 10600
rect 19330 10360 19570 10600
rect 7780 10030 8020 10270
rect 8110 10030 8350 10270
rect 8440 10030 8680 10270
rect 8770 10030 9010 10270
rect 9100 10030 9340 10270
rect 9430 10030 9670 10270
rect 9760 10030 10000 10270
rect 10090 10030 10330 10270
rect 10420 10030 10660 10270
rect 10750 10030 10990 10270
rect 11080 10030 11320 10270
rect 11410 10030 11650 10270
rect 11740 10030 11980 10270
rect 12070 10030 12310 10270
rect 12400 10030 12640 10270
rect 12730 10030 12970 10270
rect 13060 10030 13300 10270
rect 13390 10030 13630 10270
rect 13720 10030 13960 10270
rect 14050 10030 14290 10270
rect 14380 10030 14620 10270
rect 14710 10030 14950 10270
rect 15040 10030 15280 10270
rect 15370 10030 15610 10270
rect 15700 10030 15940 10270
rect 16030 10030 16270 10270
rect 16360 10030 16600 10270
rect 16690 10030 16930 10270
rect 17020 10030 17260 10270
rect 17350 10030 17590 10270
rect 17680 10030 17920 10270
rect 18010 10030 18250 10270
rect 18340 10030 18580 10270
rect 18670 10030 18910 10270
rect 19000 10030 19240 10270
rect 19330 10030 19570 10270
rect 7780 9700 8020 9940
rect 8110 9700 8350 9940
rect 8440 9700 8680 9940
rect 8770 9700 9010 9940
rect 9100 9700 9340 9940
rect 9430 9700 9670 9940
rect 9760 9700 10000 9940
rect 10090 9700 10330 9940
rect 10420 9700 10660 9940
rect 10750 9700 10990 9940
rect 11080 9700 11320 9940
rect 11410 9700 11650 9940
rect 11740 9700 11980 9940
rect 12070 9700 12310 9940
rect 12400 9700 12640 9940
rect 12730 9700 12970 9940
rect 13060 9700 13300 9940
rect 13390 9700 13630 9940
rect 13720 9700 13960 9940
rect 14050 9700 14290 9940
rect 14380 9700 14620 9940
rect 14710 9700 14950 9940
rect 15040 9700 15280 9940
rect 15370 9700 15610 9940
rect 15700 9700 15940 9940
rect 16030 9700 16270 9940
rect 16360 9700 16600 9940
rect 16690 9700 16930 9940
rect 17020 9700 17260 9940
rect 17350 9700 17590 9940
rect 17680 9700 17920 9940
rect 18010 9700 18250 9940
rect 18340 9700 18580 9940
rect 18670 9700 18910 9940
rect 19000 9700 19240 9940
rect 19330 9700 19570 9940
rect 7780 9370 8020 9610
rect 8110 9370 8350 9610
rect 8440 9370 8680 9610
rect 8770 9370 9010 9610
rect 9100 9370 9340 9610
rect 9430 9370 9670 9610
rect 9760 9370 10000 9610
rect 10090 9370 10330 9610
rect 10420 9370 10660 9610
rect 10750 9370 10990 9610
rect 11080 9370 11320 9610
rect 11410 9370 11650 9610
rect 11740 9370 11980 9610
rect 12070 9370 12310 9610
rect 12400 9370 12640 9610
rect 12730 9370 12970 9610
rect 13060 9370 13300 9610
rect 13390 9370 13630 9610
rect 13720 9370 13960 9610
rect 14050 9370 14290 9610
rect 14380 9370 14620 9610
rect 14710 9370 14950 9610
rect 15040 9370 15280 9610
rect 15370 9370 15610 9610
rect 15700 9370 15940 9610
rect 16030 9370 16270 9610
rect 16360 9370 16600 9610
rect 16690 9370 16930 9610
rect 17020 9370 17260 9610
rect 17350 9370 17590 9610
rect 17680 9370 17920 9610
rect 18010 9370 18250 9610
rect 18340 9370 18580 9610
rect 18670 9370 18910 9610
rect 19000 9370 19240 9610
rect 19330 9370 19570 9610
rect 7780 9040 8020 9280
rect 8110 9040 8350 9280
rect 8440 9040 8680 9280
rect 8770 9040 9010 9280
rect 9100 9040 9340 9280
rect 9430 9040 9670 9280
rect 9760 9040 10000 9280
rect 10090 9040 10330 9280
rect 10420 9040 10660 9280
rect 10750 9040 10990 9280
rect 11080 9040 11320 9280
rect 11410 9040 11650 9280
rect 11740 9040 11980 9280
rect 12070 9040 12310 9280
rect 12400 9040 12640 9280
rect 12730 9040 12970 9280
rect 13060 9040 13300 9280
rect 13390 9040 13630 9280
rect 13720 9040 13960 9280
rect 14050 9040 14290 9280
rect 14380 9040 14620 9280
rect 14710 9040 14950 9280
rect 15040 9040 15280 9280
rect 15370 9040 15610 9280
rect 15700 9040 15940 9280
rect 16030 9040 16270 9280
rect 16360 9040 16600 9280
rect 16690 9040 16930 9280
rect 17020 9040 17260 9280
rect 17350 9040 17590 9280
rect 17680 9040 17920 9280
rect 18010 9040 18250 9280
rect 18340 9040 18580 9280
rect 18670 9040 18910 9280
rect 19000 9040 19240 9280
rect 19330 9040 19570 9280
rect 31180 7590 31420 7830
rect 31510 7590 31750 7830
rect 31840 7590 32080 7830
rect 32170 7590 32410 7830
rect 32500 7590 32740 7830
rect 32830 7590 33070 7830
rect 33160 7590 33400 7830
rect 33490 7590 33730 7830
rect 33820 7590 34060 7830
rect 34150 7590 34390 7830
rect 34480 7590 34720 7830
rect 34810 7590 35050 7830
rect 35140 7590 35380 7830
rect 35470 7590 35710 7830
rect 35800 7590 36040 7830
rect 36130 7590 36370 7830
rect 36460 7590 36700 7830
rect 36790 7590 37030 7830
rect 37120 7590 37360 7830
rect 37450 7590 37690 7830
rect 31180 7260 31420 7500
rect 31510 7260 31750 7500
rect 31840 7260 32080 7500
rect 32170 7260 32410 7500
rect 32500 7260 32740 7500
rect 32830 7260 33070 7500
rect 33160 7260 33400 7500
rect 33490 7260 33730 7500
rect 33820 7260 34060 7500
rect 34150 7260 34390 7500
rect 34480 7260 34720 7500
rect 34810 7260 35050 7500
rect 35140 7260 35380 7500
rect 35470 7260 35710 7500
rect 35800 7260 36040 7500
rect 36130 7260 36370 7500
rect 36460 7260 36700 7500
rect 36790 7260 37030 7500
rect 37120 7260 37360 7500
rect 37450 7260 37690 7500
rect 31180 6930 31420 7170
rect 31510 6930 31750 7170
rect 31840 6930 32080 7170
rect 32170 6930 32410 7170
rect 32500 6930 32740 7170
rect 32830 6930 33070 7170
rect 33160 6930 33400 7170
rect 33490 6930 33730 7170
rect 33820 6930 34060 7170
rect 34150 6930 34390 7170
rect 34480 6930 34720 7170
rect 34810 6930 35050 7170
rect 35140 6930 35380 7170
rect 35470 6930 35710 7170
rect 35800 6930 36040 7170
rect 36130 6930 36370 7170
rect 36460 6930 36700 7170
rect 36790 6930 37030 7170
rect 37120 6930 37360 7170
rect 37450 6930 37690 7170
rect 31180 6600 31420 6840
rect 31510 6600 31750 6840
rect 31840 6600 32080 6840
rect 32170 6600 32410 6840
rect 32500 6600 32740 6840
rect 32830 6600 33070 6840
rect 33160 6600 33400 6840
rect 33490 6600 33730 6840
rect 33820 6600 34060 6840
rect 34150 6600 34390 6840
rect 34480 6600 34720 6840
rect 34810 6600 35050 6840
rect 35140 6600 35380 6840
rect 35470 6600 35710 6840
rect 35800 6600 36040 6840
rect 36130 6600 36370 6840
rect 36460 6600 36700 6840
rect 36790 6600 37030 6840
rect 37120 6600 37360 6840
rect 37450 6600 37690 6840
rect 31180 6270 31420 6510
rect 31510 6270 31750 6510
rect 31840 6270 32080 6510
rect 32170 6270 32410 6510
rect 32500 6270 32740 6510
rect 32830 6270 33070 6510
rect 33160 6270 33400 6510
rect 33490 6270 33730 6510
rect 33820 6270 34060 6510
rect 34150 6270 34390 6510
rect 34480 6270 34720 6510
rect 34810 6270 35050 6510
rect 35140 6270 35380 6510
rect 35470 6270 35710 6510
rect 35800 6270 36040 6510
rect 36130 6270 36370 6510
rect 36460 6270 36700 6510
rect 36790 6270 37030 6510
rect 37120 6270 37360 6510
rect 37450 6270 37690 6510
rect 31180 5940 31420 6180
rect 31510 5940 31750 6180
rect 31840 5940 32080 6180
rect 32170 5940 32410 6180
rect 32500 5940 32740 6180
rect 32830 5940 33070 6180
rect 33160 5940 33400 6180
rect 33490 5940 33730 6180
rect 33820 5940 34060 6180
rect 34150 5940 34390 6180
rect 34480 5940 34720 6180
rect 34810 5940 35050 6180
rect 35140 5940 35380 6180
rect 35470 5940 35710 6180
rect 35800 5940 36040 6180
rect 36130 5940 36370 6180
rect 36460 5940 36700 6180
rect 36790 5940 37030 6180
rect 37120 5940 37360 6180
rect 37450 5940 37690 6180
rect 31180 5610 31420 5850
rect 31510 5610 31750 5850
rect 31840 5610 32080 5850
rect 32170 5610 32410 5850
rect 32500 5610 32740 5850
rect 32830 5610 33070 5850
rect 33160 5610 33400 5850
rect 33490 5610 33730 5850
rect 33820 5610 34060 5850
rect 34150 5610 34390 5850
rect 34480 5610 34720 5850
rect 34810 5610 35050 5850
rect 35140 5610 35380 5850
rect 35470 5610 35710 5850
rect 35800 5610 36040 5850
rect 36130 5610 36370 5850
rect 36460 5610 36700 5850
rect 36790 5610 37030 5850
rect 37120 5610 37360 5850
rect 37450 5610 37690 5850
rect 31180 5280 31420 5520
rect 31510 5280 31750 5520
rect 31840 5280 32080 5520
rect 32170 5280 32410 5520
rect 32500 5280 32740 5520
rect 32830 5280 33070 5520
rect 33160 5280 33400 5520
rect 33490 5280 33730 5520
rect 33820 5280 34060 5520
rect 34150 5280 34390 5520
rect 34480 5280 34720 5520
rect 34810 5280 35050 5520
rect 35140 5280 35380 5520
rect 35470 5280 35710 5520
rect 35800 5280 36040 5520
rect 36130 5280 36370 5520
rect 36460 5280 36700 5520
rect 36790 5280 37030 5520
rect 37120 5280 37360 5520
rect 37450 5280 37690 5520
rect 31180 4950 31420 5190
rect 31510 4950 31750 5190
rect 31840 4950 32080 5190
rect 32170 4950 32410 5190
rect 32500 4950 32740 5190
rect 32830 4950 33070 5190
rect 33160 4950 33400 5190
rect 33490 4950 33730 5190
rect 33820 4950 34060 5190
rect 34150 4950 34390 5190
rect 34480 4950 34720 5190
rect 34810 4950 35050 5190
rect 35140 4950 35380 5190
rect 35470 4950 35710 5190
rect 35800 4950 36040 5190
rect 36130 4950 36370 5190
rect 36460 4950 36700 5190
rect 36790 4950 37030 5190
rect 37120 4950 37360 5190
rect 37450 4950 37690 5190
rect 31180 4620 31420 4860
rect 31510 4620 31750 4860
rect 31840 4620 32080 4860
rect 32170 4620 32410 4860
rect 32500 4620 32740 4860
rect 32830 4620 33070 4860
rect 33160 4620 33400 4860
rect 33490 4620 33730 4860
rect 33820 4620 34060 4860
rect 34150 4620 34390 4860
rect 34480 4620 34720 4860
rect 34810 4620 35050 4860
rect 35140 4620 35380 4860
rect 35470 4620 35710 4860
rect 35800 4620 36040 4860
rect 36130 4620 36370 4860
rect 36460 4620 36700 4860
rect 36790 4620 37030 4860
rect 37120 4620 37360 4860
rect 37450 4620 37690 4860
rect 31180 4290 31420 4530
rect 31510 4290 31750 4530
rect 31840 4290 32080 4530
rect 32170 4290 32410 4530
rect 32500 4290 32740 4530
rect 32830 4290 33070 4530
rect 33160 4290 33400 4530
rect 33490 4290 33730 4530
rect 33820 4290 34060 4530
rect 34150 4290 34390 4530
rect 34480 4290 34720 4530
rect 34810 4290 35050 4530
rect 35140 4290 35380 4530
rect 35470 4290 35710 4530
rect 35800 4290 36040 4530
rect 36130 4290 36370 4530
rect 36460 4290 36700 4530
rect 36790 4290 37030 4530
rect 37120 4290 37360 4530
rect 37450 4290 37690 4530
rect 31180 3960 31420 4200
rect 31510 3960 31750 4200
rect 31840 3960 32080 4200
rect 32170 3960 32410 4200
rect 32500 3960 32740 4200
rect 32830 3960 33070 4200
rect 33160 3960 33400 4200
rect 33490 3960 33730 4200
rect 33820 3960 34060 4200
rect 34150 3960 34390 4200
rect 34480 3960 34720 4200
rect 34810 3960 35050 4200
rect 35140 3960 35380 4200
rect 35470 3960 35710 4200
rect 35800 3960 36040 4200
rect 36130 3960 36370 4200
rect 36460 3960 36700 4200
rect 36790 3960 37030 4200
rect 37120 3960 37360 4200
rect 37450 3960 37690 4200
rect 31180 3630 31420 3870
rect 31510 3630 31750 3870
rect 31840 3630 32080 3870
rect 32170 3630 32410 3870
rect 32500 3630 32740 3870
rect 32830 3630 33070 3870
rect 33160 3630 33400 3870
rect 33490 3630 33730 3870
rect 33820 3630 34060 3870
rect 34150 3630 34390 3870
rect 34480 3630 34720 3870
rect 34810 3630 35050 3870
rect 35140 3630 35380 3870
rect 35470 3630 35710 3870
rect 35800 3630 36040 3870
rect 36130 3630 36370 3870
rect 36460 3630 36700 3870
rect 36790 3630 37030 3870
rect 37120 3630 37360 3870
rect 37450 3630 37690 3870
rect 31180 3300 31420 3540
rect 31510 3300 31750 3540
rect 31840 3300 32080 3540
rect 32170 3300 32410 3540
rect 32500 3300 32740 3540
rect 32830 3300 33070 3540
rect 33160 3300 33400 3540
rect 33490 3300 33730 3540
rect 33820 3300 34060 3540
rect 34150 3300 34390 3540
rect 34480 3300 34720 3540
rect 34810 3300 35050 3540
rect 35140 3300 35380 3540
rect 35470 3300 35710 3540
rect 35800 3300 36040 3540
rect 36130 3300 36370 3540
rect 36460 3300 36700 3540
rect 36790 3300 37030 3540
rect 37120 3300 37360 3540
rect 37450 3300 37690 3540
rect 31180 2970 31420 3210
rect 31510 2970 31750 3210
rect 31840 2970 32080 3210
rect 32170 2970 32410 3210
rect 32500 2970 32740 3210
rect 32830 2970 33070 3210
rect 33160 2970 33400 3210
rect 33490 2970 33730 3210
rect 33820 2970 34060 3210
rect 34150 2970 34390 3210
rect 34480 2970 34720 3210
rect 34810 2970 35050 3210
rect 35140 2970 35380 3210
rect 35470 2970 35710 3210
rect 35800 2970 36040 3210
rect 36130 2970 36370 3210
rect 36460 2970 36700 3210
rect 36790 2970 37030 3210
rect 37120 2970 37360 3210
rect 37450 2970 37690 3210
rect 31180 2640 31420 2880
rect 31510 2640 31750 2880
rect 31840 2640 32080 2880
rect 32170 2640 32410 2880
rect 32500 2640 32740 2880
rect 32830 2640 33070 2880
rect 33160 2640 33400 2880
rect 33490 2640 33730 2880
rect 33820 2640 34060 2880
rect 34150 2640 34390 2880
rect 34480 2640 34720 2880
rect 34810 2640 35050 2880
rect 35140 2640 35380 2880
rect 35470 2640 35710 2880
rect 35800 2640 36040 2880
rect 36130 2640 36370 2880
rect 36460 2640 36700 2880
rect 36790 2640 37030 2880
rect 37120 2640 37360 2880
rect 37450 2640 37690 2880
rect 31180 2310 31420 2550
rect 31510 2310 31750 2550
rect 31840 2310 32080 2550
rect 32170 2310 32410 2550
rect 32500 2310 32740 2550
rect 32830 2310 33070 2550
rect 33160 2310 33400 2550
rect 33490 2310 33730 2550
rect 33820 2310 34060 2550
rect 34150 2310 34390 2550
rect 34480 2310 34720 2550
rect 34810 2310 35050 2550
rect 35140 2310 35380 2550
rect 35470 2310 35710 2550
rect 35800 2310 36040 2550
rect 36130 2310 36370 2550
rect 36460 2310 36700 2550
rect 36790 2310 37030 2550
rect 37120 2310 37360 2550
rect 37450 2310 37690 2550
rect 31180 1980 31420 2220
rect 31510 1980 31750 2220
rect 31840 1980 32080 2220
rect 32170 1980 32410 2220
rect 32500 1980 32740 2220
rect 32830 1980 33070 2220
rect 33160 1980 33400 2220
rect 33490 1980 33730 2220
rect 33820 1980 34060 2220
rect 34150 1980 34390 2220
rect 34480 1980 34720 2220
rect 34810 1980 35050 2220
rect 35140 1980 35380 2220
rect 35470 1980 35710 2220
rect 35800 1980 36040 2220
rect 36130 1980 36370 2220
rect 36460 1980 36700 2220
rect 36790 1980 37030 2220
rect 37120 1980 37360 2220
rect 37450 1980 37690 2220
rect 31180 1650 31420 1890
rect 31510 1650 31750 1890
rect 31840 1650 32080 1890
rect 32170 1650 32410 1890
rect 32500 1650 32740 1890
rect 32830 1650 33070 1890
rect 33160 1650 33400 1890
rect 33490 1650 33730 1890
rect 33820 1650 34060 1890
rect 34150 1650 34390 1890
rect 34480 1650 34720 1890
rect 34810 1650 35050 1890
rect 35140 1650 35380 1890
rect 35470 1650 35710 1890
rect 35800 1650 36040 1890
rect 36130 1650 36370 1890
rect 36460 1650 36700 1890
rect 36790 1650 37030 1890
rect 37120 1650 37360 1890
rect 37450 1650 37690 1890
rect 31180 1320 31420 1560
rect 31510 1320 31750 1560
rect 31840 1320 32080 1560
rect 32170 1320 32410 1560
rect 32500 1320 32740 1560
rect 32830 1320 33070 1560
rect 33160 1320 33400 1560
rect 33490 1320 33730 1560
rect 33820 1320 34060 1560
rect 34150 1320 34390 1560
rect 34480 1320 34720 1560
rect 34810 1320 35050 1560
rect 35140 1320 35380 1560
rect 35470 1320 35710 1560
rect 35800 1320 36040 1560
rect 36130 1320 36370 1560
rect 36460 1320 36700 1560
rect 36790 1320 37030 1560
rect 37120 1320 37360 1560
rect 37450 1320 37690 1560
rect 31180 -10 31420 230
rect 31510 -10 31750 230
rect 31840 -10 32080 230
rect 32170 -10 32410 230
rect 32500 -10 32740 230
rect 32830 -10 33070 230
rect 33160 -10 33400 230
rect 33490 -10 33730 230
rect 33820 -10 34060 230
rect 34150 -10 34390 230
rect 34480 -10 34720 230
rect 34810 -10 35050 230
rect 35140 -10 35380 230
rect 35470 -10 35710 230
rect 35800 -10 36040 230
rect 36130 -10 36370 230
rect 36460 -10 36700 230
rect 36790 -10 37030 230
rect 37120 -10 37360 230
rect 37450 -10 37690 230
rect 31180 -340 31420 -100
rect 31510 -340 31750 -100
rect 31840 -340 32080 -100
rect 32170 -340 32410 -100
rect 32500 -340 32740 -100
rect 32830 -340 33070 -100
rect 33160 -340 33400 -100
rect 33490 -340 33730 -100
rect 33820 -340 34060 -100
rect 34150 -340 34390 -100
rect 34480 -340 34720 -100
rect 34810 -340 35050 -100
rect 35140 -340 35380 -100
rect 35470 -340 35710 -100
rect 35800 -340 36040 -100
rect 36130 -340 36370 -100
rect 36460 -340 36700 -100
rect 36790 -340 37030 -100
rect 37120 -340 37360 -100
rect 37450 -340 37690 -100
rect 31180 -670 31420 -430
rect 31510 -670 31750 -430
rect 31840 -670 32080 -430
rect 32170 -670 32410 -430
rect 32500 -670 32740 -430
rect 32830 -670 33070 -430
rect 33160 -670 33400 -430
rect 33490 -670 33730 -430
rect 33820 -670 34060 -430
rect 34150 -670 34390 -430
rect 34480 -670 34720 -430
rect 34810 -670 35050 -430
rect 35140 -670 35380 -430
rect 35470 -670 35710 -430
rect 35800 -670 36040 -430
rect 36130 -670 36370 -430
rect 36460 -670 36700 -430
rect 36790 -670 37030 -430
rect 37120 -670 37360 -430
rect 37450 -670 37690 -430
rect 31180 -1000 31420 -760
rect 31510 -1000 31750 -760
rect 31840 -1000 32080 -760
rect 32170 -1000 32410 -760
rect 32500 -1000 32740 -760
rect 32830 -1000 33070 -760
rect 33160 -1000 33400 -760
rect 33490 -1000 33730 -760
rect 33820 -1000 34060 -760
rect 34150 -1000 34390 -760
rect 34480 -1000 34720 -760
rect 34810 -1000 35050 -760
rect 35140 -1000 35380 -760
rect 35470 -1000 35710 -760
rect 35800 -1000 36040 -760
rect 36130 -1000 36370 -760
rect 36460 -1000 36700 -760
rect 36790 -1000 37030 -760
rect 37120 -1000 37360 -760
rect 37450 -1000 37690 -760
rect 31180 -1330 31420 -1090
rect 31510 -1330 31750 -1090
rect 31840 -1330 32080 -1090
rect 32170 -1330 32410 -1090
rect 32500 -1330 32740 -1090
rect 32830 -1330 33070 -1090
rect 33160 -1330 33400 -1090
rect 33490 -1330 33730 -1090
rect 33820 -1330 34060 -1090
rect 34150 -1330 34390 -1090
rect 34480 -1330 34720 -1090
rect 34810 -1330 35050 -1090
rect 35140 -1330 35380 -1090
rect 35470 -1330 35710 -1090
rect 35800 -1330 36040 -1090
rect 36130 -1330 36370 -1090
rect 36460 -1330 36700 -1090
rect 36790 -1330 37030 -1090
rect 37120 -1330 37360 -1090
rect 37450 -1330 37690 -1090
rect 31180 -1660 31420 -1420
rect 31510 -1660 31750 -1420
rect 31840 -1660 32080 -1420
rect 32170 -1660 32410 -1420
rect 32500 -1660 32740 -1420
rect 32830 -1660 33070 -1420
rect 33160 -1660 33400 -1420
rect 33490 -1660 33730 -1420
rect 33820 -1660 34060 -1420
rect 34150 -1660 34390 -1420
rect 34480 -1660 34720 -1420
rect 34810 -1660 35050 -1420
rect 35140 -1660 35380 -1420
rect 35470 -1660 35710 -1420
rect 35800 -1660 36040 -1420
rect 36130 -1660 36370 -1420
rect 36460 -1660 36700 -1420
rect 36790 -1660 37030 -1420
rect 37120 -1660 37360 -1420
rect 37450 -1660 37690 -1420
rect 31180 -1990 31420 -1750
rect 31510 -1990 31750 -1750
rect 31840 -1990 32080 -1750
rect 32170 -1990 32410 -1750
rect 32500 -1990 32740 -1750
rect 32830 -1990 33070 -1750
rect 33160 -1990 33400 -1750
rect 33490 -1990 33730 -1750
rect 33820 -1990 34060 -1750
rect 34150 -1990 34390 -1750
rect 34480 -1990 34720 -1750
rect 34810 -1990 35050 -1750
rect 35140 -1990 35380 -1750
rect 35470 -1990 35710 -1750
rect 35800 -1990 36040 -1750
rect 36130 -1990 36370 -1750
rect 36460 -1990 36700 -1750
rect 36790 -1990 37030 -1750
rect 37120 -1990 37360 -1750
rect 37450 -1990 37690 -1750
rect 31180 -2320 31420 -2080
rect 31510 -2320 31750 -2080
rect 31840 -2320 32080 -2080
rect 32170 -2320 32410 -2080
rect 32500 -2320 32740 -2080
rect 32830 -2320 33070 -2080
rect 33160 -2320 33400 -2080
rect 33490 -2320 33730 -2080
rect 33820 -2320 34060 -2080
rect 34150 -2320 34390 -2080
rect 34480 -2320 34720 -2080
rect 34810 -2320 35050 -2080
rect 35140 -2320 35380 -2080
rect 35470 -2320 35710 -2080
rect 35800 -2320 36040 -2080
rect 36130 -2320 36370 -2080
rect 36460 -2320 36700 -2080
rect 36790 -2320 37030 -2080
rect 37120 -2320 37360 -2080
rect 37450 -2320 37690 -2080
rect 31180 -2650 31420 -2410
rect 31510 -2650 31750 -2410
rect 31840 -2650 32080 -2410
rect 32170 -2650 32410 -2410
rect 32500 -2650 32740 -2410
rect 32830 -2650 33070 -2410
rect 33160 -2650 33400 -2410
rect 33490 -2650 33730 -2410
rect 33820 -2650 34060 -2410
rect 34150 -2650 34390 -2410
rect 34480 -2650 34720 -2410
rect 34810 -2650 35050 -2410
rect 35140 -2650 35380 -2410
rect 35470 -2650 35710 -2410
rect 35800 -2650 36040 -2410
rect 36130 -2650 36370 -2410
rect 36460 -2650 36700 -2410
rect 36790 -2650 37030 -2410
rect 37120 -2650 37360 -2410
rect 37450 -2650 37690 -2410
rect 31180 -2980 31420 -2740
rect 31510 -2980 31750 -2740
rect 31840 -2980 32080 -2740
rect 32170 -2980 32410 -2740
rect 32500 -2980 32740 -2740
rect 32830 -2980 33070 -2740
rect 33160 -2980 33400 -2740
rect 33490 -2980 33730 -2740
rect 33820 -2980 34060 -2740
rect 34150 -2980 34390 -2740
rect 34480 -2980 34720 -2740
rect 34810 -2980 35050 -2740
rect 35140 -2980 35380 -2740
rect 35470 -2980 35710 -2740
rect 35800 -2980 36040 -2740
rect 36130 -2980 36370 -2740
rect 36460 -2980 36700 -2740
rect 36790 -2980 37030 -2740
rect 37120 -2980 37360 -2740
rect 37450 -2980 37690 -2740
rect 31180 -3310 31420 -3070
rect 31510 -3310 31750 -3070
rect 31840 -3310 32080 -3070
rect 32170 -3310 32410 -3070
rect 32500 -3310 32740 -3070
rect 32830 -3310 33070 -3070
rect 33160 -3310 33400 -3070
rect 33490 -3310 33730 -3070
rect 33820 -3310 34060 -3070
rect 34150 -3310 34390 -3070
rect 34480 -3310 34720 -3070
rect 34810 -3310 35050 -3070
rect 35140 -3310 35380 -3070
rect 35470 -3310 35710 -3070
rect 35800 -3310 36040 -3070
rect 36130 -3310 36370 -3070
rect 36460 -3310 36700 -3070
rect 36790 -3310 37030 -3070
rect 37120 -3310 37360 -3070
rect 37450 -3310 37690 -3070
rect 31180 -3640 31420 -3400
rect 31510 -3640 31750 -3400
rect 31840 -3640 32080 -3400
rect 32170 -3640 32410 -3400
rect 32500 -3640 32740 -3400
rect 32830 -3640 33070 -3400
rect 33160 -3640 33400 -3400
rect 33490 -3640 33730 -3400
rect 33820 -3640 34060 -3400
rect 34150 -3640 34390 -3400
rect 34480 -3640 34720 -3400
rect 34810 -3640 35050 -3400
rect 35140 -3640 35380 -3400
rect 35470 -3640 35710 -3400
rect 35800 -3640 36040 -3400
rect 36130 -3640 36370 -3400
rect 36460 -3640 36700 -3400
rect 36790 -3640 37030 -3400
rect 37120 -3640 37360 -3400
rect 37450 -3640 37690 -3400
rect 31180 -3970 31420 -3730
rect 31510 -3970 31750 -3730
rect 31840 -3970 32080 -3730
rect 32170 -3970 32410 -3730
rect 32500 -3970 32740 -3730
rect 32830 -3970 33070 -3730
rect 33160 -3970 33400 -3730
rect 33490 -3970 33730 -3730
rect 33820 -3970 34060 -3730
rect 34150 -3970 34390 -3730
rect 34480 -3970 34720 -3730
rect 34810 -3970 35050 -3730
rect 35140 -3970 35380 -3730
rect 35470 -3970 35710 -3730
rect 35800 -3970 36040 -3730
rect 36130 -3970 36370 -3730
rect 36460 -3970 36700 -3730
rect 36790 -3970 37030 -3730
rect 37120 -3970 37360 -3730
rect 37450 -3970 37690 -3730
rect 31180 -4300 31420 -4060
rect 31510 -4300 31750 -4060
rect 31840 -4300 32080 -4060
rect 32170 -4300 32410 -4060
rect 32500 -4300 32740 -4060
rect 32830 -4300 33070 -4060
rect 33160 -4300 33400 -4060
rect 33490 -4300 33730 -4060
rect 33820 -4300 34060 -4060
rect 34150 -4300 34390 -4060
rect 34480 -4300 34720 -4060
rect 34810 -4300 35050 -4060
rect 35140 -4300 35380 -4060
rect 35470 -4300 35710 -4060
rect 35800 -4300 36040 -4060
rect 36130 -4300 36370 -4060
rect 36460 -4300 36700 -4060
rect 36790 -4300 37030 -4060
rect 37120 -4300 37360 -4060
rect 37450 -4300 37690 -4060
rect 31180 -4630 31420 -4390
rect 31510 -4630 31750 -4390
rect 31840 -4630 32080 -4390
rect 32170 -4630 32410 -4390
rect 32500 -4630 32740 -4390
rect 32830 -4630 33070 -4390
rect 33160 -4630 33400 -4390
rect 33490 -4630 33730 -4390
rect 33820 -4630 34060 -4390
rect 34150 -4630 34390 -4390
rect 34480 -4630 34720 -4390
rect 34810 -4630 35050 -4390
rect 35140 -4630 35380 -4390
rect 35470 -4630 35710 -4390
rect 35800 -4630 36040 -4390
rect 36130 -4630 36370 -4390
rect 36460 -4630 36700 -4390
rect 36790 -4630 37030 -4390
rect 37120 -4630 37360 -4390
rect 37450 -4630 37690 -4390
rect -1180 -5080 -940 -4840
rect -850 -5080 -610 -4840
rect -520 -5080 -280 -4840
rect -190 -5080 50 -4840
rect -1180 -5410 -940 -5170
rect -850 -5410 -610 -5170
rect -520 -5410 -280 -5170
rect -190 -5410 50 -5170
rect -1180 -5740 -940 -5500
rect -850 -5740 -610 -5500
rect -520 -5740 -280 -5500
rect -190 -5740 50 -5500
rect -1180 -6070 -940 -5830
rect -850 -6070 -610 -5830
rect -520 -6070 -280 -5830
rect -190 -6070 50 -5830
rect 14730 -5080 14970 -4840
rect 15060 -5080 15300 -4840
rect 15390 -5080 15630 -4840
rect 15720 -5080 15960 -4840
rect 14730 -5410 14970 -5170
rect 15060 -5410 15300 -5170
rect 15390 -5410 15630 -5170
rect 15720 -5410 15960 -5170
rect 14730 -5740 14970 -5500
rect 15060 -5740 15300 -5500
rect 15390 -5740 15630 -5500
rect 15720 -5740 15960 -5500
rect 14730 -6070 14970 -5830
rect 15060 -6070 15300 -5830
rect 15390 -6070 15630 -5830
rect 15720 -6070 15960 -5830
rect 31180 -4960 31420 -4720
rect 31510 -4960 31750 -4720
rect 31840 -4960 32080 -4720
rect 32170 -4960 32410 -4720
rect 32500 -4960 32740 -4720
rect 32830 -4960 33070 -4720
rect 33160 -4960 33400 -4720
rect 33490 -4960 33730 -4720
rect 33820 -4960 34060 -4720
rect 34150 -4960 34390 -4720
rect 34480 -4960 34720 -4720
rect 34810 -4960 35050 -4720
rect 35140 -4960 35380 -4720
rect 35470 -4960 35710 -4720
rect 35800 -4960 36040 -4720
rect 36130 -4960 36370 -4720
rect 36460 -4960 36700 -4720
rect 36790 -4960 37030 -4720
rect 37120 -4960 37360 -4720
rect 37450 -4960 37690 -4720
rect 31180 -5290 31420 -5050
rect 31510 -5290 31750 -5050
rect 31840 -5290 32080 -5050
rect 32170 -5290 32410 -5050
rect 32500 -5290 32740 -5050
rect 32830 -5290 33070 -5050
rect 33160 -5290 33400 -5050
rect 33490 -5290 33730 -5050
rect 33820 -5290 34060 -5050
rect 34150 -5290 34390 -5050
rect 34480 -5290 34720 -5050
rect 34810 -5290 35050 -5050
rect 35140 -5290 35380 -5050
rect 35470 -5290 35710 -5050
rect 35800 -5290 36040 -5050
rect 36130 -5290 36370 -5050
rect 36460 -5290 36700 -5050
rect 36790 -5290 37030 -5050
rect 37120 -5290 37360 -5050
rect 37450 -5290 37690 -5050
rect 31180 -5620 31420 -5380
rect 31510 -5620 31750 -5380
rect 31840 -5620 32080 -5380
rect 32170 -5620 32410 -5380
rect 32500 -5620 32740 -5380
rect 32830 -5620 33070 -5380
rect 33160 -5620 33400 -5380
rect 33490 -5620 33730 -5380
rect 33820 -5620 34060 -5380
rect 34150 -5620 34390 -5380
rect 34480 -5620 34720 -5380
rect 34810 -5620 35050 -5380
rect 35140 -5620 35380 -5380
rect 35470 -5620 35710 -5380
rect 35800 -5620 36040 -5380
rect 36130 -5620 36370 -5380
rect 36460 -5620 36700 -5380
rect 36790 -5620 37030 -5380
rect 37120 -5620 37360 -5380
rect 37450 -5620 37690 -5380
rect 31180 -5950 31420 -5710
rect 31510 -5950 31750 -5710
rect 31840 -5950 32080 -5710
rect 32170 -5950 32410 -5710
rect 32500 -5950 32740 -5710
rect 32830 -5950 33070 -5710
rect 33160 -5950 33400 -5710
rect 33490 -5950 33730 -5710
rect 33820 -5950 34060 -5710
rect 34150 -5950 34390 -5710
rect 34480 -5950 34720 -5710
rect 34810 -5950 35050 -5710
rect 35140 -5950 35380 -5710
rect 35470 -5950 35710 -5710
rect 35800 -5950 36040 -5710
rect 36130 -5950 36370 -5710
rect 36460 -5950 36700 -5710
rect 36790 -5950 37030 -5710
rect 37120 -5950 37360 -5710
rect 37450 -5950 37690 -5710
rect 31180 -6280 31420 -6040
rect 31510 -6280 31750 -6040
rect 31840 -6280 32080 -6040
rect 32170 -6280 32410 -6040
rect 32500 -6280 32740 -6040
rect 32830 -6280 33070 -6040
rect 33160 -6280 33400 -6040
rect 33490 -6280 33730 -6040
rect 33820 -6280 34060 -6040
rect 34150 -6280 34390 -6040
rect 34480 -6280 34720 -6040
rect 34810 -6280 35050 -6040
rect 35140 -6280 35380 -6040
rect 35470 -6280 35710 -6040
rect 35800 -6280 36040 -6040
rect 36130 -6280 36370 -6040
rect 36460 -6280 36700 -6040
rect 36790 -6280 37030 -6040
rect 37120 -6280 37360 -6040
rect 37450 -6280 37690 -6040
<< metal4 >>
rect -5020 21610 7290 21640
rect -5020 21580 -4650 21610
rect -4410 21580 -4320 21610
rect -4080 21580 -3990 21610
rect -3750 21580 -3660 21610
rect -3420 21580 -3330 21610
rect -3090 21580 -3000 21610
rect -2760 21580 -2670 21610
rect -2430 21580 -2340 21610
rect -2100 21580 -2010 21610
rect -1770 21580 -1640 21610
rect -1400 21580 -1310 21610
rect -1070 21580 -980 21610
rect -740 21580 -650 21610
rect -410 21580 -320 21610
rect -80 21580 10 21610
rect 250 21580 340 21610
rect 580 21580 670 21610
rect 910 21580 1000 21610
rect 1240 21580 1370 21610
rect 1610 21580 1700 21610
rect 1940 21580 2030 21610
rect 2270 21580 2360 21610
rect 2600 21580 2690 21610
rect 2930 21580 3020 21610
rect 3260 21580 3350 21610
rect 3590 21580 3680 21610
rect 3920 21580 4010 21610
rect 4250 21580 4380 21610
rect 4620 21580 4710 21610
rect 4950 21580 5040 21610
rect 5280 21580 5370 21610
rect 5610 21580 5700 21610
rect 5940 21580 6030 21610
rect 6270 21580 6360 21610
rect 6600 21580 6690 21610
rect 6930 21580 7020 21610
rect -5020 21510 -4730 21580
rect -4660 21510 -4650 21580
rect -4390 21510 -4370 21580
rect -4030 21510 -4010 21580
rect -3750 21510 -3740 21580
rect -3670 21510 -3660 21580
rect -3400 21510 -3380 21580
rect -3040 21510 -3020 21580
rect -2760 21510 -2750 21580
rect -2680 21510 -2670 21580
rect -2410 21510 -2390 21580
rect -2050 21510 -2030 21580
rect -1770 21510 -1720 21580
rect -1650 21510 -1640 21580
rect -1380 21510 -1360 21580
rect -1020 21510 -1000 21580
rect -740 21510 -730 21580
rect -660 21510 -650 21580
rect -390 21510 -370 21580
rect -30 21510 -10 21580
rect 250 21510 260 21580
rect 330 21510 340 21580
rect 600 21510 620 21580
rect 960 21510 980 21580
rect 1240 21510 1290 21580
rect 1360 21510 1370 21580
rect 1630 21510 1650 21580
rect 1990 21510 2010 21580
rect 2270 21510 2280 21580
rect 2350 21510 2360 21580
rect 2620 21510 2640 21580
rect 2980 21510 3000 21580
rect 3260 21510 3270 21580
rect 3340 21510 3350 21580
rect 3610 21510 3630 21580
rect 3970 21510 3990 21580
rect 4250 21510 4300 21580
rect 4370 21510 4380 21580
rect 4640 21510 4660 21580
rect 5000 21510 5020 21580
rect 5280 21510 5290 21580
rect 5360 21510 5370 21580
rect 5630 21510 5650 21580
rect 5990 21510 6010 21580
rect 6270 21510 6280 21580
rect 6350 21510 6360 21580
rect 6620 21510 6640 21580
rect 6980 21510 7000 21580
rect -5020 21490 -4650 21510
rect -4410 21490 -4320 21510
rect -4080 21490 -3990 21510
rect -3750 21490 -3660 21510
rect -3420 21490 -3330 21510
rect -3090 21490 -3000 21510
rect -2760 21490 -2670 21510
rect -2430 21490 -2340 21510
rect -2100 21490 -2010 21510
rect -1770 21490 -1640 21510
rect -1400 21490 -1310 21510
rect -1070 21490 -980 21510
rect -740 21490 -650 21510
rect -410 21490 -320 21510
rect -80 21490 10 21510
rect 250 21490 340 21510
rect 580 21490 670 21510
rect 910 21490 1000 21510
rect 1240 21490 1370 21510
rect 1610 21490 1700 21510
rect 1940 21490 2030 21510
rect 2270 21490 2360 21510
rect 2600 21490 2690 21510
rect 2930 21490 3020 21510
rect 3260 21490 3350 21510
rect 3590 21490 3680 21510
rect 3920 21490 4010 21510
rect 4250 21490 4380 21510
rect 4620 21490 4710 21510
rect 4950 21490 5040 21510
rect 5280 21490 5370 21510
rect 5610 21490 5700 21510
rect 5940 21490 6030 21510
rect 6270 21490 6360 21510
rect 6600 21490 6690 21510
rect 6930 21490 7020 21510
rect -5020 21420 -4730 21490
rect -4660 21420 -4650 21490
rect -4390 21420 -4370 21490
rect -4030 21420 -4010 21490
rect -3750 21420 -3740 21490
rect -3670 21420 -3660 21490
rect -3400 21420 -3380 21490
rect -3040 21420 -3020 21490
rect -2760 21420 -2750 21490
rect -2680 21420 -2670 21490
rect -2410 21420 -2390 21490
rect -2050 21420 -2030 21490
rect -1770 21420 -1720 21490
rect -1650 21420 -1640 21490
rect -1380 21420 -1360 21490
rect -1020 21420 -1000 21490
rect -740 21420 -730 21490
rect -660 21420 -650 21490
rect -390 21420 -370 21490
rect -30 21420 -10 21490
rect 250 21420 260 21490
rect 330 21420 340 21490
rect 600 21420 620 21490
rect 960 21420 980 21490
rect 1240 21420 1290 21490
rect 1360 21420 1370 21490
rect 1630 21420 1650 21490
rect 1990 21420 2010 21490
rect 2270 21420 2280 21490
rect 2350 21420 2360 21490
rect 2620 21420 2640 21490
rect 2980 21420 3000 21490
rect 3260 21420 3270 21490
rect 3340 21420 3350 21490
rect 3610 21420 3630 21490
rect 3970 21420 3990 21490
rect 4250 21420 4300 21490
rect 4370 21420 4380 21490
rect 4640 21420 4660 21490
rect 5000 21420 5020 21490
rect 5280 21420 5290 21490
rect 5360 21420 5370 21490
rect 5630 21420 5650 21490
rect 5990 21420 6010 21490
rect 6270 21420 6280 21490
rect 6350 21420 6360 21490
rect 6620 21420 6640 21490
rect 6980 21420 7000 21490
rect -5020 21400 -4650 21420
rect -4410 21400 -4320 21420
rect -4080 21400 -3990 21420
rect -3750 21400 -3660 21420
rect -3420 21400 -3330 21420
rect -3090 21400 -3000 21420
rect -2760 21400 -2670 21420
rect -2430 21400 -2340 21420
rect -2100 21400 -2010 21420
rect -1770 21400 -1640 21420
rect -1400 21400 -1310 21420
rect -1070 21400 -980 21420
rect -740 21400 -650 21420
rect -410 21400 -320 21420
rect -80 21400 10 21420
rect 250 21400 340 21420
rect 580 21400 670 21420
rect 910 21400 1000 21420
rect 1240 21400 1370 21420
rect 1610 21400 1700 21420
rect 1940 21400 2030 21420
rect 2270 21400 2360 21420
rect 2600 21400 2690 21420
rect 2930 21400 3020 21420
rect 3260 21400 3350 21420
rect 3590 21400 3680 21420
rect 3920 21400 4010 21420
rect 4250 21400 4380 21420
rect 4620 21400 4710 21420
rect 4950 21400 5040 21420
rect 5280 21400 5370 21420
rect 5610 21400 5700 21420
rect 5940 21400 6030 21420
rect 6270 21400 6360 21420
rect 6600 21400 6690 21420
rect 6930 21400 7020 21420
rect -5020 21330 -4730 21400
rect -4660 21370 -4650 21400
rect -4660 21330 -4640 21370
rect -4570 21330 -4550 21370
rect -4480 21330 -4460 21370
rect -4390 21330 -4370 21400
rect -4300 21330 -4280 21370
rect -4210 21330 -4190 21370
rect -4120 21330 -4100 21370
rect -4030 21330 -4010 21400
rect -3750 21370 -3740 21400
rect -3940 21330 -3920 21370
rect -3850 21330 -3830 21370
rect -3760 21330 -3740 21370
rect -3670 21370 -3660 21400
rect -3670 21330 -3650 21370
rect -3580 21330 -3560 21370
rect -3490 21330 -3470 21370
rect -3400 21330 -3380 21400
rect -3310 21330 -3290 21370
rect -3220 21330 -3200 21370
rect -3130 21330 -3110 21370
rect -3040 21330 -3020 21400
rect -2760 21370 -2750 21400
rect -2950 21330 -2930 21370
rect -2860 21330 -2840 21370
rect -2770 21330 -2750 21370
rect -2680 21370 -2670 21400
rect -2680 21330 -2660 21370
rect -2590 21330 -2570 21370
rect -2500 21330 -2480 21370
rect -2410 21330 -2390 21400
rect -2320 21330 -2300 21370
rect -2230 21330 -2210 21370
rect -2140 21330 -2120 21370
rect -2050 21330 -2030 21400
rect -1770 21370 -1720 21400
rect -1960 21330 -1940 21370
rect -1870 21330 -1850 21370
rect -1780 21330 -1720 21370
rect -1650 21370 -1640 21400
rect -1650 21330 -1630 21370
rect -1560 21330 -1540 21370
rect -1470 21330 -1450 21370
rect -1380 21330 -1360 21400
rect -1290 21330 -1270 21370
rect -1200 21330 -1180 21370
rect -1110 21330 -1090 21370
rect -1020 21330 -1000 21400
rect -740 21370 -730 21400
rect -930 21330 -910 21370
rect -840 21330 -820 21370
rect -750 21330 -730 21370
rect -660 21370 -650 21400
rect -660 21330 -640 21370
rect -570 21330 -550 21370
rect -480 21330 -460 21370
rect -390 21330 -370 21400
rect -300 21330 -280 21370
rect -210 21330 -190 21370
rect -120 21330 -100 21370
rect -30 21330 -10 21400
rect 250 21370 260 21400
rect 60 21330 80 21370
rect 150 21330 170 21370
rect 240 21330 260 21370
rect 330 21370 340 21400
rect 330 21330 350 21370
rect 420 21330 440 21370
rect 510 21330 530 21370
rect 600 21330 620 21400
rect 690 21330 710 21370
rect 780 21330 800 21370
rect 870 21330 890 21370
rect 960 21330 980 21400
rect 1240 21370 1290 21400
rect 1050 21330 1070 21370
rect 1140 21330 1160 21370
rect 1230 21330 1290 21370
rect 1360 21370 1370 21400
rect 1360 21330 1380 21370
rect 1450 21330 1470 21370
rect 1540 21330 1560 21370
rect 1630 21330 1650 21400
rect 1720 21330 1740 21370
rect 1810 21330 1830 21370
rect 1900 21330 1920 21370
rect 1990 21330 2010 21400
rect 2270 21370 2280 21400
rect 2080 21330 2100 21370
rect 2170 21330 2190 21370
rect 2260 21330 2280 21370
rect 2350 21370 2360 21400
rect 2350 21330 2370 21370
rect 2440 21330 2460 21370
rect 2530 21330 2550 21370
rect 2620 21330 2640 21400
rect 2710 21330 2730 21370
rect 2800 21330 2820 21370
rect 2890 21330 2910 21370
rect 2980 21330 3000 21400
rect 3260 21370 3270 21400
rect 3070 21330 3090 21370
rect 3160 21330 3180 21370
rect 3250 21330 3270 21370
rect 3340 21370 3350 21400
rect 3340 21330 3360 21370
rect 3430 21330 3450 21370
rect 3520 21330 3540 21370
rect 3610 21330 3630 21400
rect 3700 21330 3720 21370
rect 3790 21330 3810 21370
rect 3880 21330 3900 21370
rect 3970 21330 3990 21400
rect 4250 21370 4300 21400
rect 4060 21330 4080 21370
rect 4150 21330 4170 21370
rect 4240 21330 4300 21370
rect 4370 21370 4380 21400
rect 4370 21330 4390 21370
rect 4460 21330 4480 21370
rect 4550 21330 4570 21370
rect 4640 21330 4660 21400
rect 4730 21330 4750 21370
rect 4820 21330 4840 21370
rect 4910 21330 4930 21370
rect 5000 21330 5020 21400
rect 5280 21370 5290 21400
rect 5090 21330 5110 21370
rect 5180 21330 5200 21370
rect 5270 21330 5290 21370
rect 5360 21370 5370 21400
rect 5360 21330 5380 21370
rect 5450 21330 5470 21370
rect 5540 21330 5560 21370
rect 5630 21330 5650 21400
rect 5720 21330 5740 21370
rect 5810 21330 5830 21370
rect 5900 21330 5920 21370
rect 5990 21330 6010 21400
rect 6270 21370 6280 21400
rect 6080 21330 6100 21370
rect 6170 21330 6190 21370
rect 6260 21330 6280 21370
rect 6350 21370 6360 21400
rect 6350 21330 6370 21370
rect 6440 21330 6460 21370
rect 6530 21330 6550 21370
rect 6620 21330 6640 21400
rect 6710 21330 6730 21370
rect 6800 21330 6820 21370
rect 6890 21330 6910 21370
rect 6980 21330 7000 21400
rect 7260 21370 7290 21610
rect 7070 21330 7090 21370
rect 7160 21330 7180 21370
rect 7250 21330 7290 21370
rect -5020 21320 7290 21330
rect 7610 21610 19920 21640
rect 7610 21370 7640 21610
rect 7880 21580 7970 21610
rect 8210 21580 8300 21610
rect 8540 21580 8630 21610
rect 8870 21580 8960 21610
rect 9200 21580 9290 21610
rect 9530 21580 9620 21610
rect 9860 21580 9950 21610
rect 10190 21580 10280 21610
rect 10520 21580 10650 21610
rect 10890 21580 10980 21610
rect 11220 21580 11310 21610
rect 11550 21580 11640 21610
rect 11880 21580 11970 21610
rect 12210 21580 12300 21610
rect 12540 21580 12630 21610
rect 12870 21580 12960 21610
rect 13200 21580 13290 21610
rect 13530 21580 13660 21610
rect 13900 21580 13990 21610
rect 14230 21580 14320 21610
rect 14560 21580 14650 21610
rect 14890 21580 14980 21610
rect 15220 21580 15310 21610
rect 15550 21580 15640 21610
rect 15880 21580 15970 21610
rect 16210 21580 16300 21610
rect 16540 21580 16670 21610
rect 16910 21580 17000 21610
rect 17240 21580 17330 21610
rect 17570 21580 17660 21610
rect 17900 21580 17990 21610
rect 18230 21580 18320 21610
rect 18560 21580 18650 21610
rect 18890 21580 18980 21610
rect 19220 21580 19310 21610
rect 19550 21580 19920 21610
rect 7900 21510 7920 21580
rect 8260 21510 8280 21580
rect 8540 21510 8550 21580
rect 8620 21510 8630 21580
rect 8890 21510 8910 21580
rect 9250 21510 9270 21580
rect 9530 21510 9540 21580
rect 9610 21510 9620 21580
rect 9880 21510 9900 21580
rect 10240 21510 10260 21580
rect 10520 21510 10530 21580
rect 10600 21510 10650 21580
rect 10910 21510 10930 21580
rect 11270 21510 11290 21580
rect 11550 21510 11560 21580
rect 11630 21510 11640 21580
rect 11900 21510 11920 21580
rect 12260 21510 12280 21580
rect 12540 21510 12550 21580
rect 12620 21510 12630 21580
rect 12890 21510 12910 21580
rect 13250 21510 13270 21580
rect 13530 21510 13540 21580
rect 13610 21510 13660 21580
rect 13920 21510 13940 21580
rect 14280 21510 14300 21580
rect 14560 21510 14570 21580
rect 14640 21510 14650 21580
rect 14910 21510 14930 21580
rect 15270 21510 15290 21580
rect 15550 21510 15560 21580
rect 15630 21510 15640 21580
rect 15900 21510 15920 21580
rect 16260 21510 16280 21580
rect 16540 21510 16550 21580
rect 16620 21510 16670 21580
rect 16930 21510 16950 21580
rect 17290 21510 17310 21580
rect 17570 21510 17580 21580
rect 17650 21510 17660 21580
rect 17920 21510 17940 21580
rect 18280 21510 18300 21580
rect 18560 21510 18570 21580
rect 18640 21510 18650 21580
rect 18910 21510 18930 21580
rect 19270 21510 19290 21580
rect 19550 21510 19560 21580
rect 19630 21510 19920 21580
rect 7880 21490 7970 21510
rect 8210 21490 8300 21510
rect 8540 21490 8630 21510
rect 8870 21490 8960 21510
rect 9200 21490 9290 21510
rect 9530 21490 9620 21510
rect 9860 21490 9950 21510
rect 10190 21490 10280 21510
rect 10520 21490 10650 21510
rect 10890 21490 10980 21510
rect 11220 21490 11310 21510
rect 11550 21490 11640 21510
rect 11880 21490 11970 21510
rect 12210 21490 12300 21510
rect 12540 21490 12630 21510
rect 12870 21490 12960 21510
rect 13200 21490 13290 21510
rect 13530 21490 13660 21510
rect 13900 21490 13990 21510
rect 14230 21490 14320 21510
rect 14560 21490 14650 21510
rect 14890 21490 14980 21510
rect 15220 21490 15310 21510
rect 15550 21490 15640 21510
rect 15880 21490 15970 21510
rect 16210 21490 16300 21510
rect 16540 21490 16670 21510
rect 16910 21490 17000 21510
rect 17240 21490 17330 21510
rect 17570 21490 17660 21510
rect 17900 21490 17990 21510
rect 18230 21490 18320 21510
rect 18560 21490 18650 21510
rect 18890 21490 18980 21510
rect 19220 21490 19310 21510
rect 19550 21490 19920 21510
rect 7900 21420 7920 21490
rect 8260 21420 8280 21490
rect 8540 21420 8550 21490
rect 8620 21420 8630 21490
rect 8890 21420 8910 21490
rect 9250 21420 9270 21490
rect 9530 21420 9540 21490
rect 9610 21420 9620 21490
rect 9880 21420 9900 21490
rect 10240 21420 10260 21490
rect 10520 21420 10530 21490
rect 10600 21420 10650 21490
rect 10910 21420 10930 21490
rect 11270 21420 11290 21490
rect 11550 21420 11560 21490
rect 11630 21420 11640 21490
rect 11900 21420 11920 21490
rect 12260 21420 12280 21490
rect 12540 21420 12550 21490
rect 12620 21420 12630 21490
rect 12890 21420 12910 21490
rect 13250 21420 13270 21490
rect 13530 21420 13540 21490
rect 13610 21420 13660 21490
rect 13920 21420 13940 21490
rect 14280 21420 14300 21490
rect 14560 21420 14570 21490
rect 14640 21420 14650 21490
rect 14910 21420 14930 21490
rect 15270 21420 15290 21490
rect 15550 21420 15560 21490
rect 15630 21420 15640 21490
rect 15900 21420 15920 21490
rect 16260 21420 16280 21490
rect 16540 21420 16550 21490
rect 16620 21420 16670 21490
rect 16930 21420 16950 21490
rect 17290 21420 17310 21490
rect 17570 21420 17580 21490
rect 17650 21420 17660 21490
rect 17920 21420 17940 21490
rect 18280 21420 18300 21490
rect 18560 21420 18570 21490
rect 18640 21420 18650 21490
rect 18910 21420 18930 21490
rect 19270 21420 19290 21490
rect 19550 21420 19560 21490
rect 19630 21420 19920 21490
rect 7880 21400 7970 21420
rect 8210 21400 8300 21420
rect 8540 21400 8630 21420
rect 8870 21400 8960 21420
rect 9200 21400 9290 21420
rect 9530 21400 9620 21420
rect 9860 21400 9950 21420
rect 10190 21400 10280 21420
rect 10520 21400 10650 21420
rect 10890 21400 10980 21420
rect 11220 21400 11310 21420
rect 11550 21400 11640 21420
rect 11880 21400 11970 21420
rect 12210 21400 12300 21420
rect 12540 21400 12630 21420
rect 12870 21400 12960 21420
rect 13200 21400 13290 21420
rect 13530 21400 13660 21420
rect 13900 21400 13990 21420
rect 14230 21400 14320 21420
rect 14560 21400 14650 21420
rect 14890 21400 14980 21420
rect 15220 21400 15310 21420
rect 15550 21400 15640 21420
rect 15880 21400 15970 21420
rect 16210 21400 16300 21420
rect 16540 21400 16670 21420
rect 16910 21400 17000 21420
rect 17240 21400 17330 21420
rect 17570 21400 17660 21420
rect 17900 21400 17990 21420
rect 18230 21400 18320 21420
rect 18560 21400 18650 21420
rect 18890 21400 18980 21420
rect 19220 21400 19310 21420
rect 19550 21400 19920 21420
rect 7610 21330 7650 21370
rect 7720 21330 7740 21370
rect 7810 21330 7830 21370
rect 7900 21330 7920 21400
rect 7990 21330 8010 21370
rect 8080 21330 8100 21370
rect 8170 21330 8190 21370
rect 8260 21330 8280 21400
rect 8540 21370 8550 21400
rect 8350 21330 8370 21370
rect 8440 21330 8460 21370
rect 8530 21330 8550 21370
rect 8620 21370 8630 21400
rect 8620 21330 8640 21370
rect 8710 21330 8730 21370
rect 8800 21330 8820 21370
rect 8890 21330 8910 21400
rect 8980 21330 9000 21370
rect 9070 21330 9090 21370
rect 9160 21330 9180 21370
rect 9250 21330 9270 21400
rect 9530 21370 9540 21400
rect 9340 21330 9360 21370
rect 9430 21330 9450 21370
rect 9520 21330 9540 21370
rect 9610 21370 9620 21400
rect 9610 21330 9630 21370
rect 9700 21330 9720 21370
rect 9790 21330 9810 21370
rect 9880 21330 9900 21400
rect 9970 21330 9990 21370
rect 10060 21330 10080 21370
rect 10150 21330 10170 21370
rect 10240 21330 10260 21400
rect 10520 21370 10530 21400
rect 10330 21330 10350 21370
rect 10420 21330 10440 21370
rect 10510 21330 10530 21370
rect 10600 21370 10650 21400
rect 10600 21330 10660 21370
rect 10730 21330 10750 21370
rect 10820 21330 10840 21370
rect 10910 21330 10930 21400
rect 11000 21330 11020 21370
rect 11090 21330 11110 21370
rect 11180 21330 11200 21370
rect 11270 21330 11290 21400
rect 11550 21370 11560 21400
rect 11360 21330 11380 21370
rect 11450 21330 11470 21370
rect 11540 21330 11560 21370
rect 11630 21370 11640 21400
rect 11630 21330 11650 21370
rect 11720 21330 11740 21370
rect 11810 21330 11830 21370
rect 11900 21330 11920 21400
rect 11990 21330 12010 21370
rect 12080 21330 12100 21370
rect 12170 21330 12190 21370
rect 12260 21330 12280 21400
rect 12540 21370 12550 21400
rect 12350 21330 12370 21370
rect 12440 21330 12460 21370
rect 12530 21330 12550 21370
rect 12620 21370 12630 21400
rect 12620 21330 12640 21370
rect 12710 21330 12730 21370
rect 12800 21330 12820 21370
rect 12890 21330 12910 21400
rect 12980 21330 13000 21370
rect 13070 21330 13090 21370
rect 13160 21330 13180 21370
rect 13250 21330 13270 21400
rect 13530 21370 13540 21400
rect 13340 21330 13360 21370
rect 13430 21330 13450 21370
rect 13520 21330 13540 21370
rect 13610 21370 13660 21400
rect 13610 21330 13670 21370
rect 13740 21330 13760 21370
rect 13830 21330 13850 21370
rect 13920 21330 13940 21400
rect 14010 21330 14030 21370
rect 14100 21330 14120 21370
rect 14190 21330 14210 21370
rect 14280 21330 14300 21400
rect 14560 21370 14570 21400
rect 14370 21330 14390 21370
rect 14460 21330 14480 21370
rect 14550 21330 14570 21370
rect 14640 21370 14650 21400
rect 14640 21330 14660 21370
rect 14730 21330 14750 21370
rect 14820 21330 14840 21370
rect 14910 21330 14930 21400
rect 15000 21330 15020 21370
rect 15090 21330 15110 21370
rect 15180 21330 15200 21370
rect 15270 21330 15290 21400
rect 15550 21370 15560 21400
rect 15360 21330 15380 21370
rect 15450 21330 15470 21370
rect 15540 21330 15560 21370
rect 15630 21370 15640 21400
rect 15630 21330 15650 21370
rect 15720 21330 15740 21370
rect 15810 21330 15830 21370
rect 15900 21330 15920 21400
rect 15990 21330 16010 21370
rect 16080 21330 16100 21370
rect 16170 21330 16190 21370
rect 16260 21330 16280 21400
rect 16540 21370 16550 21400
rect 16350 21330 16370 21370
rect 16440 21330 16460 21370
rect 16530 21330 16550 21370
rect 16620 21370 16670 21400
rect 16620 21330 16680 21370
rect 16750 21330 16770 21370
rect 16840 21330 16860 21370
rect 16930 21330 16950 21400
rect 17020 21330 17040 21370
rect 17110 21330 17130 21370
rect 17200 21330 17220 21370
rect 17290 21330 17310 21400
rect 17570 21370 17580 21400
rect 17380 21330 17400 21370
rect 17470 21330 17490 21370
rect 17560 21330 17580 21370
rect 17650 21370 17660 21400
rect 17650 21330 17670 21370
rect 17740 21330 17760 21370
rect 17830 21330 17850 21370
rect 17920 21330 17940 21400
rect 18010 21330 18030 21370
rect 18100 21330 18120 21370
rect 18190 21330 18210 21370
rect 18280 21330 18300 21400
rect 18560 21370 18570 21400
rect 18370 21330 18390 21370
rect 18460 21330 18480 21370
rect 18550 21330 18570 21370
rect 18640 21370 18650 21400
rect 18640 21330 18660 21370
rect 18730 21330 18750 21370
rect 18820 21330 18840 21370
rect 18910 21330 18930 21400
rect 19000 21330 19020 21370
rect 19090 21330 19110 21370
rect 19180 21330 19200 21370
rect 19270 21330 19290 21400
rect 19550 21370 19560 21400
rect 19360 21330 19380 21370
rect 19450 21330 19470 21370
rect 19540 21330 19560 21370
rect 19630 21330 19920 21400
rect 7610 21320 19920 21330
rect -5020 20830 7290 21000
rect -5020 20590 -4670 20830
rect -4430 20590 -4340 20830
rect -4100 20590 -4010 20830
rect -3770 20590 -3680 20830
rect -3440 20590 -3350 20830
rect -3110 20590 -3020 20830
rect -2780 20590 -2690 20830
rect -2450 20590 -2360 20830
rect -2120 20590 -2030 20830
rect -1790 20590 -1700 20830
rect -1460 20590 -1370 20830
rect -1130 20590 -1040 20830
rect -800 20590 -710 20830
rect -470 20590 -380 20830
rect -140 20590 -50 20830
rect 190 20590 280 20830
rect 520 20590 610 20830
rect 850 20590 940 20830
rect 1180 20590 1270 20830
rect 1510 20590 1600 20830
rect 1840 20590 1930 20830
rect 2170 20590 2260 20830
rect 2500 20590 2590 20830
rect 2830 20590 2920 20830
rect 3160 20590 3250 20830
rect 3490 20590 3580 20830
rect 3820 20590 3910 20830
rect 4150 20590 4240 20830
rect 4480 20590 4570 20830
rect 4810 20590 4900 20830
rect 5140 20590 5230 20830
rect 5470 20590 5560 20830
rect 5800 20590 5890 20830
rect 6130 20590 6220 20830
rect 6460 20590 6550 20830
rect 6790 20590 6880 20830
rect 7120 20590 7290 20830
rect -5020 20500 7290 20590
rect -5020 20260 -4670 20500
rect -4430 20260 -4340 20500
rect -4100 20260 -4010 20500
rect -3770 20260 -3680 20500
rect -3440 20260 -3350 20500
rect -3110 20260 -3020 20500
rect -2780 20260 -2690 20500
rect -2450 20260 -2360 20500
rect -2120 20260 -2030 20500
rect -1790 20260 -1700 20500
rect -1460 20260 -1370 20500
rect -1130 20260 -1040 20500
rect -800 20260 -710 20500
rect -470 20260 -380 20500
rect -140 20260 -50 20500
rect 190 20260 280 20500
rect 520 20260 610 20500
rect 850 20260 940 20500
rect 1180 20260 1270 20500
rect 1510 20260 1600 20500
rect 1840 20260 1930 20500
rect 2170 20260 2260 20500
rect 2500 20260 2590 20500
rect 2830 20260 2920 20500
rect 3160 20260 3250 20500
rect 3490 20260 3580 20500
rect 3820 20260 3910 20500
rect 4150 20260 4240 20500
rect 4480 20260 4570 20500
rect 4810 20260 4900 20500
rect 5140 20260 5230 20500
rect 5470 20260 5560 20500
rect 5800 20260 5890 20500
rect 6130 20260 6220 20500
rect 6460 20260 6550 20500
rect 6790 20260 6880 20500
rect 7120 20260 7290 20500
rect -5020 20170 7290 20260
rect -5020 19930 -4670 20170
rect -4430 19930 -4340 20170
rect -4100 19930 -4010 20170
rect -3770 19930 -3680 20170
rect -3440 19930 -3350 20170
rect -3110 19930 -3020 20170
rect -2780 19930 -2690 20170
rect -2450 19930 -2360 20170
rect -2120 19930 -2030 20170
rect -1790 19930 -1700 20170
rect -1460 19930 -1370 20170
rect -1130 19930 -1040 20170
rect -800 19930 -710 20170
rect -470 19930 -380 20170
rect -140 19930 -50 20170
rect 190 19930 280 20170
rect 520 19930 610 20170
rect 850 19930 940 20170
rect 1180 19930 1270 20170
rect 1510 19930 1600 20170
rect 1840 19930 1930 20170
rect 2170 19930 2260 20170
rect 2500 19930 2590 20170
rect 2830 19930 2920 20170
rect 3160 19930 3250 20170
rect 3490 19930 3580 20170
rect 3820 19930 3910 20170
rect 4150 19930 4240 20170
rect 4480 19930 4570 20170
rect 4810 19930 4900 20170
rect 5140 19930 5230 20170
rect 5470 19930 5560 20170
rect 5800 19930 5890 20170
rect 6130 19930 6220 20170
rect 6460 19930 6550 20170
rect 6790 19930 6880 20170
rect 7120 19930 7290 20170
rect -5020 19840 7290 19930
rect -5020 19600 -4670 19840
rect -4430 19600 -4340 19840
rect -4100 19600 -4010 19840
rect -3770 19600 -3680 19840
rect -3440 19600 -3350 19840
rect -3110 19600 -3020 19840
rect -2780 19600 -2690 19840
rect -2450 19600 -2360 19840
rect -2120 19600 -2030 19840
rect -1790 19600 -1700 19840
rect -1460 19600 -1370 19840
rect -1130 19600 -1040 19840
rect -800 19600 -710 19840
rect -470 19600 -380 19840
rect -140 19600 -50 19840
rect 190 19600 280 19840
rect 520 19600 610 19840
rect 850 19600 940 19840
rect 1180 19600 1270 19840
rect 1510 19600 1600 19840
rect 1840 19600 1930 19840
rect 2170 19600 2260 19840
rect 2500 19600 2590 19840
rect 2830 19600 2920 19840
rect 3160 19600 3250 19840
rect 3490 19600 3580 19840
rect 3820 19600 3910 19840
rect 4150 19600 4240 19840
rect 4480 19600 4570 19840
rect 4810 19600 4900 19840
rect 5140 19600 5230 19840
rect 5470 19600 5560 19840
rect 5800 19600 5890 19840
rect 6130 19600 6220 19840
rect 6460 19600 6550 19840
rect 6790 19600 6880 19840
rect 7120 19600 7290 19840
rect -5020 19510 7290 19600
rect -5020 19270 -4670 19510
rect -4430 19270 -4340 19510
rect -4100 19270 -4010 19510
rect -3770 19270 -3680 19510
rect -3440 19270 -3350 19510
rect -3110 19270 -3020 19510
rect -2780 19270 -2690 19510
rect -2450 19270 -2360 19510
rect -2120 19270 -2030 19510
rect -1790 19270 -1700 19510
rect -1460 19270 -1370 19510
rect -1130 19270 -1040 19510
rect -800 19270 -710 19510
rect -470 19270 -380 19510
rect -140 19270 -50 19510
rect 190 19270 280 19510
rect 520 19270 610 19510
rect 850 19270 940 19510
rect 1180 19270 1270 19510
rect 1510 19270 1600 19510
rect 1840 19270 1930 19510
rect 2170 19270 2260 19510
rect 2500 19270 2590 19510
rect 2830 19270 2920 19510
rect 3160 19270 3250 19510
rect 3490 19270 3580 19510
rect 3820 19270 3910 19510
rect 4150 19270 4240 19510
rect 4480 19270 4570 19510
rect 4810 19270 4900 19510
rect 5140 19270 5230 19510
rect 5470 19270 5560 19510
rect 5800 19270 5890 19510
rect 6130 19270 6220 19510
rect 6460 19270 6550 19510
rect 6790 19270 6880 19510
rect 7120 19270 7290 19510
rect -5020 19180 7290 19270
rect -5020 18940 -4670 19180
rect -4430 18940 -4340 19180
rect -4100 18940 -4010 19180
rect -3770 18940 -3680 19180
rect -3440 18940 -3350 19180
rect -3110 18940 -3020 19180
rect -2780 18940 -2690 19180
rect -2450 18940 -2360 19180
rect -2120 18940 -2030 19180
rect -1790 18940 -1700 19180
rect -1460 18940 -1370 19180
rect -1130 18940 -1040 19180
rect -800 18940 -710 19180
rect -470 18940 -380 19180
rect -140 18940 -50 19180
rect 190 18940 280 19180
rect 520 18940 610 19180
rect 850 18940 940 19180
rect 1180 18940 1270 19180
rect 1510 18940 1600 19180
rect 1840 18940 1930 19180
rect 2170 18940 2260 19180
rect 2500 18940 2590 19180
rect 2830 18940 2920 19180
rect 3160 18940 3250 19180
rect 3490 18940 3580 19180
rect 3820 18940 3910 19180
rect 4150 18940 4240 19180
rect 4480 18940 4570 19180
rect 4810 18940 4900 19180
rect 5140 18940 5230 19180
rect 5470 18940 5560 19180
rect 5800 18940 5890 19180
rect 6130 18940 6220 19180
rect 6460 18940 6550 19180
rect 6790 18940 6880 19180
rect 7120 18940 7290 19180
rect -5020 18850 7290 18940
rect -5020 18610 -4670 18850
rect -4430 18610 -4340 18850
rect -4100 18610 -4010 18850
rect -3770 18610 -3680 18850
rect -3440 18610 -3350 18850
rect -3110 18610 -3020 18850
rect -2780 18610 -2690 18850
rect -2450 18610 -2360 18850
rect -2120 18610 -2030 18850
rect -1790 18610 -1700 18850
rect -1460 18610 -1370 18850
rect -1130 18610 -1040 18850
rect -800 18610 -710 18850
rect -470 18610 -380 18850
rect -140 18610 -50 18850
rect 190 18610 280 18850
rect 520 18610 610 18850
rect 850 18610 940 18850
rect 1180 18610 1270 18850
rect 1510 18610 1600 18850
rect 1840 18610 1930 18850
rect 2170 18610 2260 18850
rect 2500 18610 2590 18850
rect 2830 18610 2920 18850
rect 3160 18610 3250 18850
rect 3490 18610 3580 18850
rect 3820 18610 3910 18850
rect 4150 18610 4240 18850
rect 4480 18610 4570 18850
rect 4810 18610 4900 18850
rect 5140 18610 5230 18850
rect 5470 18610 5560 18850
rect 5800 18610 5890 18850
rect 6130 18610 6220 18850
rect 6460 18610 6550 18850
rect 6790 18610 6880 18850
rect 7120 18610 7290 18850
rect -5020 18520 7290 18610
rect -5020 18280 -4670 18520
rect -4430 18280 -4340 18520
rect -4100 18280 -4010 18520
rect -3770 18280 -3680 18520
rect -3440 18280 -3350 18520
rect -3110 18280 -3020 18520
rect -2780 18280 -2690 18520
rect -2450 18280 -2360 18520
rect -2120 18280 -2030 18520
rect -1790 18280 -1700 18520
rect -1460 18280 -1370 18520
rect -1130 18280 -1040 18520
rect -800 18280 -710 18520
rect -470 18280 -380 18520
rect -140 18280 -50 18520
rect 190 18280 280 18520
rect 520 18280 610 18520
rect 850 18280 940 18520
rect 1180 18280 1270 18520
rect 1510 18280 1600 18520
rect 1840 18280 1930 18520
rect 2170 18280 2260 18520
rect 2500 18280 2590 18520
rect 2830 18280 2920 18520
rect 3160 18280 3250 18520
rect 3490 18280 3580 18520
rect 3820 18280 3910 18520
rect 4150 18280 4240 18520
rect 4480 18280 4570 18520
rect 4810 18280 4900 18520
rect 5140 18280 5230 18520
rect 5470 18280 5560 18520
rect 5800 18280 5890 18520
rect 6130 18280 6220 18520
rect 6460 18280 6550 18520
rect 6790 18280 6880 18520
rect 7120 18280 7290 18520
rect -5020 18190 7290 18280
rect -5020 17950 -4670 18190
rect -4430 17950 -4340 18190
rect -4100 17950 -4010 18190
rect -3770 17950 -3680 18190
rect -3440 17950 -3350 18190
rect -3110 17950 -3020 18190
rect -2780 17950 -2690 18190
rect -2450 17950 -2360 18190
rect -2120 17950 -2030 18190
rect -1790 17950 -1700 18190
rect -1460 17950 -1370 18190
rect -1130 17950 -1040 18190
rect -800 17950 -710 18190
rect -470 17950 -380 18190
rect -140 17950 -50 18190
rect 190 17950 280 18190
rect 520 17950 610 18190
rect 850 17950 940 18190
rect 1180 17950 1270 18190
rect 1510 17950 1600 18190
rect 1840 17950 1930 18190
rect 2170 17950 2260 18190
rect 2500 17950 2590 18190
rect 2830 17950 2920 18190
rect 3160 17950 3250 18190
rect 3490 17950 3580 18190
rect 3820 17950 3910 18190
rect 4150 17950 4240 18190
rect 4480 17950 4570 18190
rect 4810 17950 4900 18190
rect 5140 17950 5230 18190
rect 5470 17950 5560 18190
rect 5800 17950 5890 18190
rect 6130 17950 6220 18190
rect 6460 17950 6550 18190
rect 6790 17950 6880 18190
rect 7120 17950 7290 18190
rect -5020 17860 7290 17950
rect -5020 17620 -4670 17860
rect -4430 17620 -4340 17860
rect -4100 17620 -4010 17860
rect -3770 17620 -3680 17860
rect -3440 17620 -3350 17860
rect -3110 17620 -3020 17860
rect -2780 17620 -2690 17860
rect -2450 17620 -2360 17860
rect -2120 17620 -2030 17860
rect -1790 17620 -1700 17860
rect -1460 17620 -1370 17860
rect -1130 17620 -1040 17860
rect -800 17620 -710 17860
rect -470 17620 -380 17860
rect -140 17620 -50 17860
rect 190 17620 280 17860
rect 520 17620 610 17860
rect 850 17620 940 17860
rect 1180 17620 1270 17860
rect 1510 17620 1600 17860
rect 1840 17620 1930 17860
rect 2170 17620 2260 17860
rect 2500 17620 2590 17860
rect 2830 17620 2920 17860
rect 3160 17620 3250 17860
rect 3490 17620 3580 17860
rect 3820 17620 3910 17860
rect 4150 17620 4240 17860
rect 4480 17620 4570 17860
rect 4810 17620 4900 17860
rect 5140 17620 5230 17860
rect 5470 17620 5560 17860
rect 5800 17620 5890 17860
rect 6130 17620 6220 17860
rect 6460 17620 6550 17860
rect 6790 17620 6880 17860
rect 7120 17620 7290 17860
rect -5020 17530 7290 17620
rect -5020 17290 -4670 17530
rect -4430 17290 -4340 17530
rect -4100 17290 -4010 17530
rect -3770 17290 -3680 17530
rect -3440 17290 -3350 17530
rect -3110 17290 -3020 17530
rect -2780 17290 -2690 17530
rect -2450 17290 -2360 17530
rect -2120 17290 -2030 17530
rect -1790 17290 -1700 17530
rect -1460 17290 -1370 17530
rect -1130 17290 -1040 17530
rect -800 17290 -710 17530
rect -470 17290 -380 17530
rect -140 17290 -50 17530
rect 190 17290 280 17530
rect 520 17290 610 17530
rect 850 17290 940 17530
rect 1180 17290 1270 17530
rect 1510 17290 1600 17530
rect 1840 17290 1930 17530
rect 2170 17290 2260 17530
rect 2500 17290 2590 17530
rect 2830 17290 2920 17530
rect 3160 17290 3250 17530
rect 3490 17290 3580 17530
rect 3820 17290 3910 17530
rect 4150 17290 4240 17530
rect 4480 17290 4570 17530
rect 4810 17290 4900 17530
rect 5140 17290 5230 17530
rect 5470 17290 5560 17530
rect 5800 17290 5890 17530
rect 6130 17290 6220 17530
rect 6460 17290 6550 17530
rect 6790 17290 6880 17530
rect 7120 17290 7290 17530
rect -5020 17200 7290 17290
rect -5020 16960 -4670 17200
rect -4430 16960 -4340 17200
rect -4100 16960 -4010 17200
rect -3770 16960 -3680 17200
rect -3440 16960 -3350 17200
rect -3110 16960 -3020 17200
rect -2780 16960 -2690 17200
rect -2450 16960 -2360 17200
rect -2120 16960 -2030 17200
rect -1790 16960 -1700 17200
rect -1460 16960 -1370 17200
rect -1130 16960 -1040 17200
rect -800 16960 -710 17200
rect -470 16960 -380 17200
rect -140 16960 -50 17200
rect 190 16960 280 17200
rect 520 16960 610 17200
rect 850 16960 940 17200
rect 1180 16960 1270 17200
rect 1510 16960 1600 17200
rect 1840 16960 1930 17200
rect 2170 16960 2260 17200
rect 2500 16960 2590 17200
rect 2830 16960 2920 17200
rect 3160 16960 3250 17200
rect 3490 16960 3580 17200
rect 3820 16960 3910 17200
rect 4150 16960 4240 17200
rect 4480 16960 4570 17200
rect 4810 16960 4900 17200
rect 5140 16960 5230 17200
rect 5470 16960 5560 17200
rect 5800 16960 5890 17200
rect 6130 16960 6220 17200
rect 6460 16960 6550 17200
rect 6790 16960 6880 17200
rect 7120 16960 7290 17200
rect -5020 16870 7290 16960
rect -5020 16630 -4670 16870
rect -4430 16630 -4340 16870
rect -4100 16630 -4010 16870
rect -3770 16630 -3680 16870
rect -3440 16630 -3350 16870
rect -3110 16630 -3020 16870
rect -2780 16630 -2690 16870
rect -2450 16630 -2360 16870
rect -2120 16630 -2030 16870
rect -1790 16630 -1700 16870
rect -1460 16630 -1370 16870
rect -1130 16630 -1040 16870
rect -800 16630 -710 16870
rect -470 16630 -380 16870
rect -140 16630 -50 16870
rect 190 16630 280 16870
rect 520 16630 610 16870
rect 850 16630 940 16870
rect 1180 16630 1270 16870
rect 1510 16630 1600 16870
rect 1840 16630 1930 16870
rect 2170 16630 2260 16870
rect 2500 16630 2590 16870
rect 2830 16630 2920 16870
rect 3160 16630 3250 16870
rect 3490 16630 3580 16870
rect 3820 16630 3910 16870
rect 4150 16630 4240 16870
rect 4480 16630 4570 16870
rect 4810 16630 4900 16870
rect 5140 16630 5230 16870
rect 5470 16630 5560 16870
rect 5800 16630 5890 16870
rect 6130 16630 6220 16870
rect 6460 16630 6550 16870
rect 6790 16630 6880 16870
rect 7120 16630 7290 16870
rect -5020 16540 7290 16630
rect -5020 16300 -4670 16540
rect -4430 16300 -4340 16540
rect -4100 16300 -4010 16540
rect -3770 16300 -3680 16540
rect -3440 16300 -3350 16540
rect -3110 16300 -3020 16540
rect -2780 16300 -2690 16540
rect -2450 16300 -2360 16540
rect -2120 16300 -2030 16540
rect -1790 16300 -1700 16540
rect -1460 16300 -1370 16540
rect -1130 16300 -1040 16540
rect -800 16300 -710 16540
rect -470 16300 -380 16540
rect -140 16300 -50 16540
rect 190 16300 280 16540
rect 520 16300 610 16540
rect 850 16300 940 16540
rect 1180 16300 1270 16540
rect 1510 16300 1600 16540
rect 1840 16300 1930 16540
rect 2170 16300 2260 16540
rect 2500 16300 2590 16540
rect 2830 16300 2920 16540
rect 3160 16300 3250 16540
rect 3490 16300 3580 16540
rect 3820 16300 3910 16540
rect 4150 16300 4240 16540
rect 4480 16300 4570 16540
rect 4810 16300 4900 16540
rect 5140 16300 5230 16540
rect 5470 16300 5560 16540
rect 5800 16300 5890 16540
rect 6130 16300 6220 16540
rect 6460 16300 6550 16540
rect 6790 16300 6880 16540
rect 7120 16300 7290 16540
rect -5020 16210 7290 16300
rect -5020 15970 -4670 16210
rect -4430 15970 -4340 16210
rect -4100 15970 -4010 16210
rect -3770 15970 -3680 16210
rect -3440 15970 -3350 16210
rect -3110 15970 -3020 16210
rect -2780 15970 -2690 16210
rect -2450 15970 -2360 16210
rect -2120 15970 -2030 16210
rect -1790 15970 -1700 16210
rect -1460 15970 -1370 16210
rect -1130 15970 -1040 16210
rect -800 15970 -710 16210
rect -470 15970 -380 16210
rect -140 15970 -50 16210
rect 190 15970 280 16210
rect 520 15970 610 16210
rect 850 15970 940 16210
rect 1180 15970 1270 16210
rect 1510 15970 1600 16210
rect 1840 15970 1930 16210
rect 2170 15970 2260 16210
rect 2500 15970 2590 16210
rect 2830 15970 2920 16210
rect 3160 15970 3250 16210
rect 3490 15970 3580 16210
rect 3820 15970 3910 16210
rect 4150 15970 4240 16210
rect 4480 15970 4570 16210
rect 4810 15970 4900 16210
rect 5140 15970 5230 16210
rect 5470 15970 5560 16210
rect 5800 15970 5890 16210
rect 6130 15970 6220 16210
rect 6460 15970 6550 16210
rect 6790 15970 6880 16210
rect 7120 15970 7290 16210
rect -5020 15880 7290 15970
rect -5020 15640 -4670 15880
rect -4430 15640 -4340 15880
rect -4100 15640 -4010 15880
rect -3770 15640 -3680 15880
rect -3440 15640 -3350 15880
rect -3110 15640 -3020 15880
rect -2780 15640 -2690 15880
rect -2450 15640 -2360 15880
rect -2120 15640 -2030 15880
rect -1790 15640 -1700 15880
rect -1460 15640 -1370 15880
rect -1130 15640 -1040 15880
rect -800 15640 -710 15880
rect -470 15640 -380 15880
rect -140 15640 -50 15880
rect 190 15640 280 15880
rect 520 15640 610 15880
rect 850 15640 940 15880
rect 1180 15640 1270 15880
rect 1510 15640 1600 15880
rect 1840 15640 1930 15880
rect 2170 15640 2260 15880
rect 2500 15640 2590 15880
rect 2830 15640 2920 15880
rect 3160 15640 3250 15880
rect 3490 15640 3580 15880
rect 3820 15640 3910 15880
rect 4150 15640 4240 15880
rect 4480 15640 4570 15880
rect 4810 15640 4900 15880
rect 5140 15640 5230 15880
rect 5470 15640 5560 15880
rect 5800 15640 5890 15880
rect 6130 15640 6220 15880
rect 6460 15640 6550 15880
rect 6790 15640 6880 15880
rect 7120 15640 7290 15880
rect -5020 15550 7290 15640
rect -5020 15310 -4670 15550
rect -4430 15310 -4340 15550
rect -4100 15310 -4010 15550
rect -3770 15310 -3680 15550
rect -3440 15310 -3350 15550
rect -3110 15310 -3020 15550
rect -2780 15310 -2690 15550
rect -2450 15310 -2360 15550
rect -2120 15310 -2030 15550
rect -1790 15310 -1700 15550
rect -1460 15310 -1370 15550
rect -1130 15310 -1040 15550
rect -800 15310 -710 15550
rect -470 15310 -380 15550
rect -140 15310 -50 15550
rect 190 15310 280 15550
rect 520 15310 610 15550
rect 850 15310 940 15550
rect 1180 15310 1270 15550
rect 1510 15310 1600 15550
rect 1840 15310 1930 15550
rect 2170 15310 2260 15550
rect 2500 15310 2590 15550
rect 2830 15310 2920 15550
rect 3160 15310 3250 15550
rect 3490 15310 3580 15550
rect 3820 15310 3910 15550
rect 4150 15310 4240 15550
rect 4480 15310 4570 15550
rect 4810 15310 4900 15550
rect 5140 15310 5230 15550
rect 5470 15310 5560 15550
rect 5800 15310 5890 15550
rect 6130 15310 6220 15550
rect 6460 15310 6550 15550
rect 6790 15310 6880 15550
rect 7120 15310 7290 15550
rect -5020 15220 7290 15310
rect -5020 14980 -4670 15220
rect -4430 14980 -4340 15220
rect -4100 14980 -4010 15220
rect -3770 14980 -3680 15220
rect -3440 14980 -3350 15220
rect -3110 14980 -3020 15220
rect -2780 14980 -2690 15220
rect -2450 14980 -2360 15220
rect -2120 14980 -2030 15220
rect -1790 14980 -1700 15220
rect -1460 14980 -1370 15220
rect -1130 14980 -1040 15220
rect -800 14980 -710 15220
rect -470 14980 -380 15220
rect -140 14980 -50 15220
rect 190 14980 280 15220
rect 520 14980 610 15220
rect 850 14980 940 15220
rect 1180 14980 1270 15220
rect 1510 14980 1600 15220
rect 1840 14980 1930 15220
rect 2170 14980 2260 15220
rect 2500 14980 2590 15220
rect 2830 14980 2920 15220
rect 3160 14980 3250 15220
rect 3490 14980 3580 15220
rect 3820 14980 3910 15220
rect 4150 14980 4240 15220
rect 4480 14980 4570 15220
rect 4810 14980 4900 15220
rect 5140 14980 5230 15220
rect 5470 14980 5560 15220
rect 5800 14980 5890 15220
rect 6130 14980 6220 15220
rect 6460 14980 6550 15220
rect 6790 14980 6880 15220
rect 7120 14980 7290 15220
rect -5020 14890 7290 14980
rect -5020 14650 -4670 14890
rect -4430 14650 -4340 14890
rect -4100 14650 -4010 14890
rect -3770 14650 -3680 14890
rect -3440 14650 -3350 14890
rect -3110 14650 -3020 14890
rect -2780 14650 -2690 14890
rect -2450 14650 -2360 14890
rect -2120 14650 -2030 14890
rect -1790 14650 -1700 14890
rect -1460 14650 -1370 14890
rect -1130 14650 -1040 14890
rect -800 14650 -710 14890
rect -470 14650 -380 14890
rect -140 14650 -50 14890
rect 190 14650 280 14890
rect 520 14650 610 14890
rect 850 14650 940 14890
rect 1180 14650 1270 14890
rect 1510 14650 1600 14890
rect 1840 14650 1930 14890
rect 2170 14650 2260 14890
rect 2500 14650 2590 14890
rect 2830 14650 2920 14890
rect 3160 14650 3250 14890
rect 3490 14650 3580 14890
rect 3820 14650 3910 14890
rect 4150 14650 4240 14890
rect 4480 14650 4570 14890
rect 4810 14650 4900 14890
rect 5140 14650 5230 14890
rect 5470 14650 5560 14890
rect 5800 14650 5890 14890
rect 6130 14650 6220 14890
rect 6460 14650 6550 14890
rect 6790 14650 6880 14890
rect 7120 14650 7290 14890
rect -5020 14560 7290 14650
rect -5020 14320 -4670 14560
rect -4430 14320 -4340 14560
rect -4100 14320 -4010 14560
rect -3770 14320 -3680 14560
rect -3440 14320 -3350 14560
rect -3110 14320 -3020 14560
rect -2780 14320 -2690 14560
rect -2450 14320 -2360 14560
rect -2120 14320 -2030 14560
rect -1790 14320 -1700 14560
rect -1460 14320 -1370 14560
rect -1130 14320 -1040 14560
rect -800 14320 -710 14560
rect -470 14320 -380 14560
rect -140 14320 -50 14560
rect 190 14320 280 14560
rect 520 14320 610 14560
rect 850 14320 940 14560
rect 1180 14320 1270 14560
rect 1510 14320 1600 14560
rect 1840 14320 1930 14560
rect 2170 14320 2260 14560
rect 2500 14320 2590 14560
rect 2830 14320 2920 14560
rect 3160 14320 3250 14560
rect 3490 14320 3580 14560
rect 3820 14320 3910 14560
rect 4150 14320 4240 14560
rect 4480 14320 4570 14560
rect 4810 14320 4900 14560
rect 5140 14320 5230 14560
rect 5470 14320 5560 14560
rect 5800 14320 5890 14560
rect 6130 14320 6220 14560
rect 6460 14320 6550 14560
rect 6790 14320 6880 14560
rect 7120 14320 7290 14560
rect -5020 14230 7290 14320
rect -5020 13990 -4670 14230
rect -4430 13990 -4340 14230
rect -4100 13990 -4010 14230
rect -3770 13990 -3680 14230
rect -3440 13990 -3350 14230
rect -3110 13990 -3020 14230
rect -2780 13990 -2690 14230
rect -2450 13990 -2360 14230
rect -2120 13990 -2030 14230
rect -1790 13990 -1700 14230
rect -1460 13990 -1370 14230
rect -1130 13990 -1040 14230
rect -800 13990 -710 14230
rect -470 13990 -380 14230
rect -140 13990 -50 14230
rect 190 13990 280 14230
rect 520 13990 610 14230
rect 850 13990 940 14230
rect 1180 13990 1270 14230
rect 1510 13990 1600 14230
rect 1840 13990 1930 14230
rect 2170 13990 2260 14230
rect 2500 13990 2590 14230
rect 2830 13990 2920 14230
rect 3160 13990 3250 14230
rect 3490 13990 3580 14230
rect 3820 13990 3910 14230
rect 4150 13990 4240 14230
rect 4480 13990 4570 14230
rect 4810 13990 4900 14230
rect 5140 13990 5230 14230
rect 5470 13990 5560 14230
rect 5800 13990 5890 14230
rect 6130 13990 6220 14230
rect 6460 13990 6550 14230
rect 6790 13990 6880 14230
rect 7120 13990 7290 14230
rect -5020 13900 7290 13990
rect -5020 13660 -4670 13900
rect -4430 13660 -4340 13900
rect -4100 13660 -4010 13900
rect -3770 13660 -3680 13900
rect -3440 13660 -3350 13900
rect -3110 13660 -3020 13900
rect -2780 13660 -2690 13900
rect -2450 13660 -2360 13900
rect -2120 13660 -2030 13900
rect -1790 13660 -1700 13900
rect -1460 13660 -1370 13900
rect -1130 13660 -1040 13900
rect -800 13660 -710 13900
rect -470 13660 -380 13900
rect -140 13660 -50 13900
rect 190 13660 280 13900
rect 520 13660 610 13900
rect 850 13660 940 13900
rect 1180 13660 1270 13900
rect 1510 13660 1600 13900
rect 1840 13660 1930 13900
rect 2170 13660 2260 13900
rect 2500 13660 2590 13900
rect 2830 13660 2920 13900
rect 3160 13660 3250 13900
rect 3490 13660 3580 13900
rect 3820 13660 3910 13900
rect 4150 13660 4240 13900
rect 4480 13660 4570 13900
rect 4810 13660 4900 13900
rect 5140 13660 5230 13900
rect 5470 13660 5560 13900
rect 5800 13660 5890 13900
rect 6130 13660 6220 13900
rect 6460 13660 6550 13900
rect 6790 13660 6880 13900
rect 7120 13660 7290 13900
rect -5020 13570 7290 13660
rect -5020 13330 -4670 13570
rect -4430 13330 -4340 13570
rect -4100 13330 -4010 13570
rect -3770 13330 -3680 13570
rect -3440 13330 -3350 13570
rect -3110 13330 -3020 13570
rect -2780 13330 -2690 13570
rect -2450 13330 -2360 13570
rect -2120 13330 -2030 13570
rect -1790 13330 -1700 13570
rect -1460 13330 -1370 13570
rect -1130 13330 -1040 13570
rect -800 13330 -710 13570
rect -470 13330 -380 13570
rect -140 13330 -50 13570
rect 190 13330 280 13570
rect 520 13330 610 13570
rect 850 13330 940 13570
rect 1180 13330 1270 13570
rect 1510 13330 1600 13570
rect 1840 13330 1930 13570
rect 2170 13330 2260 13570
rect 2500 13330 2590 13570
rect 2830 13330 2920 13570
rect 3160 13330 3250 13570
rect 3490 13330 3580 13570
rect 3820 13330 3910 13570
rect 4150 13330 4240 13570
rect 4480 13330 4570 13570
rect 4810 13330 4900 13570
rect 5140 13330 5230 13570
rect 5470 13330 5560 13570
rect 5800 13330 5890 13570
rect 6130 13330 6220 13570
rect 6460 13330 6550 13570
rect 6790 13330 6880 13570
rect 7120 13330 7290 13570
rect -5020 13240 7290 13330
rect -5020 13000 -4670 13240
rect -4430 13000 -4340 13240
rect -4100 13000 -4010 13240
rect -3770 13000 -3680 13240
rect -3440 13000 -3350 13240
rect -3110 13000 -3020 13240
rect -2780 13000 -2690 13240
rect -2450 13000 -2360 13240
rect -2120 13000 -2030 13240
rect -1790 13000 -1700 13240
rect -1460 13000 -1370 13240
rect -1130 13000 -1040 13240
rect -800 13000 -710 13240
rect -470 13000 -380 13240
rect -140 13000 -50 13240
rect 190 13000 280 13240
rect 520 13000 610 13240
rect 850 13000 940 13240
rect 1180 13000 1270 13240
rect 1510 13000 1600 13240
rect 1840 13000 1930 13240
rect 2170 13000 2260 13240
rect 2500 13000 2590 13240
rect 2830 13000 2920 13240
rect 3160 13000 3250 13240
rect 3490 13000 3580 13240
rect 3820 13000 3910 13240
rect 4150 13000 4240 13240
rect 4480 13000 4570 13240
rect 4810 13000 4900 13240
rect 5140 13000 5230 13240
rect 5470 13000 5560 13240
rect 5800 13000 5890 13240
rect 6130 13000 6220 13240
rect 6460 13000 6550 13240
rect 6790 13000 6880 13240
rect 7120 13000 7290 13240
rect -5020 12910 7290 13000
rect -5020 12670 -4670 12910
rect -4430 12670 -4340 12910
rect -4100 12670 -4010 12910
rect -3770 12670 -3680 12910
rect -3440 12670 -3350 12910
rect -3110 12670 -3020 12910
rect -2780 12670 -2690 12910
rect -2450 12670 -2360 12910
rect -2120 12670 -2030 12910
rect -1790 12670 -1700 12910
rect -1460 12670 -1370 12910
rect -1130 12670 -1040 12910
rect -800 12670 -710 12910
rect -470 12670 -380 12910
rect -140 12670 -50 12910
rect 190 12670 280 12910
rect 520 12670 610 12910
rect 850 12670 940 12910
rect 1180 12670 1270 12910
rect 1510 12670 1600 12910
rect 1840 12670 1930 12910
rect 2170 12670 2260 12910
rect 2500 12670 2590 12910
rect 2830 12670 2920 12910
rect 3160 12670 3250 12910
rect 3490 12670 3580 12910
rect 3820 12670 3910 12910
rect 4150 12670 4240 12910
rect 4480 12670 4570 12910
rect 4810 12670 4900 12910
rect 5140 12670 5230 12910
rect 5470 12670 5560 12910
rect 5800 12670 5890 12910
rect 6130 12670 6220 12910
rect 6460 12670 6550 12910
rect 6790 12670 6880 12910
rect 7120 12670 7290 12910
rect -5020 12580 7290 12670
rect -5020 12340 -4670 12580
rect -4430 12340 -4340 12580
rect -4100 12340 -4010 12580
rect -3770 12340 -3680 12580
rect -3440 12340 -3350 12580
rect -3110 12340 -3020 12580
rect -2780 12340 -2690 12580
rect -2450 12340 -2360 12580
rect -2120 12340 -2030 12580
rect -1790 12340 -1700 12580
rect -1460 12340 -1370 12580
rect -1130 12340 -1040 12580
rect -800 12340 -710 12580
rect -470 12340 -380 12580
rect -140 12340 -50 12580
rect 190 12340 280 12580
rect 520 12340 610 12580
rect 850 12340 940 12580
rect 1180 12340 1270 12580
rect 1510 12340 1600 12580
rect 1840 12340 1930 12580
rect 2170 12340 2260 12580
rect 2500 12340 2590 12580
rect 2830 12340 2920 12580
rect 3160 12340 3250 12580
rect 3490 12340 3580 12580
rect 3820 12340 3910 12580
rect 4150 12340 4240 12580
rect 4480 12340 4570 12580
rect 4810 12340 4900 12580
rect 5140 12340 5230 12580
rect 5470 12340 5560 12580
rect 5800 12340 5890 12580
rect 6130 12340 6220 12580
rect 6460 12340 6550 12580
rect 6790 12340 6880 12580
rect 7120 12340 7290 12580
rect -5020 12250 7290 12340
rect -5020 12010 -4670 12250
rect -4430 12010 -4340 12250
rect -4100 12010 -4010 12250
rect -3770 12010 -3680 12250
rect -3440 12010 -3350 12250
rect -3110 12010 -3020 12250
rect -2780 12010 -2690 12250
rect -2450 12010 -2360 12250
rect -2120 12010 -2030 12250
rect -1790 12010 -1700 12250
rect -1460 12010 -1370 12250
rect -1130 12010 -1040 12250
rect -800 12010 -710 12250
rect -470 12010 -380 12250
rect -140 12010 -50 12250
rect 190 12010 280 12250
rect 520 12010 610 12250
rect 850 12010 940 12250
rect 1180 12010 1270 12250
rect 1510 12010 1600 12250
rect 1840 12010 1930 12250
rect 2170 12010 2260 12250
rect 2500 12010 2590 12250
rect 2830 12010 2920 12250
rect 3160 12010 3250 12250
rect 3490 12010 3580 12250
rect 3820 12010 3910 12250
rect 4150 12010 4240 12250
rect 4480 12010 4570 12250
rect 4810 12010 4900 12250
rect 5140 12010 5230 12250
rect 5470 12010 5560 12250
rect 5800 12010 5890 12250
rect 6130 12010 6220 12250
rect 6460 12010 6550 12250
rect 6790 12010 6880 12250
rect 7120 12010 7290 12250
rect -5020 11920 7290 12010
rect -5020 11680 -4670 11920
rect -4430 11680 -4340 11920
rect -4100 11680 -4010 11920
rect -3770 11680 -3680 11920
rect -3440 11680 -3350 11920
rect -3110 11680 -3020 11920
rect -2780 11680 -2690 11920
rect -2450 11680 -2360 11920
rect -2120 11680 -2030 11920
rect -1790 11680 -1700 11920
rect -1460 11680 -1370 11920
rect -1130 11680 -1040 11920
rect -800 11680 -710 11920
rect -470 11680 -380 11920
rect -140 11680 -50 11920
rect 190 11680 280 11920
rect 520 11680 610 11920
rect 850 11680 940 11920
rect 1180 11680 1270 11920
rect 1510 11680 1600 11920
rect 1840 11680 1930 11920
rect 2170 11680 2260 11920
rect 2500 11680 2590 11920
rect 2830 11680 2920 11920
rect 3160 11680 3250 11920
rect 3490 11680 3580 11920
rect 3820 11680 3910 11920
rect 4150 11680 4240 11920
rect 4480 11680 4570 11920
rect 4810 11680 4900 11920
rect 5140 11680 5230 11920
rect 5470 11680 5560 11920
rect 5800 11680 5890 11920
rect 6130 11680 6220 11920
rect 6460 11680 6550 11920
rect 6790 11680 6880 11920
rect 7120 11680 7290 11920
rect -5020 11590 7290 11680
rect -5020 11350 -4670 11590
rect -4430 11350 -4340 11590
rect -4100 11350 -4010 11590
rect -3770 11350 -3680 11590
rect -3440 11350 -3350 11590
rect -3110 11350 -3020 11590
rect -2780 11350 -2690 11590
rect -2450 11350 -2360 11590
rect -2120 11350 -2030 11590
rect -1790 11350 -1700 11590
rect -1460 11350 -1370 11590
rect -1130 11350 -1040 11590
rect -800 11350 -710 11590
rect -470 11350 -380 11590
rect -140 11350 -50 11590
rect 190 11350 280 11590
rect 520 11350 610 11590
rect 850 11350 940 11590
rect 1180 11350 1270 11590
rect 1510 11350 1600 11590
rect 1840 11350 1930 11590
rect 2170 11350 2260 11590
rect 2500 11350 2590 11590
rect 2830 11350 2920 11590
rect 3160 11350 3250 11590
rect 3490 11350 3580 11590
rect 3820 11350 3910 11590
rect 4150 11350 4240 11590
rect 4480 11350 4570 11590
rect 4810 11350 4900 11590
rect 5140 11350 5230 11590
rect 5470 11350 5560 11590
rect 5800 11350 5890 11590
rect 6130 11350 6220 11590
rect 6460 11350 6550 11590
rect 6790 11350 6880 11590
rect 7120 11350 7290 11590
rect -5020 11260 7290 11350
rect -5020 11020 -4670 11260
rect -4430 11020 -4340 11260
rect -4100 11020 -4010 11260
rect -3770 11020 -3680 11260
rect -3440 11020 -3350 11260
rect -3110 11020 -3020 11260
rect -2780 11020 -2690 11260
rect -2450 11020 -2360 11260
rect -2120 11020 -2030 11260
rect -1790 11020 -1700 11260
rect -1460 11020 -1370 11260
rect -1130 11020 -1040 11260
rect -800 11020 -710 11260
rect -470 11020 -380 11260
rect -140 11020 -50 11260
rect 190 11020 280 11260
rect 520 11020 610 11260
rect 850 11020 940 11260
rect 1180 11020 1270 11260
rect 1510 11020 1600 11260
rect 1840 11020 1930 11260
rect 2170 11020 2260 11260
rect 2500 11020 2590 11260
rect 2830 11020 2920 11260
rect 3160 11020 3250 11260
rect 3490 11020 3580 11260
rect 3820 11020 3910 11260
rect 4150 11020 4240 11260
rect 4480 11020 4570 11260
rect 4810 11020 4900 11260
rect 5140 11020 5230 11260
rect 5470 11020 5560 11260
rect 5800 11020 5890 11260
rect 6130 11020 6220 11260
rect 6460 11020 6550 11260
rect 6790 11020 6880 11260
rect 7120 11020 7290 11260
rect -5020 10930 7290 11020
rect -5020 10690 -4670 10930
rect -4430 10690 -4340 10930
rect -4100 10690 -4010 10930
rect -3770 10690 -3680 10930
rect -3440 10690 -3350 10930
rect -3110 10690 -3020 10930
rect -2780 10690 -2690 10930
rect -2450 10690 -2360 10930
rect -2120 10690 -2030 10930
rect -1790 10690 -1700 10930
rect -1460 10690 -1370 10930
rect -1130 10690 -1040 10930
rect -800 10690 -710 10930
rect -470 10690 -380 10930
rect -140 10690 -50 10930
rect 190 10690 280 10930
rect 520 10690 610 10930
rect 850 10690 940 10930
rect 1180 10690 1270 10930
rect 1510 10690 1600 10930
rect 1840 10690 1930 10930
rect 2170 10690 2260 10930
rect 2500 10690 2590 10930
rect 2830 10690 2920 10930
rect 3160 10690 3250 10930
rect 3490 10690 3580 10930
rect 3820 10690 3910 10930
rect 4150 10690 4240 10930
rect 4480 10690 4570 10930
rect 4810 10690 4900 10930
rect 5140 10690 5230 10930
rect 5470 10690 5560 10930
rect 5800 10690 5890 10930
rect 6130 10690 6220 10930
rect 6460 10690 6550 10930
rect 6790 10690 6880 10930
rect 7120 10690 7290 10930
rect -5020 10600 7290 10690
rect -5020 10360 -4670 10600
rect -4430 10360 -4340 10600
rect -4100 10360 -4010 10600
rect -3770 10360 -3680 10600
rect -3440 10360 -3350 10600
rect -3110 10360 -3020 10600
rect -2780 10360 -2690 10600
rect -2450 10360 -2360 10600
rect -2120 10360 -2030 10600
rect -1790 10360 -1700 10600
rect -1460 10360 -1370 10600
rect -1130 10360 -1040 10600
rect -800 10360 -710 10600
rect -470 10360 -380 10600
rect -140 10360 -50 10600
rect 190 10360 280 10600
rect 520 10360 610 10600
rect 850 10360 940 10600
rect 1180 10360 1270 10600
rect 1510 10360 1600 10600
rect 1840 10360 1930 10600
rect 2170 10360 2260 10600
rect 2500 10360 2590 10600
rect 2830 10360 2920 10600
rect 3160 10360 3250 10600
rect 3490 10360 3580 10600
rect 3820 10360 3910 10600
rect 4150 10360 4240 10600
rect 4480 10360 4570 10600
rect 4810 10360 4900 10600
rect 5140 10360 5230 10600
rect 5470 10360 5560 10600
rect 5800 10360 5890 10600
rect 6130 10360 6220 10600
rect 6460 10360 6550 10600
rect 6790 10360 6880 10600
rect 7120 10360 7290 10600
rect -5020 10270 7290 10360
rect -5020 10030 -4670 10270
rect -4430 10030 -4340 10270
rect -4100 10030 -4010 10270
rect -3770 10030 -3680 10270
rect -3440 10030 -3350 10270
rect -3110 10030 -3020 10270
rect -2780 10030 -2690 10270
rect -2450 10030 -2360 10270
rect -2120 10030 -2030 10270
rect -1790 10030 -1700 10270
rect -1460 10030 -1370 10270
rect -1130 10030 -1040 10270
rect -800 10030 -710 10270
rect -470 10030 -380 10270
rect -140 10030 -50 10270
rect 190 10030 280 10270
rect 520 10030 610 10270
rect 850 10030 940 10270
rect 1180 10030 1270 10270
rect 1510 10030 1600 10270
rect 1840 10030 1930 10270
rect 2170 10030 2260 10270
rect 2500 10030 2590 10270
rect 2830 10030 2920 10270
rect 3160 10030 3250 10270
rect 3490 10030 3580 10270
rect 3820 10030 3910 10270
rect 4150 10030 4240 10270
rect 4480 10030 4570 10270
rect 4810 10030 4900 10270
rect 5140 10030 5230 10270
rect 5470 10030 5560 10270
rect 5800 10030 5890 10270
rect 6130 10030 6220 10270
rect 6460 10030 6550 10270
rect 6790 10030 6880 10270
rect 7120 10030 7290 10270
rect -5020 9940 7290 10030
rect -5020 9700 -4670 9940
rect -4430 9700 -4340 9940
rect -4100 9700 -4010 9940
rect -3770 9700 -3680 9940
rect -3440 9700 -3350 9940
rect -3110 9700 -3020 9940
rect -2780 9700 -2690 9940
rect -2450 9700 -2360 9940
rect -2120 9700 -2030 9940
rect -1790 9700 -1700 9940
rect -1460 9700 -1370 9940
rect -1130 9700 -1040 9940
rect -800 9700 -710 9940
rect -470 9700 -380 9940
rect -140 9700 -50 9940
rect 190 9700 280 9940
rect 520 9700 610 9940
rect 850 9700 940 9940
rect 1180 9700 1270 9940
rect 1510 9700 1600 9940
rect 1840 9700 1930 9940
rect 2170 9700 2260 9940
rect 2500 9700 2590 9940
rect 2830 9700 2920 9940
rect 3160 9700 3250 9940
rect 3490 9700 3580 9940
rect 3820 9700 3910 9940
rect 4150 9700 4240 9940
rect 4480 9700 4570 9940
rect 4810 9700 4900 9940
rect 5140 9700 5230 9940
rect 5470 9700 5560 9940
rect 5800 9700 5890 9940
rect 6130 9700 6220 9940
rect 6460 9700 6550 9940
rect 6790 9700 6880 9940
rect 7120 9700 7290 9940
rect -5020 9610 7290 9700
rect -5020 9370 -4670 9610
rect -4430 9370 -4340 9610
rect -4100 9370 -4010 9610
rect -3770 9370 -3680 9610
rect -3440 9370 -3350 9610
rect -3110 9370 -3020 9610
rect -2780 9370 -2690 9610
rect -2450 9370 -2360 9610
rect -2120 9370 -2030 9610
rect -1790 9370 -1700 9610
rect -1460 9370 -1370 9610
rect -1130 9370 -1040 9610
rect -800 9370 -710 9610
rect -470 9370 -380 9610
rect -140 9370 -50 9610
rect 190 9370 280 9610
rect 520 9370 610 9610
rect 850 9370 940 9610
rect 1180 9370 1270 9610
rect 1510 9370 1600 9610
rect 1840 9370 1930 9610
rect 2170 9370 2260 9610
rect 2500 9370 2590 9610
rect 2830 9370 2920 9610
rect 3160 9370 3250 9610
rect 3490 9370 3580 9610
rect 3820 9370 3910 9610
rect 4150 9370 4240 9610
rect 4480 9370 4570 9610
rect 4810 9370 4900 9610
rect 5140 9370 5230 9610
rect 5470 9370 5560 9610
rect 5800 9370 5890 9610
rect 6130 9370 6220 9610
rect 6460 9370 6550 9610
rect 6790 9370 6880 9610
rect 7120 9370 7290 9610
rect -5020 9280 7290 9370
rect -5020 9040 -4670 9280
rect -4430 9040 -4340 9280
rect -4100 9040 -4010 9280
rect -3770 9040 -3680 9280
rect -3440 9040 -3350 9280
rect -3110 9040 -3020 9280
rect -2780 9040 -2690 9280
rect -2450 9040 -2360 9280
rect -2120 9040 -2030 9280
rect -1790 9040 -1700 9280
rect -1460 9040 -1370 9280
rect -1130 9040 -1040 9280
rect -800 9040 -710 9280
rect -470 9040 -380 9280
rect -140 9040 -50 9280
rect 190 9040 280 9280
rect 520 9040 610 9280
rect 850 9040 940 9280
rect 1180 9040 1270 9280
rect 1510 9040 1600 9280
rect 1840 9040 1930 9280
rect 2170 9040 2260 9280
rect 2500 9040 2590 9280
rect 2830 9040 2920 9280
rect 3160 9040 3250 9280
rect 3490 9040 3580 9280
rect 3820 9040 3910 9280
rect 4150 9040 4240 9280
rect 4480 9040 4570 9280
rect 4810 9040 4900 9280
rect 5140 9040 5230 9280
rect 5470 9040 5560 9280
rect 5800 9040 5890 9280
rect 6130 9040 6220 9280
rect 6460 9040 6550 9280
rect 6790 9040 6880 9280
rect 7120 9040 7290 9280
rect -5020 8690 7290 9040
rect 7020 8410 7290 8690
rect 7020 8340 7040 8410
rect 7140 8340 7170 8410
rect 7270 8340 7290 8410
rect 7020 8320 7290 8340
rect 7020 8250 7040 8320
rect 7140 8250 7170 8320
rect 7270 8250 7290 8320
rect 7020 8230 7290 8250
rect 7610 20830 19920 21000
rect 7610 20590 7780 20830
rect 8020 20590 8110 20830
rect 8350 20590 8440 20830
rect 8680 20590 8770 20830
rect 9010 20590 9100 20830
rect 9340 20590 9430 20830
rect 9670 20590 9760 20830
rect 10000 20590 10090 20830
rect 10330 20590 10420 20830
rect 10660 20590 10750 20830
rect 10990 20590 11080 20830
rect 11320 20590 11410 20830
rect 11650 20590 11740 20830
rect 11980 20590 12070 20830
rect 12310 20590 12400 20830
rect 12640 20590 12730 20830
rect 12970 20590 13060 20830
rect 13300 20590 13390 20830
rect 13630 20590 13720 20830
rect 13960 20590 14050 20830
rect 14290 20590 14380 20830
rect 14620 20590 14710 20830
rect 14950 20590 15040 20830
rect 15280 20590 15370 20830
rect 15610 20590 15700 20830
rect 15940 20590 16030 20830
rect 16270 20590 16360 20830
rect 16600 20590 16690 20830
rect 16930 20590 17020 20830
rect 17260 20590 17350 20830
rect 17590 20590 17680 20830
rect 17920 20590 18010 20830
rect 18250 20590 18340 20830
rect 18580 20590 18670 20830
rect 18910 20590 19000 20830
rect 19240 20590 19330 20830
rect 19570 20590 19920 20830
rect 7610 20500 19920 20590
rect 7610 20260 7780 20500
rect 8020 20260 8110 20500
rect 8350 20260 8440 20500
rect 8680 20260 8770 20500
rect 9010 20260 9100 20500
rect 9340 20260 9430 20500
rect 9670 20260 9760 20500
rect 10000 20260 10090 20500
rect 10330 20260 10420 20500
rect 10660 20260 10750 20500
rect 10990 20260 11080 20500
rect 11320 20260 11410 20500
rect 11650 20260 11740 20500
rect 11980 20260 12070 20500
rect 12310 20260 12400 20500
rect 12640 20260 12730 20500
rect 12970 20260 13060 20500
rect 13300 20260 13390 20500
rect 13630 20260 13720 20500
rect 13960 20260 14050 20500
rect 14290 20260 14380 20500
rect 14620 20260 14710 20500
rect 14950 20260 15040 20500
rect 15280 20260 15370 20500
rect 15610 20260 15700 20500
rect 15940 20260 16030 20500
rect 16270 20260 16360 20500
rect 16600 20260 16690 20500
rect 16930 20260 17020 20500
rect 17260 20260 17350 20500
rect 17590 20260 17680 20500
rect 17920 20260 18010 20500
rect 18250 20260 18340 20500
rect 18580 20260 18670 20500
rect 18910 20260 19000 20500
rect 19240 20260 19330 20500
rect 19570 20260 19920 20500
rect 7610 20170 19920 20260
rect 7610 19930 7780 20170
rect 8020 19930 8110 20170
rect 8350 19930 8440 20170
rect 8680 19930 8770 20170
rect 9010 19930 9100 20170
rect 9340 19930 9430 20170
rect 9670 19930 9760 20170
rect 10000 19930 10090 20170
rect 10330 19930 10420 20170
rect 10660 19930 10750 20170
rect 10990 19930 11080 20170
rect 11320 19930 11410 20170
rect 11650 19930 11740 20170
rect 11980 19930 12070 20170
rect 12310 19930 12400 20170
rect 12640 19930 12730 20170
rect 12970 19930 13060 20170
rect 13300 19930 13390 20170
rect 13630 19930 13720 20170
rect 13960 19930 14050 20170
rect 14290 19930 14380 20170
rect 14620 19930 14710 20170
rect 14950 19930 15040 20170
rect 15280 19930 15370 20170
rect 15610 19930 15700 20170
rect 15940 19930 16030 20170
rect 16270 19930 16360 20170
rect 16600 19930 16690 20170
rect 16930 19930 17020 20170
rect 17260 19930 17350 20170
rect 17590 19930 17680 20170
rect 17920 19930 18010 20170
rect 18250 19930 18340 20170
rect 18580 19930 18670 20170
rect 18910 19930 19000 20170
rect 19240 19930 19330 20170
rect 19570 19930 19920 20170
rect 7610 19840 19920 19930
rect 7610 19600 7780 19840
rect 8020 19600 8110 19840
rect 8350 19600 8440 19840
rect 8680 19600 8770 19840
rect 9010 19600 9100 19840
rect 9340 19600 9430 19840
rect 9670 19600 9760 19840
rect 10000 19600 10090 19840
rect 10330 19600 10420 19840
rect 10660 19600 10750 19840
rect 10990 19600 11080 19840
rect 11320 19600 11410 19840
rect 11650 19600 11740 19840
rect 11980 19600 12070 19840
rect 12310 19600 12400 19840
rect 12640 19600 12730 19840
rect 12970 19600 13060 19840
rect 13300 19600 13390 19840
rect 13630 19600 13720 19840
rect 13960 19600 14050 19840
rect 14290 19600 14380 19840
rect 14620 19600 14710 19840
rect 14950 19600 15040 19840
rect 15280 19600 15370 19840
rect 15610 19600 15700 19840
rect 15940 19600 16030 19840
rect 16270 19600 16360 19840
rect 16600 19600 16690 19840
rect 16930 19600 17020 19840
rect 17260 19600 17350 19840
rect 17590 19600 17680 19840
rect 17920 19600 18010 19840
rect 18250 19600 18340 19840
rect 18580 19600 18670 19840
rect 18910 19600 19000 19840
rect 19240 19600 19330 19840
rect 19570 19600 19920 19840
rect 7610 19510 19920 19600
rect 7610 19270 7780 19510
rect 8020 19270 8110 19510
rect 8350 19270 8440 19510
rect 8680 19270 8770 19510
rect 9010 19270 9100 19510
rect 9340 19270 9430 19510
rect 9670 19270 9760 19510
rect 10000 19270 10090 19510
rect 10330 19270 10420 19510
rect 10660 19270 10750 19510
rect 10990 19270 11080 19510
rect 11320 19270 11410 19510
rect 11650 19270 11740 19510
rect 11980 19270 12070 19510
rect 12310 19270 12400 19510
rect 12640 19270 12730 19510
rect 12970 19270 13060 19510
rect 13300 19270 13390 19510
rect 13630 19270 13720 19510
rect 13960 19270 14050 19510
rect 14290 19270 14380 19510
rect 14620 19270 14710 19510
rect 14950 19270 15040 19510
rect 15280 19270 15370 19510
rect 15610 19270 15700 19510
rect 15940 19270 16030 19510
rect 16270 19270 16360 19510
rect 16600 19270 16690 19510
rect 16930 19270 17020 19510
rect 17260 19270 17350 19510
rect 17590 19270 17680 19510
rect 17920 19270 18010 19510
rect 18250 19270 18340 19510
rect 18580 19270 18670 19510
rect 18910 19270 19000 19510
rect 19240 19270 19330 19510
rect 19570 19270 19920 19510
rect 7610 19180 19920 19270
rect 7610 18940 7780 19180
rect 8020 18940 8110 19180
rect 8350 18940 8440 19180
rect 8680 18940 8770 19180
rect 9010 18940 9100 19180
rect 9340 18940 9430 19180
rect 9670 18940 9760 19180
rect 10000 18940 10090 19180
rect 10330 18940 10420 19180
rect 10660 18940 10750 19180
rect 10990 18940 11080 19180
rect 11320 18940 11410 19180
rect 11650 18940 11740 19180
rect 11980 18940 12070 19180
rect 12310 18940 12400 19180
rect 12640 18940 12730 19180
rect 12970 18940 13060 19180
rect 13300 18940 13390 19180
rect 13630 18940 13720 19180
rect 13960 18940 14050 19180
rect 14290 18940 14380 19180
rect 14620 18940 14710 19180
rect 14950 18940 15040 19180
rect 15280 18940 15370 19180
rect 15610 18940 15700 19180
rect 15940 18940 16030 19180
rect 16270 18940 16360 19180
rect 16600 18940 16690 19180
rect 16930 18940 17020 19180
rect 17260 18940 17350 19180
rect 17590 18940 17680 19180
rect 17920 18940 18010 19180
rect 18250 18940 18340 19180
rect 18580 18940 18670 19180
rect 18910 18940 19000 19180
rect 19240 18940 19330 19180
rect 19570 18940 19920 19180
rect 7610 18850 19920 18940
rect 7610 18610 7780 18850
rect 8020 18610 8110 18850
rect 8350 18610 8440 18850
rect 8680 18610 8770 18850
rect 9010 18610 9100 18850
rect 9340 18610 9430 18850
rect 9670 18610 9760 18850
rect 10000 18610 10090 18850
rect 10330 18610 10420 18850
rect 10660 18610 10750 18850
rect 10990 18610 11080 18850
rect 11320 18610 11410 18850
rect 11650 18610 11740 18850
rect 11980 18610 12070 18850
rect 12310 18610 12400 18850
rect 12640 18610 12730 18850
rect 12970 18610 13060 18850
rect 13300 18610 13390 18850
rect 13630 18610 13720 18850
rect 13960 18610 14050 18850
rect 14290 18610 14380 18850
rect 14620 18610 14710 18850
rect 14950 18610 15040 18850
rect 15280 18610 15370 18850
rect 15610 18610 15700 18850
rect 15940 18610 16030 18850
rect 16270 18610 16360 18850
rect 16600 18610 16690 18850
rect 16930 18610 17020 18850
rect 17260 18610 17350 18850
rect 17590 18610 17680 18850
rect 17920 18610 18010 18850
rect 18250 18610 18340 18850
rect 18580 18610 18670 18850
rect 18910 18610 19000 18850
rect 19240 18610 19330 18850
rect 19570 18610 19920 18850
rect 7610 18520 19920 18610
rect 7610 18280 7780 18520
rect 8020 18280 8110 18520
rect 8350 18280 8440 18520
rect 8680 18280 8770 18520
rect 9010 18280 9100 18520
rect 9340 18280 9430 18520
rect 9670 18280 9760 18520
rect 10000 18280 10090 18520
rect 10330 18280 10420 18520
rect 10660 18280 10750 18520
rect 10990 18280 11080 18520
rect 11320 18280 11410 18520
rect 11650 18280 11740 18520
rect 11980 18280 12070 18520
rect 12310 18280 12400 18520
rect 12640 18280 12730 18520
rect 12970 18280 13060 18520
rect 13300 18280 13390 18520
rect 13630 18280 13720 18520
rect 13960 18280 14050 18520
rect 14290 18280 14380 18520
rect 14620 18280 14710 18520
rect 14950 18280 15040 18520
rect 15280 18280 15370 18520
rect 15610 18280 15700 18520
rect 15940 18280 16030 18520
rect 16270 18280 16360 18520
rect 16600 18280 16690 18520
rect 16930 18280 17020 18520
rect 17260 18280 17350 18520
rect 17590 18280 17680 18520
rect 17920 18280 18010 18520
rect 18250 18280 18340 18520
rect 18580 18280 18670 18520
rect 18910 18280 19000 18520
rect 19240 18280 19330 18520
rect 19570 18280 19920 18520
rect 7610 18190 19920 18280
rect 7610 17950 7780 18190
rect 8020 17950 8110 18190
rect 8350 17950 8440 18190
rect 8680 17950 8770 18190
rect 9010 17950 9100 18190
rect 9340 17950 9430 18190
rect 9670 17950 9760 18190
rect 10000 17950 10090 18190
rect 10330 17950 10420 18190
rect 10660 17950 10750 18190
rect 10990 17950 11080 18190
rect 11320 17950 11410 18190
rect 11650 17950 11740 18190
rect 11980 17950 12070 18190
rect 12310 17950 12400 18190
rect 12640 17950 12730 18190
rect 12970 17950 13060 18190
rect 13300 17950 13390 18190
rect 13630 17950 13720 18190
rect 13960 17950 14050 18190
rect 14290 17950 14380 18190
rect 14620 17950 14710 18190
rect 14950 17950 15040 18190
rect 15280 17950 15370 18190
rect 15610 17950 15700 18190
rect 15940 17950 16030 18190
rect 16270 17950 16360 18190
rect 16600 17950 16690 18190
rect 16930 17950 17020 18190
rect 17260 17950 17350 18190
rect 17590 17950 17680 18190
rect 17920 17950 18010 18190
rect 18250 17950 18340 18190
rect 18580 17950 18670 18190
rect 18910 17950 19000 18190
rect 19240 17950 19330 18190
rect 19570 17950 19920 18190
rect 7610 17860 19920 17950
rect 7610 17620 7780 17860
rect 8020 17620 8110 17860
rect 8350 17620 8440 17860
rect 8680 17620 8770 17860
rect 9010 17620 9100 17860
rect 9340 17620 9430 17860
rect 9670 17620 9760 17860
rect 10000 17620 10090 17860
rect 10330 17620 10420 17860
rect 10660 17620 10750 17860
rect 10990 17620 11080 17860
rect 11320 17620 11410 17860
rect 11650 17620 11740 17860
rect 11980 17620 12070 17860
rect 12310 17620 12400 17860
rect 12640 17620 12730 17860
rect 12970 17620 13060 17860
rect 13300 17620 13390 17860
rect 13630 17620 13720 17860
rect 13960 17620 14050 17860
rect 14290 17620 14380 17860
rect 14620 17620 14710 17860
rect 14950 17620 15040 17860
rect 15280 17620 15370 17860
rect 15610 17620 15700 17860
rect 15940 17620 16030 17860
rect 16270 17620 16360 17860
rect 16600 17620 16690 17860
rect 16930 17620 17020 17860
rect 17260 17620 17350 17860
rect 17590 17620 17680 17860
rect 17920 17620 18010 17860
rect 18250 17620 18340 17860
rect 18580 17620 18670 17860
rect 18910 17620 19000 17860
rect 19240 17620 19330 17860
rect 19570 17620 19920 17860
rect 7610 17530 19920 17620
rect 7610 17290 7780 17530
rect 8020 17290 8110 17530
rect 8350 17290 8440 17530
rect 8680 17290 8770 17530
rect 9010 17290 9100 17530
rect 9340 17290 9430 17530
rect 9670 17290 9760 17530
rect 10000 17290 10090 17530
rect 10330 17290 10420 17530
rect 10660 17290 10750 17530
rect 10990 17290 11080 17530
rect 11320 17290 11410 17530
rect 11650 17290 11740 17530
rect 11980 17290 12070 17530
rect 12310 17290 12400 17530
rect 12640 17290 12730 17530
rect 12970 17290 13060 17530
rect 13300 17290 13390 17530
rect 13630 17290 13720 17530
rect 13960 17290 14050 17530
rect 14290 17290 14380 17530
rect 14620 17290 14710 17530
rect 14950 17290 15040 17530
rect 15280 17290 15370 17530
rect 15610 17290 15700 17530
rect 15940 17290 16030 17530
rect 16270 17290 16360 17530
rect 16600 17290 16690 17530
rect 16930 17290 17020 17530
rect 17260 17290 17350 17530
rect 17590 17290 17680 17530
rect 17920 17290 18010 17530
rect 18250 17290 18340 17530
rect 18580 17290 18670 17530
rect 18910 17290 19000 17530
rect 19240 17290 19330 17530
rect 19570 17290 19920 17530
rect 7610 17200 19920 17290
rect 7610 16960 7780 17200
rect 8020 16960 8110 17200
rect 8350 16960 8440 17200
rect 8680 16960 8770 17200
rect 9010 16960 9100 17200
rect 9340 16960 9430 17200
rect 9670 16960 9760 17200
rect 10000 16960 10090 17200
rect 10330 16960 10420 17200
rect 10660 16960 10750 17200
rect 10990 16960 11080 17200
rect 11320 16960 11410 17200
rect 11650 16960 11740 17200
rect 11980 16960 12070 17200
rect 12310 16960 12400 17200
rect 12640 16960 12730 17200
rect 12970 16960 13060 17200
rect 13300 16960 13390 17200
rect 13630 16960 13720 17200
rect 13960 16960 14050 17200
rect 14290 16960 14380 17200
rect 14620 16960 14710 17200
rect 14950 16960 15040 17200
rect 15280 16960 15370 17200
rect 15610 16960 15700 17200
rect 15940 16960 16030 17200
rect 16270 16960 16360 17200
rect 16600 16960 16690 17200
rect 16930 16960 17020 17200
rect 17260 16960 17350 17200
rect 17590 16960 17680 17200
rect 17920 16960 18010 17200
rect 18250 16960 18340 17200
rect 18580 16960 18670 17200
rect 18910 16960 19000 17200
rect 19240 16960 19330 17200
rect 19570 16960 19920 17200
rect 7610 16870 19920 16960
rect 7610 16630 7780 16870
rect 8020 16630 8110 16870
rect 8350 16630 8440 16870
rect 8680 16630 8770 16870
rect 9010 16630 9100 16870
rect 9340 16630 9430 16870
rect 9670 16630 9760 16870
rect 10000 16630 10090 16870
rect 10330 16630 10420 16870
rect 10660 16630 10750 16870
rect 10990 16630 11080 16870
rect 11320 16630 11410 16870
rect 11650 16630 11740 16870
rect 11980 16630 12070 16870
rect 12310 16630 12400 16870
rect 12640 16630 12730 16870
rect 12970 16630 13060 16870
rect 13300 16630 13390 16870
rect 13630 16630 13720 16870
rect 13960 16630 14050 16870
rect 14290 16630 14380 16870
rect 14620 16630 14710 16870
rect 14950 16630 15040 16870
rect 15280 16630 15370 16870
rect 15610 16630 15700 16870
rect 15940 16630 16030 16870
rect 16270 16630 16360 16870
rect 16600 16630 16690 16870
rect 16930 16630 17020 16870
rect 17260 16630 17350 16870
rect 17590 16630 17680 16870
rect 17920 16630 18010 16870
rect 18250 16630 18340 16870
rect 18580 16630 18670 16870
rect 18910 16630 19000 16870
rect 19240 16630 19330 16870
rect 19570 16630 19920 16870
rect 7610 16540 19920 16630
rect 7610 16300 7780 16540
rect 8020 16300 8110 16540
rect 8350 16300 8440 16540
rect 8680 16300 8770 16540
rect 9010 16300 9100 16540
rect 9340 16300 9430 16540
rect 9670 16300 9760 16540
rect 10000 16300 10090 16540
rect 10330 16300 10420 16540
rect 10660 16300 10750 16540
rect 10990 16300 11080 16540
rect 11320 16300 11410 16540
rect 11650 16300 11740 16540
rect 11980 16300 12070 16540
rect 12310 16300 12400 16540
rect 12640 16300 12730 16540
rect 12970 16300 13060 16540
rect 13300 16300 13390 16540
rect 13630 16300 13720 16540
rect 13960 16300 14050 16540
rect 14290 16300 14380 16540
rect 14620 16300 14710 16540
rect 14950 16300 15040 16540
rect 15280 16300 15370 16540
rect 15610 16300 15700 16540
rect 15940 16300 16030 16540
rect 16270 16300 16360 16540
rect 16600 16300 16690 16540
rect 16930 16300 17020 16540
rect 17260 16300 17350 16540
rect 17590 16300 17680 16540
rect 17920 16300 18010 16540
rect 18250 16300 18340 16540
rect 18580 16300 18670 16540
rect 18910 16300 19000 16540
rect 19240 16300 19330 16540
rect 19570 16300 19920 16540
rect 7610 16210 19920 16300
rect 7610 15970 7780 16210
rect 8020 15970 8110 16210
rect 8350 15970 8440 16210
rect 8680 15970 8770 16210
rect 9010 15970 9100 16210
rect 9340 15970 9430 16210
rect 9670 15970 9760 16210
rect 10000 15970 10090 16210
rect 10330 15970 10420 16210
rect 10660 15970 10750 16210
rect 10990 15970 11080 16210
rect 11320 15970 11410 16210
rect 11650 15970 11740 16210
rect 11980 15970 12070 16210
rect 12310 15970 12400 16210
rect 12640 15970 12730 16210
rect 12970 15970 13060 16210
rect 13300 15970 13390 16210
rect 13630 15970 13720 16210
rect 13960 15970 14050 16210
rect 14290 15970 14380 16210
rect 14620 15970 14710 16210
rect 14950 15970 15040 16210
rect 15280 15970 15370 16210
rect 15610 15970 15700 16210
rect 15940 15970 16030 16210
rect 16270 15970 16360 16210
rect 16600 15970 16690 16210
rect 16930 15970 17020 16210
rect 17260 15970 17350 16210
rect 17590 15970 17680 16210
rect 17920 15970 18010 16210
rect 18250 15970 18340 16210
rect 18580 15970 18670 16210
rect 18910 15970 19000 16210
rect 19240 15970 19330 16210
rect 19570 15970 19920 16210
rect 7610 15880 19920 15970
rect 7610 15640 7780 15880
rect 8020 15640 8110 15880
rect 8350 15640 8440 15880
rect 8680 15640 8770 15880
rect 9010 15640 9100 15880
rect 9340 15640 9430 15880
rect 9670 15640 9760 15880
rect 10000 15640 10090 15880
rect 10330 15640 10420 15880
rect 10660 15640 10750 15880
rect 10990 15640 11080 15880
rect 11320 15640 11410 15880
rect 11650 15640 11740 15880
rect 11980 15640 12070 15880
rect 12310 15640 12400 15880
rect 12640 15640 12730 15880
rect 12970 15640 13060 15880
rect 13300 15640 13390 15880
rect 13630 15640 13720 15880
rect 13960 15640 14050 15880
rect 14290 15640 14380 15880
rect 14620 15640 14710 15880
rect 14950 15640 15040 15880
rect 15280 15640 15370 15880
rect 15610 15640 15700 15880
rect 15940 15640 16030 15880
rect 16270 15640 16360 15880
rect 16600 15640 16690 15880
rect 16930 15640 17020 15880
rect 17260 15640 17350 15880
rect 17590 15640 17680 15880
rect 17920 15640 18010 15880
rect 18250 15640 18340 15880
rect 18580 15640 18670 15880
rect 18910 15640 19000 15880
rect 19240 15640 19330 15880
rect 19570 15640 19920 15880
rect 7610 15550 19920 15640
rect 7610 15310 7780 15550
rect 8020 15310 8110 15550
rect 8350 15310 8440 15550
rect 8680 15310 8770 15550
rect 9010 15310 9100 15550
rect 9340 15310 9430 15550
rect 9670 15310 9760 15550
rect 10000 15310 10090 15550
rect 10330 15310 10420 15550
rect 10660 15310 10750 15550
rect 10990 15310 11080 15550
rect 11320 15310 11410 15550
rect 11650 15310 11740 15550
rect 11980 15310 12070 15550
rect 12310 15310 12400 15550
rect 12640 15310 12730 15550
rect 12970 15310 13060 15550
rect 13300 15310 13390 15550
rect 13630 15310 13720 15550
rect 13960 15310 14050 15550
rect 14290 15310 14380 15550
rect 14620 15310 14710 15550
rect 14950 15310 15040 15550
rect 15280 15310 15370 15550
rect 15610 15310 15700 15550
rect 15940 15310 16030 15550
rect 16270 15310 16360 15550
rect 16600 15310 16690 15550
rect 16930 15310 17020 15550
rect 17260 15310 17350 15550
rect 17590 15310 17680 15550
rect 17920 15310 18010 15550
rect 18250 15310 18340 15550
rect 18580 15310 18670 15550
rect 18910 15310 19000 15550
rect 19240 15310 19330 15550
rect 19570 15310 19920 15550
rect 7610 15220 19920 15310
rect 7610 14980 7780 15220
rect 8020 14980 8110 15220
rect 8350 14980 8440 15220
rect 8680 14980 8770 15220
rect 9010 14980 9100 15220
rect 9340 14980 9430 15220
rect 9670 14980 9760 15220
rect 10000 14980 10090 15220
rect 10330 14980 10420 15220
rect 10660 14980 10750 15220
rect 10990 14980 11080 15220
rect 11320 14980 11410 15220
rect 11650 14980 11740 15220
rect 11980 14980 12070 15220
rect 12310 14980 12400 15220
rect 12640 14980 12730 15220
rect 12970 14980 13060 15220
rect 13300 14980 13390 15220
rect 13630 14980 13720 15220
rect 13960 14980 14050 15220
rect 14290 14980 14380 15220
rect 14620 14980 14710 15220
rect 14950 14980 15040 15220
rect 15280 14980 15370 15220
rect 15610 14980 15700 15220
rect 15940 14980 16030 15220
rect 16270 14980 16360 15220
rect 16600 14980 16690 15220
rect 16930 14980 17020 15220
rect 17260 14980 17350 15220
rect 17590 14980 17680 15220
rect 17920 14980 18010 15220
rect 18250 14980 18340 15220
rect 18580 14980 18670 15220
rect 18910 14980 19000 15220
rect 19240 14980 19330 15220
rect 19570 14980 19920 15220
rect 7610 14890 19920 14980
rect 7610 14650 7780 14890
rect 8020 14650 8110 14890
rect 8350 14650 8440 14890
rect 8680 14650 8770 14890
rect 9010 14650 9100 14890
rect 9340 14650 9430 14890
rect 9670 14650 9760 14890
rect 10000 14650 10090 14890
rect 10330 14650 10420 14890
rect 10660 14650 10750 14890
rect 10990 14650 11080 14890
rect 11320 14650 11410 14890
rect 11650 14650 11740 14890
rect 11980 14650 12070 14890
rect 12310 14650 12400 14890
rect 12640 14650 12730 14890
rect 12970 14650 13060 14890
rect 13300 14650 13390 14890
rect 13630 14650 13720 14890
rect 13960 14650 14050 14890
rect 14290 14650 14380 14890
rect 14620 14650 14710 14890
rect 14950 14650 15040 14890
rect 15280 14650 15370 14890
rect 15610 14650 15700 14890
rect 15940 14650 16030 14890
rect 16270 14650 16360 14890
rect 16600 14650 16690 14890
rect 16930 14650 17020 14890
rect 17260 14650 17350 14890
rect 17590 14650 17680 14890
rect 17920 14650 18010 14890
rect 18250 14650 18340 14890
rect 18580 14650 18670 14890
rect 18910 14650 19000 14890
rect 19240 14650 19330 14890
rect 19570 14650 19920 14890
rect 7610 14560 19920 14650
rect 7610 14320 7780 14560
rect 8020 14320 8110 14560
rect 8350 14320 8440 14560
rect 8680 14320 8770 14560
rect 9010 14320 9100 14560
rect 9340 14320 9430 14560
rect 9670 14320 9760 14560
rect 10000 14320 10090 14560
rect 10330 14320 10420 14560
rect 10660 14320 10750 14560
rect 10990 14320 11080 14560
rect 11320 14320 11410 14560
rect 11650 14320 11740 14560
rect 11980 14320 12070 14560
rect 12310 14320 12400 14560
rect 12640 14320 12730 14560
rect 12970 14320 13060 14560
rect 13300 14320 13390 14560
rect 13630 14320 13720 14560
rect 13960 14320 14050 14560
rect 14290 14320 14380 14560
rect 14620 14320 14710 14560
rect 14950 14320 15040 14560
rect 15280 14320 15370 14560
rect 15610 14320 15700 14560
rect 15940 14320 16030 14560
rect 16270 14320 16360 14560
rect 16600 14320 16690 14560
rect 16930 14320 17020 14560
rect 17260 14320 17350 14560
rect 17590 14320 17680 14560
rect 17920 14320 18010 14560
rect 18250 14320 18340 14560
rect 18580 14320 18670 14560
rect 18910 14320 19000 14560
rect 19240 14320 19330 14560
rect 19570 14320 19920 14560
rect 7610 14230 19920 14320
rect 7610 13990 7780 14230
rect 8020 13990 8110 14230
rect 8350 13990 8440 14230
rect 8680 13990 8770 14230
rect 9010 13990 9100 14230
rect 9340 13990 9430 14230
rect 9670 13990 9760 14230
rect 10000 13990 10090 14230
rect 10330 13990 10420 14230
rect 10660 13990 10750 14230
rect 10990 13990 11080 14230
rect 11320 13990 11410 14230
rect 11650 13990 11740 14230
rect 11980 13990 12070 14230
rect 12310 13990 12400 14230
rect 12640 13990 12730 14230
rect 12970 13990 13060 14230
rect 13300 13990 13390 14230
rect 13630 13990 13720 14230
rect 13960 13990 14050 14230
rect 14290 13990 14380 14230
rect 14620 13990 14710 14230
rect 14950 13990 15040 14230
rect 15280 13990 15370 14230
rect 15610 13990 15700 14230
rect 15940 13990 16030 14230
rect 16270 13990 16360 14230
rect 16600 13990 16690 14230
rect 16930 13990 17020 14230
rect 17260 13990 17350 14230
rect 17590 13990 17680 14230
rect 17920 13990 18010 14230
rect 18250 13990 18340 14230
rect 18580 13990 18670 14230
rect 18910 13990 19000 14230
rect 19240 13990 19330 14230
rect 19570 13990 19920 14230
rect 7610 13900 19920 13990
rect 7610 13660 7780 13900
rect 8020 13660 8110 13900
rect 8350 13660 8440 13900
rect 8680 13660 8770 13900
rect 9010 13660 9100 13900
rect 9340 13660 9430 13900
rect 9670 13660 9760 13900
rect 10000 13660 10090 13900
rect 10330 13660 10420 13900
rect 10660 13660 10750 13900
rect 10990 13660 11080 13900
rect 11320 13660 11410 13900
rect 11650 13660 11740 13900
rect 11980 13660 12070 13900
rect 12310 13660 12400 13900
rect 12640 13660 12730 13900
rect 12970 13660 13060 13900
rect 13300 13660 13390 13900
rect 13630 13660 13720 13900
rect 13960 13660 14050 13900
rect 14290 13660 14380 13900
rect 14620 13660 14710 13900
rect 14950 13660 15040 13900
rect 15280 13660 15370 13900
rect 15610 13660 15700 13900
rect 15940 13660 16030 13900
rect 16270 13660 16360 13900
rect 16600 13660 16690 13900
rect 16930 13660 17020 13900
rect 17260 13660 17350 13900
rect 17590 13660 17680 13900
rect 17920 13660 18010 13900
rect 18250 13660 18340 13900
rect 18580 13660 18670 13900
rect 18910 13660 19000 13900
rect 19240 13660 19330 13900
rect 19570 13660 19920 13900
rect 7610 13570 19920 13660
rect 7610 13330 7780 13570
rect 8020 13330 8110 13570
rect 8350 13330 8440 13570
rect 8680 13330 8770 13570
rect 9010 13330 9100 13570
rect 9340 13330 9430 13570
rect 9670 13330 9760 13570
rect 10000 13330 10090 13570
rect 10330 13330 10420 13570
rect 10660 13330 10750 13570
rect 10990 13330 11080 13570
rect 11320 13330 11410 13570
rect 11650 13330 11740 13570
rect 11980 13330 12070 13570
rect 12310 13330 12400 13570
rect 12640 13330 12730 13570
rect 12970 13330 13060 13570
rect 13300 13330 13390 13570
rect 13630 13330 13720 13570
rect 13960 13330 14050 13570
rect 14290 13330 14380 13570
rect 14620 13330 14710 13570
rect 14950 13330 15040 13570
rect 15280 13330 15370 13570
rect 15610 13330 15700 13570
rect 15940 13330 16030 13570
rect 16270 13330 16360 13570
rect 16600 13330 16690 13570
rect 16930 13330 17020 13570
rect 17260 13330 17350 13570
rect 17590 13330 17680 13570
rect 17920 13330 18010 13570
rect 18250 13330 18340 13570
rect 18580 13330 18670 13570
rect 18910 13330 19000 13570
rect 19240 13330 19330 13570
rect 19570 13330 19920 13570
rect 7610 13240 19920 13330
rect 7610 13000 7780 13240
rect 8020 13000 8110 13240
rect 8350 13000 8440 13240
rect 8680 13000 8770 13240
rect 9010 13000 9100 13240
rect 9340 13000 9430 13240
rect 9670 13000 9760 13240
rect 10000 13000 10090 13240
rect 10330 13000 10420 13240
rect 10660 13000 10750 13240
rect 10990 13000 11080 13240
rect 11320 13000 11410 13240
rect 11650 13000 11740 13240
rect 11980 13000 12070 13240
rect 12310 13000 12400 13240
rect 12640 13000 12730 13240
rect 12970 13000 13060 13240
rect 13300 13000 13390 13240
rect 13630 13000 13720 13240
rect 13960 13000 14050 13240
rect 14290 13000 14380 13240
rect 14620 13000 14710 13240
rect 14950 13000 15040 13240
rect 15280 13000 15370 13240
rect 15610 13000 15700 13240
rect 15940 13000 16030 13240
rect 16270 13000 16360 13240
rect 16600 13000 16690 13240
rect 16930 13000 17020 13240
rect 17260 13000 17350 13240
rect 17590 13000 17680 13240
rect 17920 13000 18010 13240
rect 18250 13000 18340 13240
rect 18580 13000 18670 13240
rect 18910 13000 19000 13240
rect 19240 13000 19330 13240
rect 19570 13000 19920 13240
rect 7610 12910 19920 13000
rect 7610 12670 7780 12910
rect 8020 12670 8110 12910
rect 8350 12670 8440 12910
rect 8680 12670 8770 12910
rect 9010 12670 9100 12910
rect 9340 12670 9430 12910
rect 9670 12670 9760 12910
rect 10000 12670 10090 12910
rect 10330 12670 10420 12910
rect 10660 12670 10750 12910
rect 10990 12670 11080 12910
rect 11320 12670 11410 12910
rect 11650 12670 11740 12910
rect 11980 12670 12070 12910
rect 12310 12670 12400 12910
rect 12640 12670 12730 12910
rect 12970 12670 13060 12910
rect 13300 12670 13390 12910
rect 13630 12670 13720 12910
rect 13960 12670 14050 12910
rect 14290 12670 14380 12910
rect 14620 12670 14710 12910
rect 14950 12670 15040 12910
rect 15280 12670 15370 12910
rect 15610 12670 15700 12910
rect 15940 12670 16030 12910
rect 16270 12670 16360 12910
rect 16600 12670 16690 12910
rect 16930 12670 17020 12910
rect 17260 12670 17350 12910
rect 17590 12670 17680 12910
rect 17920 12670 18010 12910
rect 18250 12670 18340 12910
rect 18580 12670 18670 12910
rect 18910 12670 19000 12910
rect 19240 12670 19330 12910
rect 19570 12670 19920 12910
rect 7610 12580 19920 12670
rect 7610 12340 7780 12580
rect 8020 12340 8110 12580
rect 8350 12340 8440 12580
rect 8680 12340 8770 12580
rect 9010 12340 9100 12580
rect 9340 12340 9430 12580
rect 9670 12340 9760 12580
rect 10000 12340 10090 12580
rect 10330 12340 10420 12580
rect 10660 12340 10750 12580
rect 10990 12340 11080 12580
rect 11320 12340 11410 12580
rect 11650 12340 11740 12580
rect 11980 12340 12070 12580
rect 12310 12340 12400 12580
rect 12640 12340 12730 12580
rect 12970 12340 13060 12580
rect 13300 12340 13390 12580
rect 13630 12340 13720 12580
rect 13960 12340 14050 12580
rect 14290 12340 14380 12580
rect 14620 12340 14710 12580
rect 14950 12340 15040 12580
rect 15280 12340 15370 12580
rect 15610 12340 15700 12580
rect 15940 12340 16030 12580
rect 16270 12340 16360 12580
rect 16600 12340 16690 12580
rect 16930 12340 17020 12580
rect 17260 12340 17350 12580
rect 17590 12340 17680 12580
rect 17920 12340 18010 12580
rect 18250 12340 18340 12580
rect 18580 12340 18670 12580
rect 18910 12340 19000 12580
rect 19240 12340 19330 12580
rect 19570 12340 19920 12580
rect 7610 12250 19920 12340
rect 7610 12010 7780 12250
rect 8020 12010 8110 12250
rect 8350 12010 8440 12250
rect 8680 12010 8770 12250
rect 9010 12010 9100 12250
rect 9340 12010 9430 12250
rect 9670 12010 9760 12250
rect 10000 12010 10090 12250
rect 10330 12010 10420 12250
rect 10660 12010 10750 12250
rect 10990 12010 11080 12250
rect 11320 12010 11410 12250
rect 11650 12010 11740 12250
rect 11980 12010 12070 12250
rect 12310 12010 12400 12250
rect 12640 12010 12730 12250
rect 12970 12010 13060 12250
rect 13300 12010 13390 12250
rect 13630 12010 13720 12250
rect 13960 12010 14050 12250
rect 14290 12010 14380 12250
rect 14620 12010 14710 12250
rect 14950 12010 15040 12250
rect 15280 12010 15370 12250
rect 15610 12010 15700 12250
rect 15940 12010 16030 12250
rect 16270 12010 16360 12250
rect 16600 12010 16690 12250
rect 16930 12010 17020 12250
rect 17260 12010 17350 12250
rect 17590 12010 17680 12250
rect 17920 12010 18010 12250
rect 18250 12010 18340 12250
rect 18580 12010 18670 12250
rect 18910 12010 19000 12250
rect 19240 12010 19330 12250
rect 19570 12010 19920 12250
rect 7610 11920 19920 12010
rect 7610 11680 7780 11920
rect 8020 11680 8110 11920
rect 8350 11680 8440 11920
rect 8680 11680 8770 11920
rect 9010 11680 9100 11920
rect 9340 11680 9430 11920
rect 9670 11680 9760 11920
rect 10000 11680 10090 11920
rect 10330 11680 10420 11920
rect 10660 11680 10750 11920
rect 10990 11680 11080 11920
rect 11320 11680 11410 11920
rect 11650 11680 11740 11920
rect 11980 11680 12070 11920
rect 12310 11680 12400 11920
rect 12640 11680 12730 11920
rect 12970 11680 13060 11920
rect 13300 11680 13390 11920
rect 13630 11680 13720 11920
rect 13960 11680 14050 11920
rect 14290 11680 14380 11920
rect 14620 11680 14710 11920
rect 14950 11680 15040 11920
rect 15280 11680 15370 11920
rect 15610 11680 15700 11920
rect 15940 11680 16030 11920
rect 16270 11680 16360 11920
rect 16600 11680 16690 11920
rect 16930 11680 17020 11920
rect 17260 11680 17350 11920
rect 17590 11680 17680 11920
rect 17920 11680 18010 11920
rect 18250 11680 18340 11920
rect 18580 11680 18670 11920
rect 18910 11680 19000 11920
rect 19240 11680 19330 11920
rect 19570 11680 19920 11920
rect 7610 11590 19920 11680
rect 7610 11350 7780 11590
rect 8020 11350 8110 11590
rect 8350 11350 8440 11590
rect 8680 11350 8770 11590
rect 9010 11350 9100 11590
rect 9340 11350 9430 11590
rect 9670 11350 9760 11590
rect 10000 11350 10090 11590
rect 10330 11350 10420 11590
rect 10660 11350 10750 11590
rect 10990 11350 11080 11590
rect 11320 11350 11410 11590
rect 11650 11350 11740 11590
rect 11980 11350 12070 11590
rect 12310 11350 12400 11590
rect 12640 11350 12730 11590
rect 12970 11350 13060 11590
rect 13300 11350 13390 11590
rect 13630 11350 13720 11590
rect 13960 11350 14050 11590
rect 14290 11350 14380 11590
rect 14620 11350 14710 11590
rect 14950 11350 15040 11590
rect 15280 11350 15370 11590
rect 15610 11350 15700 11590
rect 15940 11350 16030 11590
rect 16270 11350 16360 11590
rect 16600 11350 16690 11590
rect 16930 11350 17020 11590
rect 17260 11350 17350 11590
rect 17590 11350 17680 11590
rect 17920 11350 18010 11590
rect 18250 11350 18340 11590
rect 18580 11350 18670 11590
rect 18910 11350 19000 11590
rect 19240 11350 19330 11590
rect 19570 11350 19920 11590
rect 7610 11260 19920 11350
rect 7610 11020 7780 11260
rect 8020 11020 8110 11260
rect 8350 11020 8440 11260
rect 8680 11020 8770 11260
rect 9010 11020 9100 11260
rect 9340 11020 9430 11260
rect 9670 11020 9760 11260
rect 10000 11020 10090 11260
rect 10330 11020 10420 11260
rect 10660 11020 10750 11260
rect 10990 11020 11080 11260
rect 11320 11020 11410 11260
rect 11650 11020 11740 11260
rect 11980 11020 12070 11260
rect 12310 11020 12400 11260
rect 12640 11020 12730 11260
rect 12970 11020 13060 11260
rect 13300 11020 13390 11260
rect 13630 11020 13720 11260
rect 13960 11020 14050 11260
rect 14290 11020 14380 11260
rect 14620 11020 14710 11260
rect 14950 11020 15040 11260
rect 15280 11020 15370 11260
rect 15610 11020 15700 11260
rect 15940 11020 16030 11260
rect 16270 11020 16360 11260
rect 16600 11020 16690 11260
rect 16930 11020 17020 11260
rect 17260 11020 17350 11260
rect 17590 11020 17680 11260
rect 17920 11020 18010 11260
rect 18250 11020 18340 11260
rect 18580 11020 18670 11260
rect 18910 11020 19000 11260
rect 19240 11020 19330 11260
rect 19570 11020 19920 11260
rect 7610 10930 19920 11020
rect 7610 10690 7780 10930
rect 8020 10690 8110 10930
rect 8350 10690 8440 10930
rect 8680 10690 8770 10930
rect 9010 10690 9100 10930
rect 9340 10690 9430 10930
rect 9670 10690 9760 10930
rect 10000 10690 10090 10930
rect 10330 10690 10420 10930
rect 10660 10690 10750 10930
rect 10990 10690 11080 10930
rect 11320 10690 11410 10930
rect 11650 10690 11740 10930
rect 11980 10690 12070 10930
rect 12310 10690 12400 10930
rect 12640 10690 12730 10930
rect 12970 10690 13060 10930
rect 13300 10690 13390 10930
rect 13630 10690 13720 10930
rect 13960 10690 14050 10930
rect 14290 10690 14380 10930
rect 14620 10690 14710 10930
rect 14950 10690 15040 10930
rect 15280 10690 15370 10930
rect 15610 10690 15700 10930
rect 15940 10690 16030 10930
rect 16270 10690 16360 10930
rect 16600 10690 16690 10930
rect 16930 10690 17020 10930
rect 17260 10690 17350 10930
rect 17590 10690 17680 10930
rect 17920 10690 18010 10930
rect 18250 10690 18340 10930
rect 18580 10690 18670 10930
rect 18910 10690 19000 10930
rect 19240 10690 19330 10930
rect 19570 10690 19920 10930
rect 7610 10600 19920 10690
rect 7610 10360 7780 10600
rect 8020 10360 8110 10600
rect 8350 10360 8440 10600
rect 8680 10360 8770 10600
rect 9010 10360 9100 10600
rect 9340 10360 9430 10600
rect 9670 10360 9760 10600
rect 10000 10360 10090 10600
rect 10330 10360 10420 10600
rect 10660 10360 10750 10600
rect 10990 10360 11080 10600
rect 11320 10360 11410 10600
rect 11650 10360 11740 10600
rect 11980 10360 12070 10600
rect 12310 10360 12400 10600
rect 12640 10360 12730 10600
rect 12970 10360 13060 10600
rect 13300 10360 13390 10600
rect 13630 10360 13720 10600
rect 13960 10360 14050 10600
rect 14290 10360 14380 10600
rect 14620 10360 14710 10600
rect 14950 10360 15040 10600
rect 15280 10360 15370 10600
rect 15610 10360 15700 10600
rect 15940 10360 16030 10600
rect 16270 10360 16360 10600
rect 16600 10360 16690 10600
rect 16930 10360 17020 10600
rect 17260 10360 17350 10600
rect 17590 10360 17680 10600
rect 17920 10360 18010 10600
rect 18250 10360 18340 10600
rect 18580 10360 18670 10600
rect 18910 10360 19000 10600
rect 19240 10360 19330 10600
rect 19570 10360 19920 10600
rect 7610 10270 19920 10360
rect 7610 10030 7780 10270
rect 8020 10030 8110 10270
rect 8350 10030 8440 10270
rect 8680 10030 8770 10270
rect 9010 10030 9100 10270
rect 9340 10030 9430 10270
rect 9670 10030 9760 10270
rect 10000 10030 10090 10270
rect 10330 10030 10420 10270
rect 10660 10030 10750 10270
rect 10990 10030 11080 10270
rect 11320 10030 11410 10270
rect 11650 10030 11740 10270
rect 11980 10030 12070 10270
rect 12310 10030 12400 10270
rect 12640 10030 12730 10270
rect 12970 10030 13060 10270
rect 13300 10030 13390 10270
rect 13630 10030 13720 10270
rect 13960 10030 14050 10270
rect 14290 10030 14380 10270
rect 14620 10030 14710 10270
rect 14950 10030 15040 10270
rect 15280 10030 15370 10270
rect 15610 10030 15700 10270
rect 15940 10030 16030 10270
rect 16270 10030 16360 10270
rect 16600 10030 16690 10270
rect 16930 10030 17020 10270
rect 17260 10030 17350 10270
rect 17590 10030 17680 10270
rect 17920 10030 18010 10270
rect 18250 10030 18340 10270
rect 18580 10030 18670 10270
rect 18910 10030 19000 10270
rect 19240 10030 19330 10270
rect 19570 10030 19920 10270
rect 7610 9940 19920 10030
rect 7610 9700 7780 9940
rect 8020 9700 8110 9940
rect 8350 9700 8440 9940
rect 8680 9700 8770 9940
rect 9010 9700 9100 9940
rect 9340 9700 9430 9940
rect 9670 9700 9760 9940
rect 10000 9700 10090 9940
rect 10330 9700 10420 9940
rect 10660 9700 10750 9940
rect 10990 9700 11080 9940
rect 11320 9700 11410 9940
rect 11650 9700 11740 9940
rect 11980 9700 12070 9940
rect 12310 9700 12400 9940
rect 12640 9700 12730 9940
rect 12970 9700 13060 9940
rect 13300 9700 13390 9940
rect 13630 9700 13720 9940
rect 13960 9700 14050 9940
rect 14290 9700 14380 9940
rect 14620 9700 14710 9940
rect 14950 9700 15040 9940
rect 15280 9700 15370 9940
rect 15610 9700 15700 9940
rect 15940 9700 16030 9940
rect 16270 9700 16360 9940
rect 16600 9700 16690 9940
rect 16930 9700 17020 9940
rect 17260 9700 17350 9940
rect 17590 9700 17680 9940
rect 17920 9700 18010 9940
rect 18250 9700 18340 9940
rect 18580 9700 18670 9940
rect 18910 9700 19000 9940
rect 19240 9700 19330 9940
rect 19570 9700 19920 9940
rect 7610 9610 19920 9700
rect 7610 9370 7780 9610
rect 8020 9370 8110 9610
rect 8350 9370 8440 9610
rect 8680 9370 8770 9610
rect 9010 9370 9100 9610
rect 9340 9370 9430 9610
rect 9670 9370 9760 9610
rect 10000 9370 10090 9610
rect 10330 9370 10420 9610
rect 10660 9370 10750 9610
rect 10990 9370 11080 9610
rect 11320 9370 11410 9610
rect 11650 9370 11740 9610
rect 11980 9370 12070 9610
rect 12310 9370 12400 9610
rect 12640 9370 12730 9610
rect 12970 9370 13060 9610
rect 13300 9370 13390 9610
rect 13630 9370 13720 9610
rect 13960 9370 14050 9610
rect 14290 9370 14380 9610
rect 14620 9370 14710 9610
rect 14950 9370 15040 9610
rect 15280 9370 15370 9610
rect 15610 9370 15700 9610
rect 15940 9370 16030 9610
rect 16270 9370 16360 9610
rect 16600 9370 16690 9610
rect 16930 9370 17020 9610
rect 17260 9370 17350 9610
rect 17590 9370 17680 9610
rect 17920 9370 18010 9610
rect 18250 9370 18340 9610
rect 18580 9370 18670 9610
rect 18910 9370 19000 9610
rect 19240 9370 19330 9610
rect 19570 9370 19920 9610
rect 7610 9280 19920 9370
rect 7610 9040 7780 9280
rect 8020 9040 8110 9280
rect 8350 9040 8440 9280
rect 8680 9040 8770 9280
rect 9010 9040 9100 9280
rect 9340 9040 9430 9280
rect 9670 9040 9760 9280
rect 10000 9040 10090 9280
rect 10330 9040 10420 9280
rect 10660 9040 10750 9280
rect 10990 9040 11080 9280
rect 11320 9040 11410 9280
rect 11650 9040 11740 9280
rect 11980 9040 12070 9280
rect 12310 9040 12400 9280
rect 12640 9040 12730 9280
rect 12970 9040 13060 9280
rect 13300 9040 13390 9280
rect 13630 9040 13720 9280
rect 13960 9040 14050 9280
rect 14290 9040 14380 9280
rect 14620 9040 14710 9280
rect 14950 9040 15040 9280
rect 15280 9040 15370 9280
rect 15610 9040 15700 9280
rect 15940 9040 16030 9280
rect 16270 9040 16360 9280
rect 16600 9040 16690 9280
rect 16930 9040 17020 9280
rect 17260 9040 17350 9280
rect 17590 9040 17680 9280
rect 17920 9040 18010 9280
rect 18250 9040 18340 9280
rect 18580 9040 18670 9280
rect 18910 9040 19000 9280
rect 19240 9040 19330 9280
rect 19570 9040 19920 9280
rect 7610 8690 19920 9040
rect 7610 8410 7880 8690
rect 7610 8340 7630 8410
rect 7730 8340 7760 8410
rect 7860 8340 7880 8410
rect 7610 8320 7880 8340
rect 7610 8250 7630 8320
rect 7730 8250 7760 8320
rect 7860 8250 7880 8320
rect 7610 8230 7880 8250
rect 11760 6940 13360 6960
rect 1540 6910 3140 6930
rect 1540 6850 1720 6910
rect 1960 6850 2050 6910
rect 2290 6850 2390 6910
rect 2630 6850 2720 6910
rect 2960 6850 3140 6910
rect 1540 6780 1570 6850
rect 1640 6780 1680 6850
rect 1970 6780 2010 6850
rect 2300 6780 2340 6850
rect 2630 6780 2670 6850
rect 2960 6780 3000 6850
rect 3070 6780 3140 6850
rect 1540 6740 1720 6780
rect 1960 6740 2050 6780
rect 2290 6740 2390 6780
rect 2630 6740 2720 6780
rect 2960 6740 3140 6780
rect 1540 6670 1570 6740
rect 1640 6670 1680 6740
rect 1970 6670 2010 6740
rect 2300 6670 2340 6740
rect 2630 6670 2670 6740
rect 2960 6670 3000 6740
rect 3070 6670 3140 6740
rect 11760 6880 11940 6940
rect 12180 6880 12270 6940
rect 12510 6880 12610 6940
rect 12850 6880 12940 6940
rect 13180 6880 13360 6940
rect 11760 6810 11790 6880
rect 11860 6810 11900 6880
rect 12190 6810 12230 6880
rect 12520 6810 12560 6880
rect 12850 6810 12890 6880
rect 13180 6810 13220 6880
rect 13290 6810 13360 6880
rect 11760 6770 11940 6810
rect 12180 6770 12270 6810
rect 12510 6770 12610 6810
rect 12850 6770 12940 6810
rect 13180 6770 13360 6810
rect 11760 6700 11790 6770
rect 11860 6700 11900 6770
rect 12190 6700 12230 6770
rect 12520 6700 12560 6770
rect 12850 6700 12890 6770
rect 13180 6700 13220 6770
rect 13290 6700 13360 6770
rect 11760 6670 13360 6700
rect 1540 6640 3140 6670
rect 7400 5390 7490 5410
rect 7400 5320 7410 5390
rect 7480 5320 7490 5390
rect 7400 5280 7490 5320
rect 7400 5210 7410 5280
rect 7480 5240 7490 5280
rect 21120 5240 21280 8880
rect 7480 5210 21280 5240
rect 7400 5170 21280 5210
rect 7400 5100 7410 5170
rect 7480 5100 21280 5170
rect 7400 5080 21280 5100
rect 21800 8230 39650 8490
rect 21800 5670 22060 8230
rect 31100 7830 37860 7910
rect 31100 7590 31180 7830
rect 31420 7590 31510 7830
rect 31750 7590 31840 7830
rect 32080 7590 32170 7830
rect 32410 7590 32500 7830
rect 32740 7590 32830 7830
rect 33070 7590 33160 7830
rect 33400 7590 33490 7830
rect 33730 7590 33820 7830
rect 34060 7590 34150 7830
rect 34390 7590 34480 7830
rect 34720 7590 34810 7830
rect 35050 7590 35140 7830
rect 35380 7590 35470 7830
rect 35710 7590 35800 7830
rect 36040 7590 36130 7830
rect 36370 7590 36460 7830
rect 36700 7590 36790 7830
rect 37030 7590 37120 7830
rect 37360 7590 37450 7830
rect 37690 7590 37860 7830
rect 31100 7500 37860 7590
rect 23460 7270 23940 7290
rect 23460 7210 23510 7270
rect 23880 7210 23940 7270
rect 23460 7140 23490 7210
rect 23890 7140 23940 7210
rect 23460 7100 23510 7140
rect 23880 7100 23940 7140
rect 23460 7030 23490 7100
rect 23890 7030 23940 7100
rect 23460 7000 23940 7030
rect 25860 7270 26340 7290
rect 25860 7210 25910 7270
rect 26280 7210 26340 7270
rect 25860 7140 25890 7210
rect 26290 7140 26340 7210
rect 25860 7100 25910 7140
rect 26280 7100 26340 7140
rect 25860 7030 25890 7100
rect 26290 7030 26340 7100
rect 25860 7000 26340 7030
rect 31100 7260 31180 7500
rect 31420 7260 31510 7500
rect 31750 7260 31840 7500
rect 32080 7260 32170 7500
rect 32410 7260 32500 7500
rect 32740 7260 32830 7500
rect 33070 7260 33160 7500
rect 33400 7260 33490 7500
rect 33730 7260 33820 7500
rect 34060 7260 34150 7500
rect 34390 7260 34480 7500
rect 34720 7260 34810 7500
rect 35050 7260 35140 7500
rect 35380 7260 35470 7500
rect 35710 7260 35800 7500
rect 36040 7260 36130 7500
rect 36370 7260 36460 7500
rect 36700 7260 36790 7500
rect 37030 7260 37120 7500
rect 37360 7260 37450 7500
rect 37690 7260 37860 7500
rect 31100 7170 37860 7260
rect 31100 6930 31180 7170
rect 31420 6930 31510 7170
rect 31750 6930 31840 7170
rect 32080 6930 32170 7170
rect 32410 6930 32500 7170
rect 32740 6930 32830 7170
rect 33070 6930 33160 7170
rect 33400 6930 33490 7170
rect 33730 6930 33820 7170
rect 34060 6930 34150 7170
rect 34390 6930 34480 7170
rect 34720 6930 34810 7170
rect 35050 6930 35140 7170
rect 35380 6930 35470 7170
rect 35710 6930 35800 7170
rect 36040 6930 36130 7170
rect 36370 6930 36460 7170
rect 36700 6930 36790 7170
rect 37030 6930 37120 7170
rect 37360 6930 37450 7170
rect 37690 6930 37860 7170
rect 31100 6840 37860 6930
rect 31100 6600 31180 6840
rect 31420 6600 31510 6840
rect 31750 6600 31840 6840
rect 32080 6600 32170 6840
rect 32410 6600 32500 6840
rect 32740 6600 32830 6840
rect 33070 6600 33160 6840
rect 33400 6600 33490 6840
rect 33730 6600 33820 6840
rect 34060 6600 34150 6840
rect 34390 6600 34480 6840
rect 34720 6600 34810 6840
rect 35050 6600 35140 6840
rect 35380 6600 35470 6840
rect 35710 6600 35800 6840
rect 36040 6600 36130 6840
rect 36370 6600 36460 6840
rect 36700 6600 36790 6840
rect 37030 6600 37120 6840
rect 37360 6600 37450 6840
rect 37690 6600 37860 6840
rect 31100 6510 37860 6600
rect 31100 6320 31180 6510
rect 30720 6300 31180 6320
rect 30720 6230 30740 6300
rect 30810 6230 30850 6300
rect 30920 6270 31180 6300
rect 31420 6270 31510 6510
rect 31750 6270 31840 6510
rect 32080 6270 32170 6510
rect 32410 6270 32500 6510
rect 32740 6270 32830 6510
rect 33070 6270 33160 6510
rect 33400 6270 33490 6510
rect 33730 6270 33820 6510
rect 34060 6270 34150 6510
rect 34390 6270 34480 6510
rect 34720 6270 34810 6510
rect 35050 6270 35140 6510
rect 35380 6270 35470 6510
rect 35710 6270 35800 6510
rect 36040 6270 36130 6510
rect 36370 6270 36460 6510
rect 36700 6270 36790 6510
rect 37030 6270 37120 6510
rect 37360 6270 37450 6510
rect 37690 6270 37860 6510
rect 30920 6230 37860 6270
rect 30720 6180 37860 6230
rect 30720 6170 31180 6180
rect 30720 6100 30740 6170
rect 30810 6100 30850 6170
rect 30920 6100 31180 6170
rect 30720 6040 31180 6100
rect 30720 5970 30740 6040
rect 30810 5970 30850 6040
rect 30920 5970 31180 6040
rect 30720 5950 31180 5970
rect 21800 5600 21820 5670
rect 21890 5600 21930 5670
rect 22000 5600 22060 5670
rect 21800 5560 22060 5600
rect 21800 5490 21820 5560
rect 21890 5490 21930 5560
rect 22000 5490 22060 5560
rect 21800 5450 22060 5490
rect 21800 5380 21820 5450
rect 21890 5380 21930 5450
rect 22000 5380 22060 5450
rect 21800 5340 22060 5380
rect 21800 5270 21820 5340
rect 21890 5270 21930 5340
rect 22000 5270 22060 5340
rect 21800 5230 22060 5270
rect 21800 5160 21820 5230
rect 21890 5160 21930 5230
rect 22000 5160 22060 5230
rect 21800 5120 22060 5160
rect 7400 5060 7490 5080
rect 7400 4990 7410 5060
rect 7480 4990 7490 5060
rect 7400 4950 7490 4990
rect 7400 4880 7410 4950
rect 7480 4880 7490 4950
rect 7400 4860 7490 4880
rect 1080 -790 2680 -760
rect 1080 -860 1150 -790
rect 1220 -860 1260 -790
rect 1550 -860 1590 -790
rect 1880 -860 1920 -790
rect 2210 -860 2250 -790
rect 2540 -860 2580 -790
rect 2650 -860 2680 -790
rect 1080 -900 1260 -860
rect 1500 -900 1590 -860
rect 1830 -900 1930 -860
rect 2170 -900 2260 -860
rect 2500 -900 2680 -860
rect 1080 -970 1150 -900
rect 1220 -970 1260 -900
rect 1550 -970 1590 -900
rect 1880 -970 1920 -900
rect 2210 -970 2250 -900
rect 2540 -970 2580 -900
rect 2650 -970 2680 -900
rect 1080 -1030 1260 -970
rect 1500 -1030 1590 -970
rect 1830 -1030 1930 -970
rect 2170 -1030 2260 -970
rect 2500 -1030 2680 -970
rect 1080 -1050 2680 -1030
rect 12220 -790 13820 -760
rect 12220 -860 12250 -790
rect 12320 -860 12360 -790
rect 12650 -860 12690 -790
rect 12980 -860 13020 -790
rect 13310 -860 13350 -790
rect 13640 -860 13680 -790
rect 13750 -860 13820 -790
rect 12220 -900 12400 -860
rect 12640 -900 12730 -860
rect 12970 -900 13070 -860
rect 13310 -900 13400 -860
rect 13640 -900 13820 -860
rect 12220 -970 12250 -900
rect 12320 -970 12360 -900
rect 12650 -970 12690 -900
rect 12980 -970 13020 -900
rect 13310 -970 13350 -900
rect 13640 -970 13680 -900
rect 13750 -970 13820 -900
rect 12220 -1030 12400 -970
rect 12640 -1030 12730 -970
rect 12970 -1030 13070 -970
rect 13310 -1030 13400 -970
rect 13640 -1030 13820 -970
rect 12220 -1050 13820 -1030
rect 1540 -2720 3140 -2700
rect 1540 -2780 1720 -2720
rect 1960 -2780 2050 -2720
rect 2290 -2780 2390 -2720
rect 2630 -2780 2720 -2720
rect 2960 -2780 3140 -2720
rect 1540 -2850 1570 -2780
rect 1640 -2850 1680 -2780
rect 1970 -2850 2010 -2780
rect 2300 -2850 2340 -2780
rect 2630 -2850 2670 -2780
rect 2960 -2850 3000 -2780
rect 3070 -2850 3140 -2780
rect 1540 -2890 1720 -2850
rect 1960 -2890 2050 -2850
rect 2290 -2890 2390 -2850
rect 2630 -2890 2720 -2850
rect 2960 -2890 3140 -2850
rect 1540 -2960 1570 -2890
rect 1640 -2960 1680 -2890
rect 1970 -2960 2010 -2890
rect 2300 -2960 2340 -2890
rect 2630 -2960 2670 -2890
rect 2960 -2960 3000 -2890
rect 3070 -2960 3140 -2890
rect 1540 -2990 3140 -2960
rect 11760 -2720 13360 -2700
rect 11760 -2780 11940 -2720
rect 12180 -2780 12270 -2720
rect 12510 -2780 12610 -2720
rect 12850 -2780 12940 -2720
rect 13180 -2780 13360 -2720
rect 11760 -2850 11790 -2780
rect 11860 -2850 11900 -2780
rect 12190 -2850 12230 -2780
rect 12520 -2850 12560 -2780
rect 12850 -2850 12890 -2780
rect 13180 -2850 13220 -2780
rect 13290 -2850 13360 -2780
rect 11760 -2890 11940 -2850
rect 12180 -2890 12270 -2850
rect 12510 -2890 12610 -2850
rect 12850 -2890 12940 -2850
rect 13180 -2890 13360 -2850
rect 11760 -2960 11790 -2890
rect 11860 -2960 11900 -2890
rect 12190 -2960 12230 -2890
rect 12520 -2960 12560 -2890
rect 12850 -2960 12890 -2890
rect 13180 -2960 13220 -2890
rect 13290 -2960 13360 -2890
rect 11760 -2990 13360 -2960
rect 7290 -3880 7620 -3860
rect 7290 -3950 7310 -3880
rect 7380 -3950 7420 -3880
rect 7490 -3950 7530 -3880
rect 7600 -3920 7620 -3880
rect 17190 -3920 17350 5080
rect 21800 5050 21820 5120
rect 21890 5050 21930 5120
rect 22000 5050 22060 5120
rect 21800 5010 22060 5050
rect 21800 4940 21820 5010
rect 21890 4940 21930 5010
rect 22000 4940 22060 5010
rect 21800 4900 22060 4940
rect 21800 4830 21820 4900
rect 21890 4830 21930 4900
rect 22000 4830 22060 4900
rect 21800 4790 22060 4830
rect 21800 4720 21820 4790
rect 21890 4720 21930 4790
rect 22000 4720 22060 4790
rect 21800 4680 22060 4720
rect 21800 4610 21820 4680
rect 21890 4610 21930 4680
rect 22000 4610 22060 4680
rect 21800 4570 22060 4610
rect 21800 4500 21820 4570
rect 21890 4500 21930 4570
rect 22000 4500 22060 4570
rect 17450 1160 17580 1180
rect 17450 1090 17480 1160
rect 17550 1090 17580 1160
rect 17450 1050 19085 1090
rect 17450 980 17480 1050
rect 17550 980 19085 1050
rect 17450 960 19085 980
rect 17450 940 17580 960
rect 17450 870 17480 940
rect 17550 870 17580 940
rect 17450 850 17580 870
rect 7600 -3950 17350 -3920
rect 7290 -3990 17350 -3950
rect 7290 -4060 7310 -3990
rect 7380 -4060 7420 -3990
rect 7490 -4060 7530 -3990
rect 7600 -4060 17350 -3990
rect 7290 -4080 17350 -4060
rect 7290 -4100 7620 -4080
rect 7290 -4170 7310 -4100
rect 7380 -4170 7420 -4100
rect 7490 -4170 7530 -4100
rect 7600 -4170 7620 -4100
rect 7290 -4190 7620 -4170
rect -1350 -4350 -870 -4270
rect -1350 -4420 -1330 -4350
rect -1260 -4420 -1220 -4350
rect -1150 -4420 -1110 -4350
rect -1040 -4420 -1000 -4350
rect -930 -4420 -870 -4350
rect -1350 -4460 -870 -4420
rect -1350 -4530 -1330 -4460
rect -1260 -4530 -1220 -4460
rect -1150 -4530 -1110 -4460
rect -1040 -4530 -1000 -4460
rect -930 -4530 -870 -4460
rect -1350 -4630 -870 -4530
rect 15650 -4350 16130 -4270
rect 15650 -4420 15710 -4350
rect 15780 -4420 15820 -4350
rect 15890 -4420 15930 -4350
rect 16000 -4420 16040 -4350
rect 16110 -4420 16130 -4350
rect 15650 -4460 16130 -4420
rect 15650 -4530 15710 -4460
rect 15780 -4530 15820 -4460
rect 15890 -4530 15930 -4460
rect 16000 -4530 16040 -4460
rect 16110 -4530 16130 -4460
rect 15650 -4630 16130 -4530
rect -1350 -4840 260 -4630
rect -1350 -5080 -1180 -4840
rect -940 -5080 -850 -4840
rect -610 -5080 -520 -4840
rect -280 -5080 -190 -4840
rect 50 -5080 260 -4840
rect -1350 -5170 260 -5080
rect -1350 -5410 -1180 -5170
rect -940 -5410 -850 -5170
rect -610 -5410 -520 -5170
rect -280 -5410 -190 -5170
rect 50 -5410 260 -5170
rect -1350 -5500 260 -5410
rect -1350 -5740 -1180 -5500
rect -940 -5740 -850 -5500
rect -610 -5740 -520 -5500
rect -280 -5740 -190 -5500
rect 50 -5740 260 -5500
rect -1350 -5830 260 -5740
rect -1350 -6070 -1180 -5830
rect -940 -6070 -850 -5830
rect -610 -6070 -520 -5830
rect -280 -6070 -190 -5830
rect 50 -6070 260 -5830
rect -1350 -6240 260 -6070
rect 14520 -4840 16130 -4630
rect 14520 -5080 14730 -4840
rect 14970 -5080 15060 -4840
rect 15300 -5080 15390 -4840
rect 15630 -5080 15720 -4840
rect 15960 -5080 16130 -4840
rect 14520 -5170 16130 -5080
rect 14520 -5410 14730 -5170
rect 14970 -5410 15060 -5170
rect 15300 -5410 15390 -5170
rect 15630 -5410 15720 -5170
rect 15960 -5410 16130 -5170
rect 14520 -5500 16130 -5410
rect 14520 -5740 14730 -5500
rect 14970 -5740 15060 -5500
rect 15300 -5740 15390 -5500
rect 15630 -5740 15720 -5500
rect 15960 -5740 16130 -5500
rect 14520 -5830 16130 -5740
rect 14520 -6070 14730 -5830
rect 14970 -6070 15060 -5830
rect 15300 -6070 15390 -5830
rect 15630 -6070 15720 -5830
rect 15960 -6070 16130 -5830
rect 14520 -6240 16130 -6070
rect 18975 -5915 19085 960
rect 21800 -850 22060 4500
rect 31100 5940 31180 5950
rect 31420 5940 31510 6180
rect 31750 5940 31840 6180
rect 32080 5940 32170 6180
rect 32410 5940 32500 6180
rect 32740 5940 32830 6180
rect 33070 5940 33160 6180
rect 33400 5940 33490 6180
rect 33730 5940 33820 6180
rect 34060 5940 34150 6180
rect 34390 5940 34480 6180
rect 34720 5940 34810 6180
rect 35050 5940 35140 6180
rect 35380 5940 35470 6180
rect 35710 5940 35800 6180
rect 36040 5940 36130 6180
rect 36370 5940 36460 6180
rect 36700 5940 36790 6180
rect 37030 5940 37120 6180
rect 37360 5940 37450 6180
rect 37690 5940 37860 6180
rect 31100 5850 37860 5940
rect 31100 5610 31180 5850
rect 31420 5610 31510 5850
rect 31750 5610 31840 5850
rect 32080 5610 32170 5850
rect 32410 5610 32500 5850
rect 32740 5610 32830 5850
rect 33070 5610 33160 5850
rect 33400 5610 33490 5850
rect 33730 5610 33820 5850
rect 34060 5610 34150 5850
rect 34390 5610 34480 5850
rect 34720 5610 34810 5850
rect 35050 5610 35140 5850
rect 35380 5610 35470 5850
rect 35710 5610 35800 5850
rect 36040 5610 36130 5850
rect 36370 5610 36460 5850
rect 36700 5610 36790 5850
rect 37030 5610 37120 5850
rect 37360 5610 37450 5850
rect 37690 5610 37860 5850
rect 31100 5520 37860 5610
rect 31100 5280 31180 5520
rect 31420 5280 31510 5520
rect 31750 5280 31840 5520
rect 32080 5280 32170 5520
rect 32410 5280 32500 5520
rect 32740 5280 32830 5520
rect 33070 5280 33160 5520
rect 33400 5280 33490 5520
rect 33730 5280 33820 5520
rect 34060 5280 34150 5520
rect 34390 5280 34480 5520
rect 34720 5280 34810 5520
rect 35050 5280 35140 5520
rect 35380 5280 35470 5520
rect 35710 5280 35800 5520
rect 36040 5280 36130 5520
rect 36370 5280 36460 5520
rect 36700 5280 36790 5520
rect 37030 5280 37120 5520
rect 37360 5280 37450 5520
rect 37690 5280 37860 5520
rect 31100 5190 37860 5280
rect 31100 4950 31180 5190
rect 31420 4950 31510 5190
rect 31750 4950 31840 5190
rect 32080 4950 32170 5190
rect 32410 4950 32500 5190
rect 32740 4950 32830 5190
rect 33070 4950 33160 5190
rect 33400 4950 33490 5190
rect 33730 4950 33820 5190
rect 34060 4950 34150 5190
rect 34390 4950 34480 5190
rect 34720 4950 34810 5190
rect 35050 4950 35140 5190
rect 35380 4950 35470 5190
rect 35710 4950 35800 5190
rect 36040 4950 36130 5190
rect 36370 4950 36460 5190
rect 36700 4950 36790 5190
rect 37030 4950 37120 5190
rect 37360 4950 37450 5190
rect 37690 4950 37860 5190
rect 31100 4860 37860 4950
rect 31100 4620 31180 4860
rect 31420 4620 31510 4860
rect 31750 4620 31840 4860
rect 32080 4620 32170 4860
rect 32410 4620 32500 4860
rect 32740 4620 32830 4860
rect 33070 4620 33160 4860
rect 33400 4620 33490 4860
rect 33730 4620 33820 4860
rect 34060 4620 34150 4860
rect 34390 4620 34480 4860
rect 34720 4620 34810 4860
rect 35050 4620 35140 4860
rect 35380 4620 35470 4860
rect 35710 4620 35800 4860
rect 36040 4620 36130 4860
rect 36370 4620 36460 4860
rect 36700 4620 36790 4860
rect 37030 4620 37120 4860
rect 37360 4620 37450 4860
rect 37690 4620 37860 4860
rect 31100 4530 37860 4620
rect 31100 4290 31180 4530
rect 31420 4290 31510 4530
rect 31750 4290 31840 4530
rect 32080 4290 32170 4530
rect 32410 4290 32500 4530
rect 32740 4290 32830 4530
rect 33070 4290 33160 4530
rect 33400 4290 33490 4530
rect 33730 4290 33820 4530
rect 34060 4290 34150 4530
rect 34390 4290 34480 4530
rect 34720 4290 34810 4530
rect 35050 4290 35140 4530
rect 35380 4290 35470 4530
rect 35710 4290 35800 4530
rect 36040 4290 36130 4530
rect 36370 4290 36460 4530
rect 36700 4290 36790 4530
rect 37030 4290 37120 4530
rect 37360 4290 37450 4530
rect 37690 4290 37860 4530
rect 31100 4200 37860 4290
rect 31100 3960 31180 4200
rect 31420 3960 31510 4200
rect 31750 3960 31840 4200
rect 32080 3960 32170 4200
rect 32410 3960 32500 4200
rect 32740 3960 32830 4200
rect 33070 3960 33160 4200
rect 33400 3960 33490 4200
rect 33730 3960 33820 4200
rect 34060 3960 34150 4200
rect 34390 3960 34480 4200
rect 34720 3960 34810 4200
rect 35050 3960 35140 4200
rect 35380 3960 35470 4200
rect 35710 3960 35800 4200
rect 36040 3960 36130 4200
rect 36370 3960 36460 4200
rect 36700 3960 36790 4200
rect 37030 3960 37120 4200
rect 37360 3960 37450 4200
rect 37690 3960 37860 4200
rect 31100 3870 37860 3960
rect 31100 3630 31180 3870
rect 31420 3630 31510 3870
rect 31750 3630 31840 3870
rect 32080 3630 32170 3870
rect 32410 3630 32500 3870
rect 32740 3630 32830 3870
rect 33070 3630 33160 3870
rect 33400 3630 33490 3870
rect 33730 3630 33820 3870
rect 34060 3630 34150 3870
rect 34390 3630 34480 3870
rect 34720 3630 34810 3870
rect 35050 3630 35140 3870
rect 35380 3630 35470 3870
rect 35710 3630 35800 3870
rect 36040 3630 36130 3870
rect 36370 3630 36460 3870
rect 36700 3630 36790 3870
rect 37030 3630 37120 3870
rect 37360 3630 37450 3870
rect 37690 3630 37860 3870
rect 31100 3540 37860 3630
rect 24700 3360 25030 3380
rect 24700 3290 24720 3360
rect 24790 3290 24830 3360
rect 24900 3290 24940 3360
rect 25010 3290 25030 3360
rect 24700 3250 25030 3290
rect 24700 3236 24720 3250
rect 24684 3180 24720 3236
rect 24790 3180 24830 3250
rect 24900 3180 24940 3250
rect 25010 3236 25030 3250
rect 31100 3300 31180 3540
rect 31420 3300 31510 3540
rect 31750 3300 31840 3540
rect 32080 3300 32170 3540
rect 32410 3300 32500 3540
rect 32740 3300 32830 3540
rect 33070 3300 33160 3540
rect 33400 3300 33490 3540
rect 33730 3300 33820 3540
rect 34060 3300 34150 3540
rect 34390 3300 34480 3540
rect 34720 3300 34810 3540
rect 35050 3300 35140 3540
rect 35380 3300 35470 3540
rect 35710 3300 35800 3540
rect 36040 3300 36130 3540
rect 36370 3300 36460 3540
rect 36700 3300 36790 3540
rect 37030 3300 37120 3540
rect 37360 3300 37450 3540
rect 37690 3300 37860 3540
rect 25010 3180 30477 3236
rect 24684 3140 30477 3180
rect 24684 3103 24720 3140
rect 24700 3070 24720 3103
rect 24790 3070 24830 3140
rect 24900 3070 24940 3140
rect 25010 3103 30477 3140
rect 25010 3070 25030 3103
rect 24700 3050 25030 3070
rect 22420 2600 22900 2630
rect 22420 2530 22470 2600
rect 22870 2530 22900 2600
rect 22420 2490 22480 2530
rect 22850 2490 22900 2530
rect 22420 2420 22470 2490
rect 22870 2420 22900 2490
rect 22420 2360 22480 2420
rect 22850 2360 22900 2420
rect 22420 2340 22900 2360
rect 26900 2600 27380 2630
rect 26900 2530 26950 2600
rect 27350 2530 27380 2600
rect 26900 2490 26960 2530
rect 27330 2490 27380 2530
rect 26900 2420 26950 2490
rect 27350 2420 27380 2490
rect 26900 2360 26960 2420
rect 27330 2360 27380 2420
rect 26900 2340 27380 2360
rect 23460 980 23940 1000
rect 23460 920 23510 980
rect 23880 920 23940 980
rect 23460 850 23490 920
rect 23890 850 23940 920
rect 23460 810 23510 850
rect 23880 810 23940 850
rect 23460 740 23490 810
rect 23890 740 23940 810
rect 23460 710 23940 740
rect 25860 980 26340 1000
rect 25860 920 25910 980
rect 26280 920 26340 980
rect 25860 850 25890 920
rect 26290 850 26340 920
rect 25860 810 25910 850
rect 26280 810 26340 850
rect 25860 740 25890 810
rect 26290 740 26340 810
rect 25860 710 26340 740
rect 21800 -920 21820 -850
rect 21890 -920 21930 -850
rect 22000 -920 22060 -850
rect 21800 -960 22060 -920
rect 21800 -1030 21820 -960
rect 21890 -1030 21930 -960
rect 22000 -1030 22060 -960
rect 21800 -1070 22060 -1030
rect 21800 -1140 21820 -1070
rect 21890 -1140 21930 -1070
rect 22000 -1140 22060 -1070
rect 21800 -1180 22060 -1140
rect 21800 -1250 21820 -1180
rect 21890 -1250 21930 -1180
rect 22000 -1250 22060 -1180
rect 21800 -1290 22060 -1250
rect 21800 -1360 21820 -1290
rect 21890 -1360 21930 -1290
rect 22000 -1360 22060 -1290
rect 21800 -1400 22060 -1360
rect 21800 -1470 21820 -1400
rect 21890 -1470 21930 -1400
rect 22000 -1470 22060 -1400
rect 21800 -1510 22060 -1470
rect 21800 -1580 21820 -1510
rect 21890 -1580 21930 -1510
rect 22000 -1580 22060 -1510
rect 21800 -1620 22060 -1580
rect 21800 -1690 21820 -1620
rect 21890 -1690 21930 -1620
rect 22000 -1690 22060 -1620
rect 21800 -1730 22060 -1690
rect 21800 -1800 21820 -1730
rect 21890 -1800 21930 -1730
rect 22000 -1800 22060 -1730
rect 21800 -1840 22060 -1800
rect 21800 -1910 21820 -1840
rect 21890 -1910 21930 -1840
rect 22000 -1910 22060 -1840
rect 21800 -1950 22060 -1910
rect 21800 -2020 21820 -1950
rect 21890 -2020 21930 -1950
rect 22000 -2020 22060 -1950
rect 21800 -2040 22060 -2020
rect 24720 -3050 25050 -3030
rect 24720 -3120 24740 -3050
rect 24810 -3120 24850 -3050
rect 24920 -3120 24960 -3050
rect 25030 -3120 25050 -3050
rect 24720 -3125 25050 -3120
rect 30344 -3125 30477 3103
rect 31100 3210 37860 3300
rect 31100 2970 31180 3210
rect 31420 2970 31510 3210
rect 31750 2970 31840 3210
rect 32080 2970 32170 3210
rect 32410 2970 32500 3210
rect 32740 2970 32830 3210
rect 33070 2970 33160 3210
rect 33400 2970 33490 3210
rect 33730 2970 33820 3210
rect 34060 2970 34150 3210
rect 34390 2970 34480 3210
rect 34720 2970 34810 3210
rect 35050 2970 35140 3210
rect 35380 2970 35470 3210
rect 35710 2970 35800 3210
rect 36040 2970 36130 3210
rect 36370 2970 36460 3210
rect 36700 2970 36790 3210
rect 37030 2970 37120 3210
rect 37360 2970 37450 3210
rect 37690 2970 37860 3210
rect 31100 2880 37860 2970
rect 31100 2640 31180 2880
rect 31420 2640 31510 2880
rect 31750 2640 31840 2880
rect 32080 2640 32170 2880
rect 32410 2640 32500 2880
rect 32740 2640 32830 2880
rect 33070 2640 33160 2880
rect 33400 2640 33490 2880
rect 33730 2640 33820 2880
rect 34060 2640 34150 2880
rect 34390 2640 34480 2880
rect 34720 2640 34810 2880
rect 35050 2640 35140 2880
rect 35380 2640 35470 2880
rect 35710 2640 35800 2880
rect 36040 2640 36130 2880
rect 36370 2640 36460 2880
rect 36700 2640 36790 2880
rect 37030 2640 37120 2880
rect 37360 2640 37450 2880
rect 37690 2640 37860 2880
rect 31100 2550 37860 2640
rect 31100 2310 31180 2550
rect 31420 2310 31510 2550
rect 31750 2310 31840 2550
rect 32080 2310 32170 2550
rect 32410 2310 32500 2550
rect 32740 2310 32830 2550
rect 33070 2310 33160 2550
rect 33400 2310 33490 2550
rect 33730 2310 33820 2550
rect 34060 2310 34150 2550
rect 34390 2310 34480 2550
rect 34720 2310 34810 2550
rect 35050 2310 35140 2550
rect 35380 2310 35470 2550
rect 35710 2310 35800 2550
rect 36040 2310 36130 2550
rect 36370 2310 36460 2550
rect 36700 2310 36790 2550
rect 37030 2310 37120 2550
rect 37360 2310 37450 2550
rect 37690 2310 37860 2550
rect 31100 2220 37860 2310
rect 31100 1980 31180 2220
rect 31420 1980 31510 2220
rect 31750 1980 31840 2220
rect 32080 1980 32170 2220
rect 32410 1980 32500 2220
rect 32740 1980 32830 2220
rect 33070 1980 33160 2220
rect 33400 1980 33490 2220
rect 33730 1980 33820 2220
rect 34060 1980 34150 2220
rect 34390 1980 34480 2220
rect 34720 1980 34810 2220
rect 35050 1980 35140 2220
rect 35380 1980 35470 2220
rect 35710 1980 35800 2220
rect 36040 1980 36130 2220
rect 36370 1980 36460 2220
rect 36700 1980 36790 2220
rect 37030 1980 37120 2220
rect 37360 1980 37450 2220
rect 37690 1980 37860 2220
rect 31100 1890 37860 1980
rect 31100 1650 31180 1890
rect 31420 1650 31510 1890
rect 31750 1650 31840 1890
rect 32080 1650 32170 1890
rect 32410 1650 32500 1890
rect 32740 1650 32830 1890
rect 33070 1650 33160 1890
rect 33400 1650 33490 1890
rect 33730 1650 33820 1890
rect 34060 1650 34150 1890
rect 34390 1650 34480 1890
rect 34720 1650 34810 1890
rect 35050 1650 35140 1890
rect 35380 1650 35470 1890
rect 35710 1650 35800 1890
rect 36040 1650 36130 1890
rect 36370 1650 36460 1890
rect 36700 1650 36790 1890
rect 37030 1650 37120 1890
rect 37360 1650 37450 1890
rect 37690 1650 37860 1890
rect 31100 1560 37860 1650
rect 31100 1320 31180 1560
rect 31420 1320 31510 1560
rect 31750 1320 31840 1560
rect 32080 1320 32170 1560
rect 32410 1320 32500 1560
rect 32740 1320 32830 1560
rect 33070 1320 33160 1560
rect 33400 1320 33490 1560
rect 33730 1320 33820 1560
rect 34060 1320 34150 1560
rect 34390 1320 34480 1560
rect 34720 1320 34810 1560
rect 35050 1320 35140 1560
rect 35380 1320 35470 1560
rect 35710 1320 35800 1560
rect 36040 1320 36130 1560
rect 36370 1320 36460 1560
rect 36700 1320 36790 1560
rect 37030 1320 37120 1560
rect 37360 1320 37450 1560
rect 37690 1320 37860 1560
rect 31100 1150 37860 1320
rect 38180 7820 38500 7910
rect 38180 7750 38190 7820
rect 38260 7770 38280 7820
rect 38350 7770 38370 7820
rect 38440 7770 38500 7820
rect 38180 7730 38230 7750
rect 38180 7660 38190 7730
rect 38180 7640 38230 7660
rect 38180 7570 38190 7640
rect 38180 7550 38230 7570
rect 38180 7480 38190 7550
rect 38470 7530 38500 7770
rect 38260 7480 38280 7530
rect 38350 7480 38370 7530
rect 38440 7480 38500 7530
rect 38180 7460 38500 7480
rect 38180 7390 38190 7460
rect 38260 7440 38280 7460
rect 38350 7440 38370 7460
rect 38440 7440 38500 7460
rect 38180 7370 38230 7390
rect 38180 7300 38190 7370
rect 38180 7280 38230 7300
rect 38180 7210 38190 7280
rect 38180 7200 38230 7210
rect 38470 7200 38500 7440
rect 38180 7150 38500 7200
rect 38180 7080 38190 7150
rect 38260 7080 38280 7150
rect 38350 7080 38370 7150
rect 38440 7080 38500 7150
rect 38180 7070 38500 7080
rect 38180 7060 38230 7070
rect 38180 6990 38190 7060
rect 38180 6970 38230 6990
rect 38180 6900 38190 6970
rect 38180 6880 38230 6900
rect 38180 6810 38190 6880
rect 38470 6830 38500 7070
rect 38260 6810 38280 6830
rect 38350 6810 38370 6830
rect 38440 6810 38500 6830
rect 38180 6790 38500 6810
rect 38180 6720 38190 6790
rect 38260 6740 38280 6790
rect 38350 6740 38370 6790
rect 38440 6740 38500 6790
rect 38180 6700 38230 6720
rect 38180 6630 38190 6700
rect 38180 6610 38230 6630
rect 38180 6540 38190 6610
rect 38180 6520 38230 6540
rect 38180 6450 38190 6520
rect 38470 6500 38500 6740
rect 38260 6450 38280 6500
rect 38350 6450 38370 6500
rect 38440 6450 38500 6500
rect 38180 6430 38500 6450
rect 38180 6360 38190 6430
rect 38260 6410 38280 6430
rect 38350 6410 38370 6430
rect 38440 6410 38500 6430
rect 38180 6340 38230 6360
rect 38180 6270 38190 6340
rect 38180 6250 38230 6270
rect 38180 6180 38190 6250
rect 38180 6170 38230 6180
rect 38470 6170 38500 6410
rect 38180 6160 38500 6170
rect 38180 6090 38190 6160
rect 38260 6090 38280 6160
rect 38350 6090 38370 6160
rect 38440 6090 38500 6160
rect 38180 6080 38500 6090
rect 38180 6070 38230 6080
rect 38180 6000 38190 6070
rect 38180 5980 38230 6000
rect 38180 5910 38190 5980
rect 38180 5890 38230 5910
rect 38180 5820 38190 5890
rect 38470 5840 38500 6080
rect 38260 5820 38280 5840
rect 38350 5820 38370 5840
rect 38440 5820 38500 5840
rect 38180 5800 38500 5820
rect 38180 5730 38190 5800
rect 38260 5750 38280 5800
rect 38350 5750 38370 5800
rect 38440 5750 38500 5800
rect 38180 5710 38230 5730
rect 38180 5640 38190 5710
rect 38180 5620 38230 5640
rect 38180 5550 38190 5620
rect 38180 5530 38230 5550
rect 38180 5460 38190 5530
rect 38470 5510 38500 5750
rect 38260 5460 38280 5510
rect 38350 5460 38370 5510
rect 38440 5460 38500 5510
rect 38180 5440 38500 5460
rect 38180 5370 38190 5440
rect 38260 5420 38280 5440
rect 38350 5420 38370 5440
rect 38440 5420 38500 5440
rect 38180 5350 38230 5370
rect 38180 5280 38190 5350
rect 38180 5260 38230 5280
rect 38180 5190 38190 5260
rect 38180 5180 38230 5190
rect 38470 5180 38500 5420
rect 38180 5170 38500 5180
rect 38180 5100 38190 5170
rect 38260 5100 38280 5170
rect 38350 5100 38370 5170
rect 38440 5100 38500 5170
rect 38180 5090 38500 5100
rect 38180 5080 38230 5090
rect 38180 5010 38190 5080
rect 38180 4990 38230 5010
rect 38180 4920 38190 4990
rect 38180 4900 38230 4920
rect 38180 4830 38190 4900
rect 38470 4850 38500 5090
rect 38260 4830 38280 4850
rect 38350 4830 38370 4850
rect 38440 4830 38500 4850
rect 38180 4810 38500 4830
rect 38180 4740 38190 4810
rect 38260 4760 38280 4810
rect 38350 4760 38370 4810
rect 38440 4760 38500 4810
rect 38180 4720 38230 4740
rect 38180 4650 38190 4720
rect 38180 4630 38230 4650
rect 38180 4560 38190 4630
rect 38180 4540 38230 4560
rect 38180 4470 38190 4540
rect 38470 4520 38500 4760
rect 38260 4470 38280 4520
rect 38350 4470 38370 4520
rect 38440 4470 38500 4520
rect 38180 4450 38500 4470
rect 38180 4380 38190 4450
rect 38260 4430 38280 4450
rect 38350 4430 38370 4450
rect 38440 4430 38500 4450
rect 38180 4360 38230 4380
rect 38180 4290 38190 4360
rect 38180 4270 38230 4290
rect 38180 4200 38190 4270
rect 38180 4190 38230 4200
rect 38470 4190 38500 4430
rect 38180 4140 38500 4190
rect 38180 4070 38190 4140
rect 38260 4070 38280 4140
rect 38350 4070 38370 4140
rect 38440 4070 38500 4140
rect 38180 4060 38500 4070
rect 38180 4050 38230 4060
rect 38180 3980 38190 4050
rect 38180 3960 38230 3980
rect 38180 3890 38190 3960
rect 38180 3870 38230 3890
rect 38180 3800 38190 3870
rect 38470 3820 38500 4060
rect 38260 3800 38280 3820
rect 38350 3800 38370 3820
rect 38440 3800 38500 3820
rect 38180 3780 38500 3800
rect 38180 3710 38190 3780
rect 38260 3730 38280 3780
rect 38350 3730 38370 3780
rect 38440 3730 38500 3780
rect 38180 3690 38230 3710
rect 38180 3620 38190 3690
rect 38180 3600 38230 3620
rect 38180 3530 38190 3600
rect 38180 3510 38230 3530
rect 38180 3440 38190 3510
rect 38470 3490 38500 3730
rect 38260 3440 38280 3490
rect 38350 3440 38370 3490
rect 38440 3440 38500 3490
rect 38180 3420 38500 3440
rect 38180 3350 38190 3420
rect 38260 3400 38280 3420
rect 38350 3400 38370 3420
rect 38440 3400 38500 3420
rect 38180 3330 38230 3350
rect 38180 3260 38190 3330
rect 38180 3240 38230 3260
rect 38180 3170 38190 3240
rect 38180 3160 38230 3170
rect 38470 3160 38500 3400
rect 38180 3150 38500 3160
rect 38180 3080 38190 3150
rect 38260 3080 38280 3150
rect 38350 3080 38370 3150
rect 38440 3080 38500 3150
rect 38180 3070 38500 3080
rect 38180 3060 38230 3070
rect 38180 2990 38190 3060
rect 38180 2970 38230 2990
rect 38180 2900 38190 2970
rect 38180 2880 38230 2900
rect 38180 2810 38190 2880
rect 38470 2830 38500 3070
rect 38260 2810 38280 2830
rect 38350 2810 38370 2830
rect 38440 2810 38500 2830
rect 38180 2790 38500 2810
rect 38180 2720 38190 2790
rect 38260 2740 38280 2790
rect 38350 2740 38370 2790
rect 38440 2740 38500 2790
rect 38180 2700 38230 2720
rect 38180 2630 38190 2700
rect 38180 2610 38230 2630
rect 38180 2540 38190 2610
rect 38180 2520 38230 2540
rect 38180 2450 38190 2520
rect 38470 2500 38500 2740
rect 38260 2450 38280 2500
rect 38350 2450 38370 2500
rect 38440 2450 38500 2500
rect 38180 2430 38500 2450
rect 38180 2360 38190 2430
rect 38260 2410 38280 2430
rect 38350 2410 38370 2430
rect 38440 2410 38500 2430
rect 38180 2340 38230 2360
rect 38180 2270 38190 2340
rect 38180 2250 38230 2270
rect 38180 2180 38190 2250
rect 38180 2170 38230 2180
rect 38470 2170 38500 2410
rect 38180 2160 38500 2170
rect 38180 2090 38190 2160
rect 38260 2090 38280 2160
rect 38350 2090 38370 2160
rect 38440 2090 38500 2160
rect 38180 2080 38500 2090
rect 38180 2070 38230 2080
rect 38180 2000 38190 2070
rect 38180 1980 38230 2000
rect 38180 1910 38190 1980
rect 38180 1890 38230 1910
rect 38180 1820 38190 1890
rect 38470 1840 38500 2080
rect 38260 1820 38280 1840
rect 38350 1820 38370 1840
rect 38440 1820 38500 1840
rect 38180 1800 38500 1820
rect 38180 1730 38190 1800
rect 38260 1750 38280 1800
rect 38350 1750 38370 1800
rect 38440 1750 38500 1800
rect 38180 1710 38230 1730
rect 38180 1640 38190 1710
rect 38180 1620 38230 1640
rect 38180 1550 38190 1620
rect 38180 1530 38230 1550
rect 38180 1460 38190 1530
rect 38470 1510 38500 1750
rect 38260 1460 38280 1510
rect 38350 1460 38370 1510
rect 38440 1460 38500 1510
rect 38180 1440 38500 1460
rect 38180 1370 38190 1440
rect 38260 1420 38280 1440
rect 38350 1420 38370 1440
rect 38440 1420 38500 1440
rect 38180 1350 38230 1370
rect 38180 1280 38190 1350
rect 38180 1260 38230 1280
rect 38180 1190 38190 1260
rect 38180 1180 38230 1190
rect 38470 1180 38500 1420
rect 38180 1150 38500 1180
rect 31100 230 37860 310
rect 31100 20 31180 230
rect 30720 0 31180 20
rect 30720 -70 30740 0
rect 30810 -70 30850 0
rect 30920 -10 31180 0
rect 31420 -10 31510 230
rect 31750 -10 31840 230
rect 32080 -10 32170 230
rect 32410 -10 32500 230
rect 32740 -10 32830 230
rect 33070 -10 33160 230
rect 33400 -10 33490 230
rect 33730 -10 33820 230
rect 34060 -10 34150 230
rect 34390 -10 34480 230
rect 34720 -10 34810 230
rect 35050 -10 35140 230
rect 35380 -10 35470 230
rect 35710 -10 35800 230
rect 36040 -10 36130 230
rect 36370 -10 36460 230
rect 36700 -10 36790 230
rect 37030 -10 37120 230
rect 37360 -10 37450 230
rect 37690 -10 37860 230
rect 30920 -70 37860 -10
rect 30720 -100 37860 -70
rect 30720 -130 31180 -100
rect 30720 -200 30740 -130
rect 30810 -200 30850 -130
rect 30920 -200 31180 -130
rect 30720 -260 31180 -200
rect 30720 -330 30740 -260
rect 30810 -330 30850 -260
rect 30920 -330 31180 -260
rect 30720 -340 31180 -330
rect 31420 -340 31510 -100
rect 31750 -340 31840 -100
rect 32080 -340 32170 -100
rect 32410 -340 32500 -100
rect 32740 -340 32830 -100
rect 33070 -340 33160 -100
rect 33400 -340 33490 -100
rect 33730 -340 33820 -100
rect 34060 -340 34150 -100
rect 34390 -340 34480 -100
rect 34720 -340 34810 -100
rect 35050 -340 35140 -100
rect 35380 -340 35470 -100
rect 35710 -340 35800 -100
rect 36040 -340 36130 -100
rect 36370 -340 36460 -100
rect 36700 -340 36790 -100
rect 37030 -340 37120 -100
rect 37360 -340 37450 -100
rect 37690 -340 37860 -100
rect 30720 -350 37860 -340
rect 24720 -3160 30477 -3125
rect 24720 -3230 24740 -3160
rect 24810 -3230 24850 -3160
rect 24920 -3230 24960 -3160
rect 25030 -3230 30477 -3160
rect 24720 -3258 30477 -3230
rect 24720 -3270 25050 -3258
rect 24720 -3340 24740 -3270
rect 24810 -3340 24850 -3270
rect 24920 -3340 24960 -3270
rect 25030 -3340 25050 -3270
rect 24720 -3360 25050 -3340
rect 22420 -3690 22900 -3660
rect 22420 -3760 22470 -3690
rect 22870 -3760 22900 -3690
rect 22420 -3800 22480 -3760
rect 22850 -3800 22900 -3760
rect 22420 -3870 22470 -3800
rect 22870 -3870 22900 -3800
rect 22420 -3930 22480 -3870
rect 22850 -3930 22900 -3870
rect 22420 -3950 22900 -3930
rect 26900 -3690 27380 -3660
rect 26900 -3760 26950 -3690
rect 27350 -3760 27380 -3690
rect 26900 -3800 26960 -3760
rect 27330 -3800 27380 -3760
rect 26900 -3870 26950 -3800
rect 27350 -3870 27380 -3800
rect 26900 -3930 26960 -3870
rect 27330 -3930 27380 -3870
rect 26900 -3950 27380 -3930
rect 26400 -5890 26880 -5780
rect 26400 -5915 26510 -5890
rect 18975 -6025 26510 -5915
rect -1200 -6330 90 -6320
rect -1200 -6370 -1160 -6330
rect -1090 -6370 -1070 -6330
rect -1000 -6370 -980 -6330
rect -1200 -6610 -1170 -6370
rect -910 -6400 -890 -6330
rect -820 -6370 -800 -6330
rect -730 -6370 -710 -6330
rect -640 -6370 -620 -6330
rect -550 -6400 -530 -6330
rect -460 -6370 -440 -6330
rect -370 -6370 -350 -6330
rect -280 -6370 -260 -6330
rect -270 -6400 -260 -6370
rect -190 -6370 -170 -6330
rect -100 -6370 -80 -6330
rect -10 -6370 10 -6330
rect -190 -6400 -180 -6370
rect 80 -6400 90 -6330
rect -930 -6420 -840 -6400
rect -600 -6420 -510 -6400
rect -270 -6420 -180 -6400
rect 60 -6420 90 -6400
rect -910 -6490 -890 -6420
rect -550 -6490 -530 -6420
rect -270 -6490 -260 -6420
rect -190 -6490 -180 -6420
rect 80 -6490 90 -6420
rect -930 -6510 -840 -6490
rect -600 -6510 -510 -6490
rect -270 -6510 -180 -6490
rect 60 -6510 90 -6490
rect -910 -6580 -890 -6510
rect -550 -6580 -530 -6510
rect -270 -6580 -260 -6510
rect -190 -6580 -180 -6510
rect 80 -6580 90 -6510
rect -930 -6610 -840 -6580
rect -600 -6610 -510 -6580
rect -270 -6610 -180 -6580
rect 60 -6610 90 -6580
rect -1200 -6640 90 -6610
rect 14690 -6330 15980 -6320
rect 14690 -6400 14700 -6330
rect 14770 -6370 14790 -6330
rect 14860 -6370 14880 -6330
rect 14950 -6370 14970 -6330
rect 14960 -6400 14970 -6370
rect 15040 -6370 15060 -6330
rect 15130 -6370 15150 -6330
rect 15220 -6370 15240 -6330
rect 15040 -6400 15050 -6370
rect 15310 -6400 15330 -6330
rect 15400 -6370 15420 -6330
rect 15490 -6370 15510 -6330
rect 15580 -6370 15600 -6330
rect 15670 -6400 15690 -6330
rect 15760 -6370 15780 -6330
rect 15850 -6370 15870 -6330
rect 15940 -6370 15980 -6330
rect 14690 -6420 14720 -6400
rect 14960 -6420 15050 -6400
rect 15290 -6420 15380 -6400
rect 15620 -6420 15710 -6400
rect 14690 -6490 14700 -6420
rect 14960 -6490 14970 -6420
rect 15040 -6490 15050 -6420
rect 15310 -6490 15330 -6420
rect 15670 -6490 15690 -6420
rect 14690 -6510 14720 -6490
rect 14960 -6510 15050 -6490
rect 15290 -6510 15380 -6490
rect 15620 -6510 15710 -6490
rect 14690 -6580 14700 -6510
rect 14960 -6580 14970 -6510
rect 15040 -6580 15050 -6510
rect 15310 -6580 15330 -6510
rect 15670 -6580 15690 -6510
rect 14690 -6610 14720 -6580
rect 14960 -6610 15050 -6580
rect 15290 -6610 15380 -6580
rect 15620 -6610 15710 -6580
rect 15950 -6610 15980 -6370
rect 14690 -6640 15980 -6610
rect 14590 -8230 14900 -8210
rect 14590 -8300 14600 -8230
rect 14670 -8300 14700 -8230
rect 14770 -8300 14810 -8230
rect 14880 -8300 14900 -8230
rect 14590 -8325 14900 -8300
rect 18975 -8325 19085 -6025
rect 14590 -8340 19085 -8325
rect 14590 -8410 14600 -8340
rect 14670 -8410 14700 -8340
rect 14770 -8410 14810 -8340
rect 14880 -8410 19085 -8340
rect 14590 -8435 19085 -8410
rect 21610 -8360 21930 -8330
rect 21610 -8430 21630 -8360
rect 21700 -8370 21730 -8360
rect 21800 -8370 21830 -8360
rect 21900 -8430 21930 -8360
rect 14590 -8450 14900 -8435
rect 14590 -8520 14600 -8450
rect 14670 -8520 14700 -8450
rect 14770 -8520 14810 -8450
rect 14880 -8520 14900 -8450
rect 14590 -8540 14900 -8520
rect 21610 -8460 21650 -8430
rect 21890 -8460 21930 -8430
rect 21610 -8530 21630 -8460
rect 21900 -8530 21930 -8460
rect 21610 -8560 21650 -8530
rect 21890 -8560 21930 -8530
rect 21610 -8630 21630 -8560
rect 21700 -8630 21730 -8610
rect 21800 -8630 21830 -8610
rect 21900 -8630 21930 -8560
rect 21610 -8650 21930 -8630
rect 22630 -9010 22950 -8980
rect 22630 -9080 22650 -9010
rect 22720 -9080 22750 -9010
rect 22820 -9080 22850 -9010
rect 22920 -9080 22950 -9010
rect 22630 -9110 22950 -9080
rect 22630 -9180 22650 -9110
rect 22720 -9180 22750 -9110
rect 22820 -9180 22850 -9110
rect 22920 -9180 22950 -9110
rect 22630 -9210 22950 -9180
rect 22630 -9280 22650 -9210
rect 22720 -9280 22750 -9210
rect 22820 -9280 22850 -9210
rect 22920 -9280 22950 -9210
rect 1080 -10340 2680 -10310
rect 1080 -10410 1150 -10340
rect 1220 -10410 1260 -10340
rect 1550 -10410 1590 -10340
rect 1880 -10410 1920 -10340
rect 2210 -10410 2250 -10340
rect 2540 -10410 2580 -10340
rect 2650 -10410 2680 -10340
rect 1080 -10450 1260 -10410
rect 1500 -10450 1590 -10410
rect 1830 -10450 1930 -10410
rect 2170 -10450 2260 -10410
rect 2500 -10450 2680 -10410
rect 1080 -10520 1150 -10450
rect 1220 -10520 1260 -10450
rect 1550 -10520 1590 -10450
rect 1880 -10520 1920 -10450
rect 2210 -10520 2250 -10450
rect 2540 -10520 2580 -10450
rect 2650 -10520 2680 -10450
rect 1080 -10580 1260 -10520
rect 1500 -10580 1590 -10520
rect 1830 -10580 1930 -10520
rect 2170 -10580 2260 -10520
rect 2500 -10580 2680 -10520
rect 1080 -10600 2680 -10580
rect 12220 -10370 13820 -10340
rect 12220 -10440 12290 -10370
rect 12360 -10440 12400 -10370
rect 12690 -10440 12730 -10370
rect 13020 -10440 13060 -10370
rect 13350 -10440 13390 -10370
rect 13680 -10440 13720 -10370
rect 13790 -10440 13820 -10370
rect 12220 -10480 12400 -10440
rect 12640 -10480 12730 -10440
rect 12970 -10480 13070 -10440
rect 13310 -10480 13400 -10440
rect 13640 -10480 13820 -10440
rect 12220 -10550 12290 -10480
rect 12360 -10550 12400 -10480
rect 12690 -10550 12730 -10480
rect 13020 -10550 13060 -10480
rect 13350 -10550 13390 -10480
rect 13680 -10550 13720 -10480
rect 13790 -10550 13820 -10480
rect 12220 -10610 12400 -10550
rect 12640 -10610 12730 -10550
rect 12970 -10610 13070 -10550
rect 13310 -10610 13400 -10550
rect 13640 -10610 13820 -10550
rect 12220 -10620 13820 -10610
rect 22630 -10510 22950 -9280
rect 22630 -10520 30080 -10510
rect 22630 -10590 29990 -10520
rect 30060 -10590 30080 -10520
rect 22630 -10630 30080 -10590
rect 22630 -10700 29990 -10630
rect 30060 -10700 30080 -10630
rect 22630 -10740 30080 -10700
rect 22630 -10810 29990 -10740
rect 30060 -10810 30080 -10740
rect 22630 -10830 30080 -10810
rect 30344 -10995 30477 -3258
rect 31100 -430 37860 -350
rect 31100 -670 31180 -430
rect 31420 -670 31510 -430
rect 31750 -670 31840 -430
rect 32080 -670 32170 -430
rect 32410 -670 32500 -430
rect 32740 -670 32830 -430
rect 33070 -670 33160 -430
rect 33400 -670 33490 -430
rect 33730 -670 33820 -430
rect 34060 -670 34150 -430
rect 34390 -670 34480 -430
rect 34720 -670 34810 -430
rect 35050 -670 35140 -430
rect 35380 -670 35470 -430
rect 35710 -670 35800 -430
rect 36040 -670 36130 -430
rect 36370 -670 36460 -430
rect 36700 -670 36790 -430
rect 37030 -670 37120 -430
rect 37360 -670 37450 -430
rect 37690 -670 37860 -430
rect 31100 -760 37860 -670
rect 31100 -1000 31180 -760
rect 31420 -1000 31510 -760
rect 31750 -1000 31840 -760
rect 32080 -1000 32170 -760
rect 32410 -1000 32500 -760
rect 32740 -1000 32830 -760
rect 33070 -1000 33160 -760
rect 33400 -1000 33490 -760
rect 33730 -1000 33820 -760
rect 34060 -1000 34150 -760
rect 34390 -1000 34480 -760
rect 34720 -1000 34810 -760
rect 35050 -1000 35140 -760
rect 35380 -1000 35470 -760
rect 35710 -1000 35800 -760
rect 36040 -1000 36130 -760
rect 36370 -1000 36460 -760
rect 36700 -1000 36790 -760
rect 37030 -1000 37120 -760
rect 37360 -1000 37450 -760
rect 37690 -1000 37860 -760
rect 31100 -1090 37860 -1000
rect 31100 -1330 31180 -1090
rect 31420 -1330 31510 -1090
rect 31750 -1330 31840 -1090
rect 32080 -1330 32170 -1090
rect 32410 -1330 32500 -1090
rect 32740 -1330 32830 -1090
rect 33070 -1330 33160 -1090
rect 33400 -1330 33490 -1090
rect 33730 -1330 33820 -1090
rect 34060 -1330 34150 -1090
rect 34390 -1330 34480 -1090
rect 34720 -1330 34810 -1090
rect 35050 -1330 35140 -1090
rect 35380 -1330 35470 -1090
rect 35710 -1330 35800 -1090
rect 36040 -1330 36130 -1090
rect 36370 -1330 36460 -1090
rect 36700 -1330 36790 -1090
rect 37030 -1330 37120 -1090
rect 37360 -1330 37450 -1090
rect 37690 -1330 37860 -1090
rect 31100 -1420 37860 -1330
rect 31100 -1660 31180 -1420
rect 31420 -1660 31510 -1420
rect 31750 -1660 31840 -1420
rect 32080 -1660 32170 -1420
rect 32410 -1660 32500 -1420
rect 32740 -1660 32830 -1420
rect 33070 -1660 33160 -1420
rect 33400 -1660 33490 -1420
rect 33730 -1660 33820 -1420
rect 34060 -1660 34150 -1420
rect 34390 -1660 34480 -1420
rect 34720 -1660 34810 -1420
rect 35050 -1660 35140 -1420
rect 35380 -1660 35470 -1420
rect 35710 -1660 35800 -1420
rect 36040 -1660 36130 -1420
rect 36370 -1660 36460 -1420
rect 36700 -1660 36790 -1420
rect 37030 -1660 37120 -1420
rect 37360 -1660 37450 -1420
rect 37690 -1660 37860 -1420
rect 31100 -1750 37860 -1660
rect 31100 -1990 31180 -1750
rect 31420 -1990 31510 -1750
rect 31750 -1990 31840 -1750
rect 32080 -1990 32170 -1750
rect 32410 -1990 32500 -1750
rect 32740 -1990 32830 -1750
rect 33070 -1990 33160 -1750
rect 33400 -1990 33490 -1750
rect 33730 -1990 33820 -1750
rect 34060 -1990 34150 -1750
rect 34390 -1990 34480 -1750
rect 34720 -1990 34810 -1750
rect 35050 -1990 35140 -1750
rect 35380 -1990 35470 -1750
rect 35710 -1990 35800 -1750
rect 36040 -1990 36130 -1750
rect 36370 -1990 36460 -1750
rect 36700 -1990 36790 -1750
rect 37030 -1990 37120 -1750
rect 37360 -1990 37450 -1750
rect 37690 -1990 37860 -1750
rect 31100 -2080 37860 -1990
rect 31100 -2320 31180 -2080
rect 31420 -2320 31510 -2080
rect 31750 -2320 31840 -2080
rect 32080 -2320 32170 -2080
rect 32410 -2320 32500 -2080
rect 32740 -2320 32830 -2080
rect 33070 -2320 33160 -2080
rect 33400 -2320 33490 -2080
rect 33730 -2320 33820 -2080
rect 34060 -2320 34150 -2080
rect 34390 -2320 34480 -2080
rect 34720 -2320 34810 -2080
rect 35050 -2320 35140 -2080
rect 35380 -2320 35470 -2080
rect 35710 -2320 35800 -2080
rect 36040 -2320 36130 -2080
rect 36370 -2320 36460 -2080
rect 36700 -2320 36790 -2080
rect 37030 -2320 37120 -2080
rect 37360 -2320 37450 -2080
rect 37690 -2320 37860 -2080
rect 31100 -2410 37860 -2320
rect 31100 -2650 31180 -2410
rect 31420 -2650 31510 -2410
rect 31750 -2650 31840 -2410
rect 32080 -2650 32170 -2410
rect 32410 -2650 32500 -2410
rect 32740 -2650 32830 -2410
rect 33070 -2650 33160 -2410
rect 33400 -2650 33490 -2410
rect 33730 -2650 33820 -2410
rect 34060 -2650 34150 -2410
rect 34390 -2650 34480 -2410
rect 34720 -2650 34810 -2410
rect 35050 -2650 35140 -2410
rect 35380 -2650 35470 -2410
rect 35710 -2650 35800 -2410
rect 36040 -2650 36130 -2410
rect 36370 -2650 36460 -2410
rect 36700 -2650 36790 -2410
rect 37030 -2650 37120 -2410
rect 37360 -2650 37450 -2410
rect 37690 -2650 37860 -2410
rect 31100 -2740 37860 -2650
rect 31100 -2980 31180 -2740
rect 31420 -2980 31510 -2740
rect 31750 -2980 31840 -2740
rect 32080 -2980 32170 -2740
rect 32410 -2980 32500 -2740
rect 32740 -2980 32830 -2740
rect 33070 -2980 33160 -2740
rect 33400 -2980 33490 -2740
rect 33730 -2980 33820 -2740
rect 34060 -2980 34150 -2740
rect 34390 -2980 34480 -2740
rect 34720 -2980 34810 -2740
rect 35050 -2980 35140 -2740
rect 35380 -2980 35470 -2740
rect 35710 -2980 35800 -2740
rect 36040 -2980 36130 -2740
rect 36370 -2980 36460 -2740
rect 36700 -2980 36790 -2740
rect 37030 -2980 37120 -2740
rect 37360 -2980 37450 -2740
rect 37690 -2980 37860 -2740
rect 31100 -3070 37860 -2980
rect 31100 -3310 31180 -3070
rect 31420 -3310 31510 -3070
rect 31750 -3310 31840 -3070
rect 32080 -3310 32170 -3070
rect 32410 -3310 32500 -3070
rect 32740 -3310 32830 -3070
rect 33070 -3310 33160 -3070
rect 33400 -3310 33490 -3070
rect 33730 -3310 33820 -3070
rect 34060 -3310 34150 -3070
rect 34390 -3310 34480 -3070
rect 34720 -3310 34810 -3070
rect 35050 -3310 35140 -3070
rect 35380 -3310 35470 -3070
rect 35710 -3310 35800 -3070
rect 36040 -3310 36130 -3070
rect 36370 -3310 36460 -3070
rect 36700 -3310 36790 -3070
rect 37030 -3310 37120 -3070
rect 37360 -3310 37450 -3070
rect 37690 -3310 37860 -3070
rect 31100 -3400 37860 -3310
rect 31100 -3640 31180 -3400
rect 31420 -3640 31510 -3400
rect 31750 -3640 31840 -3400
rect 32080 -3640 32170 -3400
rect 32410 -3640 32500 -3400
rect 32740 -3640 32830 -3400
rect 33070 -3640 33160 -3400
rect 33400 -3640 33490 -3400
rect 33730 -3640 33820 -3400
rect 34060 -3640 34150 -3400
rect 34390 -3640 34480 -3400
rect 34720 -3640 34810 -3400
rect 35050 -3640 35140 -3400
rect 35380 -3640 35470 -3400
rect 35710 -3640 35800 -3400
rect 36040 -3640 36130 -3400
rect 36370 -3640 36460 -3400
rect 36700 -3640 36790 -3400
rect 37030 -3640 37120 -3400
rect 37360 -3640 37450 -3400
rect 37690 -3640 37860 -3400
rect 31100 -3730 37860 -3640
rect 31100 -3970 31180 -3730
rect 31420 -3970 31510 -3730
rect 31750 -3970 31840 -3730
rect 32080 -3970 32170 -3730
rect 32410 -3970 32500 -3730
rect 32740 -3970 32830 -3730
rect 33070 -3970 33160 -3730
rect 33400 -3970 33490 -3730
rect 33730 -3970 33820 -3730
rect 34060 -3970 34150 -3730
rect 34390 -3970 34480 -3730
rect 34720 -3970 34810 -3730
rect 35050 -3970 35140 -3730
rect 35380 -3970 35470 -3730
rect 35710 -3970 35800 -3730
rect 36040 -3970 36130 -3730
rect 36370 -3970 36460 -3730
rect 36700 -3970 36790 -3730
rect 37030 -3970 37120 -3730
rect 37360 -3970 37450 -3730
rect 37690 -3970 37860 -3730
rect 31100 -4060 37860 -3970
rect 31100 -4300 31180 -4060
rect 31420 -4300 31510 -4060
rect 31750 -4300 31840 -4060
rect 32080 -4300 32170 -4060
rect 32410 -4300 32500 -4060
rect 32740 -4300 32830 -4060
rect 33070 -4300 33160 -4060
rect 33400 -4300 33490 -4060
rect 33730 -4300 33820 -4060
rect 34060 -4300 34150 -4060
rect 34390 -4300 34480 -4060
rect 34720 -4300 34810 -4060
rect 35050 -4300 35140 -4060
rect 35380 -4300 35470 -4060
rect 35710 -4300 35800 -4060
rect 36040 -4300 36130 -4060
rect 36370 -4300 36460 -4060
rect 36700 -4300 36790 -4060
rect 37030 -4300 37120 -4060
rect 37360 -4300 37450 -4060
rect 37690 -4300 37860 -4060
rect 31100 -4390 37860 -4300
rect 31100 -4630 31180 -4390
rect 31420 -4630 31510 -4390
rect 31750 -4630 31840 -4390
rect 32080 -4630 32170 -4390
rect 32410 -4630 32500 -4390
rect 32740 -4630 32830 -4390
rect 33070 -4630 33160 -4390
rect 33400 -4630 33490 -4390
rect 33730 -4630 33820 -4390
rect 34060 -4630 34150 -4390
rect 34390 -4630 34480 -4390
rect 34720 -4630 34810 -4390
rect 35050 -4630 35140 -4390
rect 35380 -4630 35470 -4390
rect 35710 -4630 35800 -4390
rect 36040 -4630 36130 -4390
rect 36370 -4630 36460 -4390
rect 36700 -4630 36790 -4390
rect 37030 -4630 37120 -4390
rect 37360 -4630 37450 -4390
rect 37690 -4630 37860 -4390
rect 31100 -4720 37860 -4630
rect 31100 -4960 31180 -4720
rect 31420 -4960 31510 -4720
rect 31750 -4960 31840 -4720
rect 32080 -4960 32170 -4720
rect 32410 -4960 32500 -4720
rect 32740 -4960 32830 -4720
rect 33070 -4960 33160 -4720
rect 33400 -4960 33490 -4720
rect 33730 -4960 33820 -4720
rect 34060 -4960 34150 -4720
rect 34390 -4960 34480 -4720
rect 34720 -4960 34810 -4720
rect 35050 -4960 35140 -4720
rect 35380 -4960 35470 -4720
rect 35710 -4960 35800 -4720
rect 36040 -4960 36130 -4720
rect 36370 -4960 36460 -4720
rect 36700 -4960 36790 -4720
rect 37030 -4960 37120 -4720
rect 37360 -4960 37450 -4720
rect 37690 -4960 37860 -4720
rect 31100 -5050 37860 -4960
rect 31100 -5290 31180 -5050
rect 31420 -5290 31510 -5050
rect 31750 -5290 31840 -5050
rect 32080 -5290 32170 -5050
rect 32410 -5290 32500 -5050
rect 32740 -5290 32830 -5050
rect 33070 -5290 33160 -5050
rect 33400 -5290 33490 -5050
rect 33730 -5290 33820 -5050
rect 34060 -5290 34150 -5050
rect 34390 -5290 34480 -5050
rect 34720 -5290 34810 -5050
rect 35050 -5290 35140 -5050
rect 35380 -5290 35470 -5050
rect 35710 -5290 35800 -5050
rect 36040 -5290 36130 -5050
rect 36370 -5290 36460 -5050
rect 36700 -5290 36790 -5050
rect 37030 -5290 37120 -5050
rect 37360 -5290 37450 -5050
rect 37690 -5290 37860 -5050
rect 31100 -5380 37860 -5290
rect 31100 -5620 31180 -5380
rect 31420 -5620 31510 -5380
rect 31750 -5620 31840 -5380
rect 32080 -5620 32170 -5380
rect 32410 -5620 32500 -5380
rect 32740 -5620 32830 -5380
rect 33070 -5620 33160 -5380
rect 33400 -5620 33490 -5380
rect 33730 -5620 33820 -5380
rect 34060 -5620 34150 -5380
rect 34390 -5620 34480 -5380
rect 34720 -5620 34810 -5380
rect 35050 -5620 35140 -5380
rect 35380 -5620 35470 -5380
rect 35710 -5620 35800 -5380
rect 36040 -5620 36130 -5380
rect 36370 -5620 36460 -5380
rect 36700 -5620 36790 -5380
rect 37030 -5620 37120 -5380
rect 37360 -5620 37450 -5380
rect 37690 -5620 37860 -5380
rect 31100 -5710 37860 -5620
rect 31100 -5950 31180 -5710
rect 31420 -5950 31510 -5710
rect 31750 -5950 31840 -5710
rect 32080 -5950 32170 -5710
rect 32410 -5950 32500 -5710
rect 32740 -5950 32830 -5710
rect 33070 -5950 33160 -5710
rect 33400 -5950 33490 -5710
rect 33730 -5950 33820 -5710
rect 34060 -5950 34150 -5710
rect 34390 -5950 34480 -5710
rect 34720 -5950 34810 -5710
rect 35050 -5950 35140 -5710
rect 35380 -5950 35470 -5710
rect 35710 -5950 35800 -5710
rect 36040 -5950 36130 -5710
rect 36370 -5950 36460 -5710
rect 36700 -5950 36790 -5710
rect 37030 -5950 37120 -5710
rect 37360 -5950 37450 -5710
rect 37690 -5950 37860 -5710
rect 31100 -6040 37860 -5950
rect 31100 -6280 31180 -6040
rect 31420 -6280 31510 -6040
rect 31750 -6280 31840 -6040
rect 32080 -6280 32170 -6040
rect 32410 -6280 32500 -6040
rect 32740 -6280 32830 -6040
rect 33070 -6280 33160 -6040
rect 33400 -6280 33490 -6040
rect 33730 -6280 33820 -6040
rect 34060 -6280 34150 -6040
rect 34390 -6280 34480 -6040
rect 34720 -6280 34810 -6040
rect 35050 -6280 35140 -6040
rect 35380 -6280 35470 -6040
rect 35710 -6280 35800 -6040
rect 36040 -6280 36130 -6040
rect 36370 -6280 36460 -6040
rect 36700 -6280 36790 -6040
rect 37030 -6280 37120 -6040
rect 37360 -6280 37450 -6040
rect 37690 -6280 37860 -6040
rect 31100 -6450 37860 -6280
rect 38180 220 38500 310
rect 38180 150 38190 220
rect 38260 170 38280 220
rect 38350 170 38370 220
rect 38440 170 38500 220
rect 38180 130 38230 150
rect 38180 60 38190 130
rect 38180 40 38230 60
rect 38180 -30 38190 40
rect 38180 -50 38230 -30
rect 38180 -120 38190 -50
rect 38470 -70 38500 170
rect 38260 -120 38280 -70
rect 38350 -120 38370 -70
rect 38440 -120 38500 -70
rect 38180 -140 38500 -120
rect 38180 -210 38190 -140
rect 38260 -160 38280 -140
rect 38350 -160 38370 -140
rect 38440 -160 38500 -140
rect 38180 -230 38230 -210
rect 38180 -300 38190 -230
rect 38180 -320 38230 -300
rect 38180 -390 38190 -320
rect 38180 -400 38230 -390
rect 38470 -400 38500 -160
rect 38180 -450 38500 -400
rect 38180 -520 38190 -450
rect 38260 -520 38280 -450
rect 38350 -520 38370 -450
rect 38440 -520 38500 -450
rect 38180 -530 38500 -520
rect 38180 -540 38230 -530
rect 38180 -610 38190 -540
rect 38180 -630 38230 -610
rect 38180 -700 38190 -630
rect 38180 -720 38230 -700
rect 38180 -790 38190 -720
rect 38470 -770 38500 -530
rect 38260 -790 38280 -770
rect 38350 -790 38370 -770
rect 38440 -790 38500 -770
rect 38180 -810 38500 -790
rect 38180 -880 38190 -810
rect 38260 -860 38280 -810
rect 38350 -860 38370 -810
rect 38440 -860 38500 -810
rect 38180 -900 38230 -880
rect 38180 -970 38190 -900
rect 38180 -990 38230 -970
rect 38180 -1060 38190 -990
rect 38180 -1080 38230 -1060
rect 38180 -1150 38190 -1080
rect 38470 -1100 38500 -860
rect 38260 -1150 38280 -1100
rect 38350 -1150 38370 -1100
rect 38440 -1150 38500 -1100
rect 38180 -1170 38500 -1150
rect 38180 -1240 38190 -1170
rect 38260 -1190 38280 -1170
rect 38350 -1190 38370 -1170
rect 38440 -1190 38500 -1170
rect 38180 -1260 38230 -1240
rect 38180 -1330 38190 -1260
rect 38180 -1350 38230 -1330
rect 38180 -1420 38190 -1350
rect 38180 -1430 38230 -1420
rect 38470 -1430 38500 -1190
rect 38180 -1440 38500 -1430
rect 38180 -1510 38190 -1440
rect 38260 -1510 38280 -1440
rect 38350 -1510 38370 -1440
rect 38440 -1510 38500 -1440
rect 38180 -1520 38500 -1510
rect 38180 -1530 38230 -1520
rect 38180 -1600 38190 -1530
rect 38180 -1620 38230 -1600
rect 38180 -1690 38190 -1620
rect 38180 -1710 38230 -1690
rect 38180 -1780 38190 -1710
rect 38470 -1760 38500 -1520
rect 38260 -1780 38280 -1760
rect 38350 -1780 38370 -1760
rect 38440 -1780 38500 -1760
rect 38180 -1800 38500 -1780
rect 38180 -1870 38190 -1800
rect 38260 -1850 38280 -1800
rect 38350 -1850 38370 -1800
rect 38440 -1850 38500 -1800
rect 38180 -1890 38230 -1870
rect 38180 -1960 38190 -1890
rect 38180 -1980 38230 -1960
rect 38180 -2050 38190 -1980
rect 38180 -2070 38230 -2050
rect 38180 -2140 38190 -2070
rect 38470 -2090 38500 -1850
rect 38260 -2140 38280 -2090
rect 38350 -2140 38370 -2090
rect 38440 -2140 38500 -2090
rect 38180 -2160 38500 -2140
rect 38180 -2230 38190 -2160
rect 38260 -2180 38280 -2160
rect 38350 -2180 38370 -2160
rect 38440 -2180 38500 -2160
rect 38180 -2250 38230 -2230
rect 38180 -2320 38190 -2250
rect 38180 -2340 38230 -2320
rect 38180 -2410 38190 -2340
rect 38180 -2420 38230 -2410
rect 38470 -2420 38500 -2180
rect 38180 -2430 38500 -2420
rect 38180 -2500 38190 -2430
rect 38260 -2500 38280 -2430
rect 38350 -2500 38370 -2430
rect 38440 -2500 38500 -2430
rect 38180 -2510 38500 -2500
rect 38180 -2520 38230 -2510
rect 38180 -2590 38190 -2520
rect 38180 -2610 38230 -2590
rect 38180 -2680 38190 -2610
rect 38180 -2700 38230 -2680
rect 38180 -2770 38190 -2700
rect 38470 -2750 38500 -2510
rect 38260 -2770 38280 -2750
rect 38350 -2770 38370 -2750
rect 38440 -2770 38500 -2750
rect 38180 -2790 38500 -2770
rect 38180 -2860 38190 -2790
rect 38260 -2840 38280 -2790
rect 38350 -2840 38370 -2790
rect 38440 -2840 38500 -2790
rect 38180 -2880 38230 -2860
rect 38180 -2950 38190 -2880
rect 38180 -2970 38230 -2950
rect 38180 -3040 38190 -2970
rect 38180 -3060 38230 -3040
rect 38180 -3130 38190 -3060
rect 38470 -3080 38500 -2840
rect 38260 -3130 38280 -3080
rect 38350 -3130 38370 -3080
rect 38440 -3130 38500 -3080
rect 38180 -3150 38500 -3130
rect 38180 -3220 38190 -3150
rect 38260 -3170 38280 -3150
rect 38350 -3170 38370 -3150
rect 38440 -3170 38500 -3150
rect 38180 -3240 38230 -3220
rect 38180 -3310 38190 -3240
rect 38180 -3330 38230 -3310
rect 38180 -3400 38190 -3330
rect 38180 -3410 38230 -3400
rect 38470 -3410 38500 -3170
rect 38180 -3460 38500 -3410
rect 38180 -3530 38190 -3460
rect 38260 -3530 38280 -3460
rect 38350 -3530 38370 -3460
rect 38440 -3530 38500 -3460
rect 38180 -3540 38500 -3530
rect 38180 -3550 38230 -3540
rect 38180 -3620 38190 -3550
rect 38180 -3640 38230 -3620
rect 38180 -3710 38190 -3640
rect 38180 -3730 38230 -3710
rect 38180 -3800 38190 -3730
rect 38470 -3780 38500 -3540
rect 38260 -3800 38280 -3780
rect 38350 -3800 38370 -3780
rect 38440 -3800 38500 -3780
rect 38180 -3820 38500 -3800
rect 38180 -3890 38190 -3820
rect 38260 -3870 38280 -3820
rect 38350 -3870 38370 -3820
rect 38440 -3870 38500 -3820
rect 38180 -3910 38230 -3890
rect 38180 -3980 38190 -3910
rect 38180 -4000 38230 -3980
rect 38180 -4070 38190 -4000
rect 38180 -4090 38230 -4070
rect 38180 -4160 38190 -4090
rect 38470 -4110 38500 -3870
rect 38260 -4160 38280 -4110
rect 38350 -4160 38370 -4110
rect 38440 -4160 38500 -4110
rect 38180 -4180 38500 -4160
rect 38180 -4250 38190 -4180
rect 38260 -4200 38280 -4180
rect 38350 -4200 38370 -4180
rect 38440 -4200 38500 -4180
rect 38180 -4270 38230 -4250
rect 38180 -4340 38190 -4270
rect 38180 -4360 38230 -4340
rect 38180 -4430 38190 -4360
rect 38180 -4440 38230 -4430
rect 38470 -4440 38500 -4200
rect 38180 -4450 38500 -4440
rect 38180 -4520 38190 -4450
rect 38260 -4520 38280 -4450
rect 38350 -4520 38370 -4450
rect 38440 -4520 38500 -4450
rect 38180 -4530 38500 -4520
rect 38180 -4540 38230 -4530
rect 38180 -4610 38190 -4540
rect 38180 -4630 38230 -4610
rect 38180 -4700 38190 -4630
rect 38180 -4720 38230 -4700
rect 38180 -4790 38190 -4720
rect 38470 -4770 38500 -4530
rect 38260 -4790 38280 -4770
rect 38350 -4790 38370 -4770
rect 38440 -4790 38500 -4770
rect 38180 -4810 38500 -4790
rect 38180 -4880 38190 -4810
rect 38260 -4860 38280 -4810
rect 38350 -4860 38370 -4810
rect 38440 -4860 38500 -4810
rect 38180 -4900 38230 -4880
rect 38180 -4970 38190 -4900
rect 38180 -4990 38230 -4970
rect 38180 -5060 38190 -4990
rect 38180 -5080 38230 -5060
rect 38180 -5150 38190 -5080
rect 38470 -5100 38500 -4860
rect 38260 -5150 38280 -5100
rect 38350 -5150 38370 -5100
rect 38440 -5150 38500 -5100
rect 38180 -5170 38500 -5150
rect 38180 -5240 38190 -5170
rect 38260 -5190 38280 -5170
rect 38350 -5190 38370 -5170
rect 38440 -5190 38500 -5170
rect 38180 -5260 38230 -5240
rect 38180 -5330 38190 -5260
rect 38180 -5350 38230 -5330
rect 38180 -5420 38190 -5350
rect 38180 -5430 38230 -5420
rect 38470 -5430 38500 -5190
rect 38180 -5440 38500 -5430
rect 38180 -5510 38190 -5440
rect 38260 -5510 38280 -5440
rect 38350 -5510 38370 -5440
rect 38440 -5510 38500 -5440
rect 38180 -5520 38500 -5510
rect 38180 -5530 38230 -5520
rect 38180 -5600 38190 -5530
rect 38180 -5620 38230 -5600
rect 38180 -5690 38190 -5620
rect 38180 -5710 38230 -5690
rect 38180 -5780 38190 -5710
rect 38470 -5760 38500 -5520
rect 38260 -5780 38280 -5760
rect 38350 -5780 38370 -5760
rect 38440 -5780 38500 -5760
rect 38180 -5800 38500 -5780
rect 38180 -5870 38190 -5800
rect 38260 -5850 38280 -5800
rect 38350 -5850 38370 -5800
rect 38440 -5850 38500 -5800
rect 38180 -5890 38230 -5870
rect 38180 -5960 38190 -5890
rect 38180 -5980 38230 -5960
rect 38180 -6050 38190 -5980
rect 38180 -6070 38230 -6050
rect 38180 -6140 38190 -6070
rect 38470 -6090 38500 -5850
rect 38260 -6140 38280 -6090
rect 38350 -6140 38370 -6090
rect 38440 -6140 38500 -6090
rect 38180 -6160 38500 -6140
rect 38180 -6230 38190 -6160
rect 38260 -6180 38280 -6160
rect 38350 -6180 38370 -6160
rect 38440 -6180 38500 -6160
rect 38180 -6250 38230 -6230
rect 38180 -6320 38190 -6250
rect 38180 -6340 38230 -6320
rect 38180 -6410 38190 -6340
rect 38180 -6420 38230 -6410
rect 38470 -6420 38500 -6180
rect 38180 -6450 38500 -6420
rect 30680 -10520 31010 -10510
rect 30680 -10590 30700 -10520
rect 30770 -10590 31010 -10520
rect 30680 -10630 31010 -10590
rect 30680 -10700 30700 -10630
rect 30770 -10700 31010 -10630
rect 30680 -10740 31010 -10700
rect 30680 -10810 30700 -10740
rect 30770 -10810 31010 -10740
rect 30680 -10830 31010 -10810
rect 27015 -11105 30477 -10995
rect 27015 -11600 27125 -11105
rect 26680 -11710 27160 -11600
rect 2210 -12240 3810 -12220
rect 2210 -12300 2390 -12240
rect 2630 -12300 2720 -12240
rect 2960 -12300 3060 -12240
rect 3300 -12300 3390 -12240
rect 3630 -12300 3810 -12240
rect 2210 -12370 2240 -12300
rect 2310 -12370 2350 -12300
rect 2640 -12370 2680 -12300
rect 2970 -12370 3010 -12300
rect 3300 -12370 3340 -12300
rect 3630 -12370 3670 -12300
rect 3740 -12370 3810 -12300
rect 2210 -12410 2390 -12370
rect 2630 -12410 2720 -12370
rect 2960 -12410 3060 -12370
rect 3300 -12410 3390 -12370
rect 3630 -12410 3810 -12370
rect 2210 -12480 2240 -12410
rect 2310 -12480 2350 -12410
rect 2640 -12480 2680 -12410
rect 2970 -12480 3010 -12410
rect 3300 -12480 3340 -12410
rect 3630 -12480 3670 -12410
rect 3740 -12480 3810 -12410
rect 2210 -12510 3810 -12480
rect 11090 -12240 12690 -12220
rect 11090 -12300 11270 -12240
rect 11510 -12300 11600 -12240
rect 11840 -12300 11940 -12240
rect 12180 -12300 12270 -12240
rect 12510 -12300 12690 -12240
rect 11090 -12370 11120 -12300
rect 11190 -12370 11230 -12300
rect 11520 -12370 11560 -12300
rect 11850 -12370 11890 -12300
rect 12180 -12370 12220 -12300
rect 12510 -12370 12550 -12300
rect 12620 -12370 12690 -12300
rect 11090 -12410 11270 -12370
rect 11510 -12410 11600 -12370
rect 11840 -12410 11940 -12370
rect 12180 -12410 12270 -12370
rect 12510 -12410 12690 -12370
rect 11090 -12480 11120 -12410
rect 11190 -12480 11230 -12410
rect 11520 -12480 11560 -12410
rect 11850 -12480 11890 -12410
rect 12180 -12480 12220 -12410
rect 12510 -12480 12550 -12410
rect 12620 -12480 12690 -12410
rect 11090 -12510 12690 -12480
rect 21610 -14020 21930 -13990
rect 21610 -14090 21630 -14020
rect 21700 -14030 21730 -14020
rect 21800 -14030 21830 -14020
rect 21900 -14090 21930 -14020
rect 21610 -14120 21650 -14090
rect 21890 -14120 21930 -14090
rect 21610 -14190 21630 -14120
rect 21900 -14190 21930 -14120
rect 21610 -14220 21650 -14190
rect 21890 -14220 21930 -14190
rect 21610 -14290 21630 -14220
rect 21700 -14290 21730 -14270
rect 21800 -14290 21830 -14270
rect 21900 -14290 21930 -14220
rect 21610 -14310 21930 -14290
rect 22900 -14870 23220 -14840
rect 22900 -14940 22920 -14870
rect 22990 -14940 23020 -14870
rect 23090 -14940 23120 -14870
rect 23190 -14940 23220 -14870
rect 22900 -14970 23220 -14940
rect 22900 -15040 22920 -14970
rect 22990 -15040 23020 -14970
rect 23090 -15040 23120 -14970
rect 23190 -15040 23220 -14970
rect 22900 -15070 23220 -15040
rect 22900 -15140 22920 -15070
rect 22990 -15140 23020 -15070
rect 23090 -15140 23120 -15070
rect 23190 -15140 23220 -15070
rect 22900 -16370 23220 -15140
rect 22900 -16690 30930 -16370
rect 7210 -17600 7650 -17580
rect 7210 -17670 7230 -17600
rect 7300 -17670 7340 -17600
rect 7410 -17670 7450 -17600
rect 7520 -17670 7560 -17600
rect 7630 -17670 7650 -17600
rect 7210 -17680 7650 -17670
rect 26480 -17620 26960 -17500
rect 26480 -17680 26600 -17620
rect 7210 -17710 26600 -17680
rect 7210 -17780 7230 -17710
rect 7300 -17780 7340 -17710
rect 7410 -17780 7450 -17710
rect 7520 -17780 7560 -17710
rect 7630 -17780 26600 -17710
rect 7210 -17800 26600 -17780
rect 7210 -17820 7650 -17800
rect 7210 -17890 7230 -17820
rect 7300 -17890 7340 -17820
rect 7410 -17890 7450 -17820
rect 7520 -17890 7560 -17820
rect 7630 -17890 7650 -17820
rect 7210 -17930 7650 -17890
rect 7210 -18000 7230 -17930
rect 7300 -18000 7340 -17930
rect 7410 -18000 7450 -17930
rect 7520 -18000 7560 -17930
rect 7630 -18000 7650 -17930
rect 7210 -18020 7650 -18000
rect 21610 -20100 21930 -20070
rect 21610 -20170 21630 -20100
rect 21700 -20110 21730 -20100
rect 21800 -20110 21830 -20100
rect 21900 -20170 21930 -20100
rect 21610 -20200 21650 -20170
rect 21890 -20200 21930 -20170
rect 21610 -20270 21630 -20200
rect 21900 -20270 21930 -20200
rect 21610 -20300 21650 -20270
rect 21890 -20300 21930 -20270
rect 21610 -20370 21630 -20300
rect 21700 -20370 21730 -20350
rect 21800 -20370 21830 -20350
rect 21900 -20370 21930 -20300
rect 21610 -20390 21930 -20370
rect 22680 -20730 23000 -20700
rect 22680 -20800 22700 -20730
rect 22770 -20800 22800 -20730
rect 22870 -20800 22900 -20730
rect 22970 -20800 23000 -20730
rect 22680 -20830 23000 -20800
rect 22680 -20900 22700 -20830
rect 22770 -20900 22800 -20830
rect 22870 -20900 22900 -20830
rect 22970 -20900 23000 -20830
rect 22680 -20930 23000 -20900
rect 22680 -21000 22700 -20930
rect 22770 -21000 22800 -20930
rect 22870 -21000 22900 -20930
rect 22970 -21000 23000 -20930
rect 22680 -22230 23000 -21000
rect 22680 -22550 30710 -22230
rect 2210 -22660 3810 -22630
rect 2210 -22730 2280 -22660
rect 2350 -22730 2390 -22660
rect 2680 -22730 2720 -22660
rect 3010 -22730 3050 -22660
rect 3340 -22730 3380 -22660
rect 3670 -22730 3710 -22660
rect 3780 -22730 3810 -22660
rect 2210 -22770 2390 -22730
rect 2630 -22770 2720 -22730
rect 2960 -22770 3060 -22730
rect 3300 -22770 3390 -22730
rect 3630 -22770 3810 -22730
rect 2210 -22840 2280 -22770
rect 2350 -22840 2390 -22770
rect 2680 -22840 2720 -22770
rect 3010 -22840 3050 -22770
rect 3340 -22840 3380 -22770
rect 3670 -22840 3710 -22770
rect 3780 -22840 3810 -22770
rect 2210 -22900 2390 -22840
rect 2630 -22900 2720 -22840
rect 2960 -22900 3060 -22840
rect 3300 -22900 3390 -22840
rect 3630 -22900 3810 -22840
rect 2210 -22910 3810 -22900
rect 11090 -22660 12690 -22630
rect 11090 -22730 11160 -22660
rect 11230 -22730 11270 -22660
rect 11560 -22730 11600 -22660
rect 11890 -22730 11930 -22660
rect 12220 -22730 12260 -22660
rect 12550 -22730 12590 -22660
rect 12660 -22730 12690 -22660
rect 11090 -22770 11270 -22730
rect 11510 -22770 11600 -22730
rect 11840 -22770 11940 -22730
rect 12180 -22770 12270 -22730
rect 12510 -22770 12690 -22730
rect 11090 -22840 11160 -22770
rect 11230 -22840 11270 -22770
rect 11560 -22840 11600 -22770
rect 11890 -22840 11930 -22770
rect 12220 -22840 12260 -22770
rect 12550 -22840 12590 -22770
rect 12660 -22840 12690 -22770
rect 11090 -22900 11270 -22840
rect 11510 -22900 11600 -22840
rect 11840 -22900 11940 -22840
rect 12180 -22900 12270 -22840
rect 12510 -22900 12690 -22840
rect 11090 -22910 12690 -22900
<< via4 >>
rect -4650 21580 -4410 21610
rect -4320 21580 -4080 21610
rect -3990 21580 -3750 21610
rect -3660 21580 -3420 21610
rect -3330 21580 -3090 21610
rect -3000 21580 -2760 21610
rect -2670 21580 -2430 21610
rect -2340 21580 -2100 21610
rect -2010 21580 -1770 21610
rect -1640 21580 -1400 21610
rect -1310 21580 -1070 21610
rect -980 21580 -740 21610
rect -650 21580 -410 21610
rect -320 21580 -80 21610
rect 10 21580 250 21610
rect 340 21580 580 21610
rect 670 21580 910 21610
rect 1000 21580 1240 21610
rect 1370 21580 1610 21610
rect 1700 21580 1940 21610
rect 2030 21580 2270 21610
rect 2360 21580 2600 21610
rect 2690 21580 2930 21610
rect 3020 21580 3260 21610
rect 3350 21580 3590 21610
rect 3680 21580 3920 21610
rect 4010 21580 4250 21610
rect 4380 21580 4620 21610
rect 4710 21580 4950 21610
rect 5040 21580 5280 21610
rect 5370 21580 5610 21610
rect 5700 21580 5940 21610
rect 6030 21580 6270 21610
rect 6360 21580 6600 21610
rect 6690 21580 6930 21610
rect 7020 21580 7260 21610
rect -4650 21510 -4640 21580
rect -4640 21510 -4570 21580
rect -4570 21510 -4550 21580
rect -4550 21510 -4480 21580
rect -4480 21510 -4460 21580
rect -4460 21510 -4410 21580
rect -4320 21510 -4300 21580
rect -4300 21510 -4280 21580
rect -4280 21510 -4210 21580
rect -4210 21510 -4190 21580
rect -4190 21510 -4120 21580
rect -4120 21510 -4100 21580
rect -4100 21510 -4080 21580
rect -3990 21510 -3940 21580
rect -3940 21510 -3920 21580
rect -3920 21510 -3850 21580
rect -3850 21510 -3830 21580
rect -3830 21510 -3760 21580
rect -3760 21510 -3750 21580
rect -3660 21510 -3650 21580
rect -3650 21510 -3580 21580
rect -3580 21510 -3560 21580
rect -3560 21510 -3490 21580
rect -3490 21510 -3470 21580
rect -3470 21510 -3420 21580
rect -3330 21510 -3310 21580
rect -3310 21510 -3290 21580
rect -3290 21510 -3220 21580
rect -3220 21510 -3200 21580
rect -3200 21510 -3130 21580
rect -3130 21510 -3110 21580
rect -3110 21510 -3090 21580
rect -3000 21510 -2950 21580
rect -2950 21510 -2930 21580
rect -2930 21510 -2860 21580
rect -2860 21510 -2840 21580
rect -2840 21510 -2770 21580
rect -2770 21510 -2760 21580
rect -2670 21510 -2660 21580
rect -2660 21510 -2590 21580
rect -2590 21510 -2570 21580
rect -2570 21510 -2500 21580
rect -2500 21510 -2480 21580
rect -2480 21510 -2430 21580
rect -2340 21510 -2320 21580
rect -2320 21510 -2300 21580
rect -2300 21510 -2230 21580
rect -2230 21510 -2210 21580
rect -2210 21510 -2140 21580
rect -2140 21510 -2120 21580
rect -2120 21510 -2100 21580
rect -2010 21510 -1960 21580
rect -1960 21510 -1940 21580
rect -1940 21510 -1870 21580
rect -1870 21510 -1850 21580
rect -1850 21510 -1780 21580
rect -1780 21510 -1770 21580
rect -1640 21510 -1630 21580
rect -1630 21510 -1560 21580
rect -1560 21510 -1540 21580
rect -1540 21510 -1470 21580
rect -1470 21510 -1450 21580
rect -1450 21510 -1400 21580
rect -1310 21510 -1290 21580
rect -1290 21510 -1270 21580
rect -1270 21510 -1200 21580
rect -1200 21510 -1180 21580
rect -1180 21510 -1110 21580
rect -1110 21510 -1090 21580
rect -1090 21510 -1070 21580
rect -980 21510 -930 21580
rect -930 21510 -910 21580
rect -910 21510 -840 21580
rect -840 21510 -820 21580
rect -820 21510 -750 21580
rect -750 21510 -740 21580
rect -650 21510 -640 21580
rect -640 21510 -570 21580
rect -570 21510 -550 21580
rect -550 21510 -480 21580
rect -480 21510 -460 21580
rect -460 21510 -410 21580
rect -320 21510 -300 21580
rect -300 21510 -280 21580
rect -280 21510 -210 21580
rect -210 21510 -190 21580
rect -190 21510 -120 21580
rect -120 21510 -100 21580
rect -100 21510 -80 21580
rect 10 21510 60 21580
rect 60 21510 80 21580
rect 80 21510 150 21580
rect 150 21510 170 21580
rect 170 21510 240 21580
rect 240 21510 250 21580
rect 340 21510 350 21580
rect 350 21510 420 21580
rect 420 21510 440 21580
rect 440 21510 510 21580
rect 510 21510 530 21580
rect 530 21510 580 21580
rect 670 21510 690 21580
rect 690 21510 710 21580
rect 710 21510 780 21580
rect 780 21510 800 21580
rect 800 21510 870 21580
rect 870 21510 890 21580
rect 890 21510 910 21580
rect 1000 21510 1050 21580
rect 1050 21510 1070 21580
rect 1070 21510 1140 21580
rect 1140 21510 1160 21580
rect 1160 21510 1230 21580
rect 1230 21510 1240 21580
rect 1370 21510 1380 21580
rect 1380 21510 1450 21580
rect 1450 21510 1470 21580
rect 1470 21510 1540 21580
rect 1540 21510 1560 21580
rect 1560 21510 1610 21580
rect 1700 21510 1720 21580
rect 1720 21510 1740 21580
rect 1740 21510 1810 21580
rect 1810 21510 1830 21580
rect 1830 21510 1900 21580
rect 1900 21510 1920 21580
rect 1920 21510 1940 21580
rect 2030 21510 2080 21580
rect 2080 21510 2100 21580
rect 2100 21510 2170 21580
rect 2170 21510 2190 21580
rect 2190 21510 2260 21580
rect 2260 21510 2270 21580
rect 2360 21510 2370 21580
rect 2370 21510 2440 21580
rect 2440 21510 2460 21580
rect 2460 21510 2530 21580
rect 2530 21510 2550 21580
rect 2550 21510 2600 21580
rect 2690 21510 2710 21580
rect 2710 21510 2730 21580
rect 2730 21510 2800 21580
rect 2800 21510 2820 21580
rect 2820 21510 2890 21580
rect 2890 21510 2910 21580
rect 2910 21510 2930 21580
rect 3020 21510 3070 21580
rect 3070 21510 3090 21580
rect 3090 21510 3160 21580
rect 3160 21510 3180 21580
rect 3180 21510 3250 21580
rect 3250 21510 3260 21580
rect 3350 21510 3360 21580
rect 3360 21510 3430 21580
rect 3430 21510 3450 21580
rect 3450 21510 3520 21580
rect 3520 21510 3540 21580
rect 3540 21510 3590 21580
rect 3680 21510 3700 21580
rect 3700 21510 3720 21580
rect 3720 21510 3790 21580
rect 3790 21510 3810 21580
rect 3810 21510 3880 21580
rect 3880 21510 3900 21580
rect 3900 21510 3920 21580
rect 4010 21510 4060 21580
rect 4060 21510 4080 21580
rect 4080 21510 4150 21580
rect 4150 21510 4170 21580
rect 4170 21510 4240 21580
rect 4240 21510 4250 21580
rect 4380 21510 4390 21580
rect 4390 21510 4460 21580
rect 4460 21510 4480 21580
rect 4480 21510 4550 21580
rect 4550 21510 4570 21580
rect 4570 21510 4620 21580
rect 4710 21510 4730 21580
rect 4730 21510 4750 21580
rect 4750 21510 4820 21580
rect 4820 21510 4840 21580
rect 4840 21510 4910 21580
rect 4910 21510 4930 21580
rect 4930 21510 4950 21580
rect 5040 21510 5090 21580
rect 5090 21510 5110 21580
rect 5110 21510 5180 21580
rect 5180 21510 5200 21580
rect 5200 21510 5270 21580
rect 5270 21510 5280 21580
rect 5370 21510 5380 21580
rect 5380 21510 5450 21580
rect 5450 21510 5470 21580
rect 5470 21510 5540 21580
rect 5540 21510 5560 21580
rect 5560 21510 5610 21580
rect 5700 21510 5720 21580
rect 5720 21510 5740 21580
rect 5740 21510 5810 21580
rect 5810 21510 5830 21580
rect 5830 21510 5900 21580
rect 5900 21510 5920 21580
rect 5920 21510 5940 21580
rect 6030 21510 6080 21580
rect 6080 21510 6100 21580
rect 6100 21510 6170 21580
rect 6170 21510 6190 21580
rect 6190 21510 6260 21580
rect 6260 21510 6270 21580
rect 6360 21510 6370 21580
rect 6370 21510 6440 21580
rect 6440 21510 6460 21580
rect 6460 21510 6530 21580
rect 6530 21510 6550 21580
rect 6550 21510 6600 21580
rect 6690 21510 6710 21580
rect 6710 21510 6730 21580
rect 6730 21510 6800 21580
rect 6800 21510 6820 21580
rect 6820 21510 6890 21580
rect 6890 21510 6910 21580
rect 6910 21510 6930 21580
rect 7020 21510 7070 21580
rect 7070 21510 7090 21580
rect 7090 21510 7160 21580
rect 7160 21510 7180 21580
rect 7180 21510 7250 21580
rect 7250 21510 7260 21580
rect -4650 21490 -4410 21510
rect -4320 21490 -4080 21510
rect -3990 21490 -3750 21510
rect -3660 21490 -3420 21510
rect -3330 21490 -3090 21510
rect -3000 21490 -2760 21510
rect -2670 21490 -2430 21510
rect -2340 21490 -2100 21510
rect -2010 21490 -1770 21510
rect -1640 21490 -1400 21510
rect -1310 21490 -1070 21510
rect -980 21490 -740 21510
rect -650 21490 -410 21510
rect -320 21490 -80 21510
rect 10 21490 250 21510
rect 340 21490 580 21510
rect 670 21490 910 21510
rect 1000 21490 1240 21510
rect 1370 21490 1610 21510
rect 1700 21490 1940 21510
rect 2030 21490 2270 21510
rect 2360 21490 2600 21510
rect 2690 21490 2930 21510
rect 3020 21490 3260 21510
rect 3350 21490 3590 21510
rect 3680 21490 3920 21510
rect 4010 21490 4250 21510
rect 4380 21490 4620 21510
rect 4710 21490 4950 21510
rect 5040 21490 5280 21510
rect 5370 21490 5610 21510
rect 5700 21490 5940 21510
rect 6030 21490 6270 21510
rect 6360 21490 6600 21510
rect 6690 21490 6930 21510
rect 7020 21490 7260 21510
rect -4650 21420 -4640 21490
rect -4640 21420 -4570 21490
rect -4570 21420 -4550 21490
rect -4550 21420 -4480 21490
rect -4480 21420 -4460 21490
rect -4460 21420 -4410 21490
rect -4320 21420 -4300 21490
rect -4300 21420 -4280 21490
rect -4280 21420 -4210 21490
rect -4210 21420 -4190 21490
rect -4190 21420 -4120 21490
rect -4120 21420 -4100 21490
rect -4100 21420 -4080 21490
rect -3990 21420 -3940 21490
rect -3940 21420 -3920 21490
rect -3920 21420 -3850 21490
rect -3850 21420 -3830 21490
rect -3830 21420 -3760 21490
rect -3760 21420 -3750 21490
rect -3660 21420 -3650 21490
rect -3650 21420 -3580 21490
rect -3580 21420 -3560 21490
rect -3560 21420 -3490 21490
rect -3490 21420 -3470 21490
rect -3470 21420 -3420 21490
rect -3330 21420 -3310 21490
rect -3310 21420 -3290 21490
rect -3290 21420 -3220 21490
rect -3220 21420 -3200 21490
rect -3200 21420 -3130 21490
rect -3130 21420 -3110 21490
rect -3110 21420 -3090 21490
rect -3000 21420 -2950 21490
rect -2950 21420 -2930 21490
rect -2930 21420 -2860 21490
rect -2860 21420 -2840 21490
rect -2840 21420 -2770 21490
rect -2770 21420 -2760 21490
rect -2670 21420 -2660 21490
rect -2660 21420 -2590 21490
rect -2590 21420 -2570 21490
rect -2570 21420 -2500 21490
rect -2500 21420 -2480 21490
rect -2480 21420 -2430 21490
rect -2340 21420 -2320 21490
rect -2320 21420 -2300 21490
rect -2300 21420 -2230 21490
rect -2230 21420 -2210 21490
rect -2210 21420 -2140 21490
rect -2140 21420 -2120 21490
rect -2120 21420 -2100 21490
rect -2010 21420 -1960 21490
rect -1960 21420 -1940 21490
rect -1940 21420 -1870 21490
rect -1870 21420 -1850 21490
rect -1850 21420 -1780 21490
rect -1780 21420 -1770 21490
rect -1640 21420 -1630 21490
rect -1630 21420 -1560 21490
rect -1560 21420 -1540 21490
rect -1540 21420 -1470 21490
rect -1470 21420 -1450 21490
rect -1450 21420 -1400 21490
rect -1310 21420 -1290 21490
rect -1290 21420 -1270 21490
rect -1270 21420 -1200 21490
rect -1200 21420 -1180 21490
rect -1180 21420 -1110 21490
rect -1110 21420 -1090 21490
rect -1090 21420 -1070 21490
rect -980 21420 -930 21490
rect -930 21420 -910 21490
rect -910 21420 -840 21490
rect -840 21420 -820 21490
rect -820 21420 -750 21490
rect -750 21420 -740 21490
rect -650 21420 -640 21490
rect -640 21420 -570 21490
rect -570 21420 -550 21490
rect -550 21420 -480 21490
rect -480 21420 -460 21490
rect -460 21420 -410 21490
rect -320 21420 -300 21490
rect -300 21420 -280 21490
rect -280 21420 -210 21490
rect -210 21420 -190 21490
rect -190 21420 -120 21490
rect -120 21420 -100 21490
rect -100 21420 -80 21490
rect 10 21420 60 21490
rect 60 21420 80 21490
rect 80 21420 150 21490
rect 150 21420 170 21490
rect 170 21420 240 21490
rect 240 21420 250 21490
rect 340 21420 350 21490
rect 350 21420 420 21490
rect 420 21420 440 21490
rect 440 21420 510 21490
rect 510 21420 530 21490
rect 530 21420 580 21490
rect 670 21420 690 21490
rect 690 21420 710 21490
rect 710 21420 780 21490
rect 780 21420 800 21490
rect 800 21420 870 21490
rect 870 21420 890 21490
rect 890 21420 910 21490
rect 1000 21420 1050 21490
rect 1050 21420 1070 21490
rect 1070 21420 1140 21490
rect 1140 21420 1160 21490
rect 1160 21420 1230 21490
rect 1230 21420 1240 21490
rect 1370 21420 1380 21490
rect 1380 21420 1450 21490
rect 1450 21420 1470 21490
rect 1470 21420 1540 21490
rect 1540 21420 1560 21490
rect 1560 21420 1610 21490
rect 1700 21420 1720 21490
rect 1720 21420 1740 21490
rect 1740 21420 1810 21490
rect 1810 21420 1830 21490
rect 1830 21420 1900 21490
rect 1900 21420 1920 21490
rect 1920 21420 1940 21490
rect 2030 21420 2080 21490
rect 2080 21420 2100 21490
rect 2100 21420 2170 21490
rect 2170 21420 2190 21490
rect 2190 21420 2260 21490
rect 2260 21420 2270 21490
rect 2360 21420 2370 21490
rect 2370 21420 2440 21490
rect 2440 21420 2460 21490
rect 2460 21420 2530 21490
rect 2530 21420 2550 21490
rect 2550 21420 2600 21490
rect 2690 21420 2710 21490
rect 2710 21420 2730 21490
rect 2730 21420 2800 21490
rect 2800 21420 2820 21490
rect 2820 21420 2890 21490
rect 2890 21420 2910 21490
rect 2910 21420 2930 21490
rect 3020 21420 3070 21490
rect 3070 21420 3090 21490
rect 3090 21420 3160 21490
rect 3160 21420 3180 21490
rect 3180 21420 3250 21490
rect 3250 21420 3260 21490
rect 3350 21420 3360 21490
rect 3360 21420 3430 21490
rect 3430 21420 3450 21490
rect 3450 21420 3520 21490
rect 3520 21420 3540 21490
rect 3540 21420 3590 21490
rect 3680 21420 3700 21490
rect 3700 21420 3720 21490
rect 3720 21420 3790 21490
rect 3790 21420 3810 21490
rect 3810 21420 3880 21490
rect 3880 21420 3900 21490
rect 3900 21420 3920 21490
rect 4010 21420 4060 21490
rect 4060 21420 4080 21490
rect 4080 21420 4150 21490
rect 4150 21420 4170 21490
rect 4170 21420 4240 21490
rect 4240 21420 4250 21490
rect 4380 21420 4390 21490
rect 4390 21420 4460 21490
rect 4460 21420 4480 21490
rect 4480 21420 4550 21490
rect 4550 21420 4570 21490
rect 4570 21420 4620 21490
rect 4710 21420 4730 21490
rect 4730 21420 4750 21490
rect 4750 21420 4820 21490
rect 4820 21420 4840 21490
rect 4840 21420 4910 21490
rect 4910 21420 4930 21490
rect 4930 21420 4950 21490
rect 5040 21420 5090 21490
rect 5090 21420 5110 21490
rect 5110 21420 5180 21490
rect 5180 21420 5200 21490
rect 5200 21420 5270 21490
rect 5270 21420 5280 21490
rect 5370 21420 5380 21490
rect 5380 21420 5450 21490
rect 5450 21420 5470 21490
rect 5470 21420 5540 21490
rect 5540 21420 5560 21490
rect 5560 21420 5610 21490
rect 5700 21420 5720 21490
rect 5720 21420 5740 21490
rect 5740 21420 5810 21490
rect 5810 21420 5830 21490
rect 5830 21420 5900 21490
rect 5900 21420 5920 21490
rect 5920 21420 5940 21490
rect 6030 21420 6080 21490
rect 6080 21420 6100 21490
rect 6100 21420 6170 21490
rect 6170 21420 6190 21490
rect 6190 21420 6260 21490
rect 6260 21420 6270 21490
rect 6360 21420 6370 21490
rect 6370 21420 6440 21490
rect 6440 21420 6460 21490
rect 6460 21420 6530 21490
rect 6530 21420 6550 21490
rect 6550 21420 6600 21490
rect 6690 21420 6710 21490
rect 6710 21420 6730 21490
rect 6730 21420 6800 21490
rect 6800 21420 6820 21490
rect 6820 21420 6890 21490
rect 6890 21420 6910 21490
rect 6910 21420 6930 21490
rect 7020 21420 7070 21490
rect 7070 21420 7090 21490
rect 7090 21420 7160 21490
rect 7160 21420 7180 21490
rect 7180 21420 7250 21490
rect 7250 21420 7260 21490
rect -4650 21400 -4410 21420
rect -4320 21400 -4080 21420
rect -3990 21400 -3750 21420
rect -3660 21400 -3420 21420
rect -3330 21400 -3090 21420
rect -3000 21400 -2760 21420
rect -2670 21400 -2430 21420
rect -2340 21400 -2100 21420
rect -2010 21400 -1770 21420
rect -1640 21400 -1400 21420
rect -1310 21400 -1070 21420
rect -980 21400 -740 21420
rect -650 21400 -410 21420
rect -320 21400 -80 21420
rect 10 21400 250 21420
rect 340 21400 580 21420
rect 670 21400 910 21420
rect 1000 21400 1240 21420
rect 1370 21400 1610 21420
rect 1700 21400 1940 21420
rect 2030 21400 2270 21420
rect 2360 21400 2600 21420
rect 2690 21400 2930 21420
rect 3020 21400 3260 21420
rect 3350 21400 3590 21420
rect 3680 21400 3920 21420
rect 4010 21400 4250 21420
rect 4380 21400 4620 21420
rect 4710 21400 4950 21420
rect 5040 21400 5280 21420
rect 5370 21400 5610 21420
rect 5700 21400 5940 21420
rect 6030 21400 6270 21420
rect 6360 21400 6600 21420
rect 6690 21400 6930 21420
rect 7020 21400 7260 21420
rect -4650 21370 -4640 21400
rect -4640 21370 -4570 21400
rect -4570 21370 -4550 21400
rect -4550 21370 -4480 21400
rect -4480 21370 -4460 21400
rect -4460 21370 -4410 21400
rect -4320 21370 -4300 21400
rect -4300 21370 -4280 21400
rect -4280 21370 -4210 21400
rect -4210 21370 -4190 21400
rect -4190 21370 -4120 21400
rect -4120 21370 -4100 21400
rect -4100 21370 -4080 21400
rect -3990 21370 -3940 21400
rect -3940 21370 -3920 21400
rect -3920 21370 -3850 21400
rect -3850 21370 -3830 21400
rect -3830 21370 -3760 21400
rect -3760 21370 -3750 21400
rect -3660 21370 -3650 21400
rect -3650 21370 -3580 21400
rect -3580 21370 -3560 21400
rect -3560 21370 -3490 21400
rect -3490 21370 -3470 21400
rect -3470 21370 -3420 21400
rect -3330 21370 -3310 21400
rect -3310 21370 -3290 21400
rect -3290 21370 -3220 21400
rect -3220 21370 -3200 21400
rect -3200 21370 -3130 21400
rect -3130 21370 -3110 21400
rect -3110 21370 -3090 21400
rect -3000 21370 -2950 21400
rect -2950 21370 -2930 21400
rect -2930 21370 -2860 21400
rect -2860 21370 -2840 21400
rect -2840 21370 -2770 21400
rect -2770 21370 -2760 21400
rect -2670 21370 -2660 21400
rect -2660 21370 -2590 21400
rect -2590 21370 -2570 21400
rect -2570 21370 -2500 21400
rect -2500 21370 -2480 21400
rect -2480 21370 -2430 21400
rect -2340 21370 -2320 21400
rect -2320 21370 -2300 21400
rect -2300 21370 -2230 21400
rect -2230 21370 -2210 21400
rect -2210 21370 -2140 21400
rect -2140 21370 -2120 21400
rect -2120 21370 -2100 21400
rect -2010 21370 -1960 21400
rect -1960 21370 -1940 21400
rect -1940 21370 -1870 21400
rect -1870 21370 -1850 21400
rect -1850 21370 -1780 21400
rect -1780 21370 -1770 21400
rect -1640 21370 -1630 21400
rect -1630 21370 -1560 21400
rect -1560 21370 -1540 21400
rect -1540 21370 -1470 21400
rect -1470 21370 -1450 21400
rect -1450 21370 -1400 21400
rect -1310 21370 -1290 21400
rect -1290 21370 -1270 21400
rect -1270 21370 -1200 21400
rect -1200 21370 -1180 21400
rect -1180 21370 -1110 21400
rect -1110 21370 -1090 21400
rect -1090 21370 -1070 21400
rect -980 21370 -930 21400
rect -930 21370 -910 21400
rect -910 21370 -840 21400
rect -840 21370 -820 21400
rect -820 21370 -750 21400
rect -750 21370 -740 21400
rect -650 21370 -640 21400
rect -640 21370 -570 21400
rect -570 21370 -550 21400
rect -550 21370 -480 21400
rect -480 21370 -460 21400
rect -460 21370 -410 21400
rect -320 21370 -300 21400
rect -300 21370 -280 21400
rect -280 21370 -210 21400
rect -210 21370 -190 21400
rect -190 21370 -120 21400
rect -120 21370 -100 21400
rect -100 21370 -80 21400
rect 10 21370 60 21400
rect 60 21370 80 21400
rect 80 21370 150 21400
rect 150 21370 170 21400
rect 170 21370 240 21400
rect 240 21370 250 21400
rect 340 21370 350 21400
rect 350 21370 420 21400
rect 420 21370 440 21400
rect 440 21370 510 21400
rect 510 21370 530 21400
rect 530 21370 580 21400
rect 670 21370 690 21400
rect 690 21370 710 21400
rect 710 21370 780 21400
rect 780 21370 800 21400
rect 800 21370 870 21400
rect 870 21370 890 21400
rect 890 21370 910 21400
rect 1000 21370 1050 21400
rect 1050 21370 1070 21400
rect 1070 21370 1140 21400
rect 1140 21370 1160 21400
rect 1160 21370 1230 21400
rect 1230 21370 1240 21400
rect 1370 21370 1380 21400
rect 1380 21370 1450 21400
rect 1450 21370 1470 21400
rect 1470 21370 1540 21400
rect 1540 21370 1560 21400
rect 1560 21370 1610 21400
rect 1700 21370 1720 21400
rect 1720 21370 1740 21400
rect 1740 21370 1810 21400
rect 1810 21370 1830 21400
rect 1830 21370 1900 21400
rect 1900 21370 1920 21400
rect 1920 21370 1940 21400
rect 2030 21370 2080 21400
rect 2080 21370 2100 21400
rect 2100 21370 2170 21400
rect 2170 21370 2190 21400
rect 2190 21370 2260 21400
rect 2260 21370 2270 21400
rect 2360 21370 2370 21400
rect 2370 21370 2440 21400
rect 2440 21370 2460 21400
rect 2460 21370 2530 21400
rect 2530 21370 2550 21400
rect 2550 21370 2600 21400
rect 2690 21370 2710 21400
rect 2710 21370 2730 21400
rect 2730 21370 2800 21400
rect 2800 21370 2820 21400
rect 2820 21370 2890 21400
rect 2890 21370 2910 21400
rect 2910 21370 2930 21400
rect 3020 21370 3070 21400
rect 3070 21370 3090 21400
rect 3090 21370 3160 21400
rect 3160 21370 3180 21400
rect 3180 21370 3250 21400
rect 3250 21370 3260 21400
rect 3350 21370 3360 21400
rect 3360 21370 3430 21400
rect 3430 21370 3450 21400
rect 3450 21370 3520 21400
rect 3520 21370 3540 21400
rect 3540 21370 3590 21400
rect 3680 21370 3700 21400
rect 3700 21370 3720 21400
rect 3720 21370 3790 21400
rect 3790 21370 3810 21400
rect 3810 21370 3880 21400
rect 3880 21370 3900 21400
rect 3900 21370 3920 21400
rect 4010 21370 4060 21400
rect 4060 21370 4080 21400
rect 4080 21370 4150 21400
rect 4150 21370 4170 21400
rect 4170 21370 4240 21400
rect 4240 21370 4250 21400
rect 4380 21370 4390 21400
rect 4390 21370 4460 21400
rect 4460 21370 4480 21400
rect 4480 21370 4550 21400
rect 4550 21370 4570 21400
rect 4570 21370 4620 21400
rect 4710 21370 4730 21400
rect 4730 21370 4750 21400
rect 4750 21370 4820 21400
rect 4820 21370 4840 21400
rect 4840 21370 4910 21400
rect 4910 21370 4930 21400
rect 4930 21370 4950 21400
rect 5040 21370 5090 21400
rect 5090 21370 5110 21400
rect 5110 21370 5180 21400
rect 5180 21370 5200 21400
rect 5200 21370 5270 21400
rect 5270 21370 5280 21400
rect 5370 21370 5380 21400
rect 5380 21370 5450 21400
rect 5450 21370 5470 21400
rect 5470 21370 5540 21400
rect 5540 21370 5560 21400
rect 5560 21370 5610 21400
rect 5700 21370 5720 21400
rect 5720 21370 5740 21400
rect 5740 21370 5810 21400
rect 5810 21370 5830 21400
rect 5830 21370 5900 21400
rect 5900 21370 5920 21400
rect 5920 21370 5940 21400
rect 6030 21370 6080 21400
rect 6080 21370 6100 21400
rect 6100 21370 6170 21400
rect 6170 21370 6190 21400
rect 6190 21370 6260 21400
rect 6260 21370 6270 21400
rect 6360 21370 6370 21400
rect 6370 21370 6440 21400
rect 6440 21370 6460 21400
rect 6460 21370 6530 21400
rect 6530 21370 6550 21400
rect 6550 21370 6600 21400
rect 6690 21370 6710 21400
rect 6710 21370 6730 21400
rect 6730 21370 6800 21400
rect 6800 21370 6820 21400
rect 6820 21370 6890 21400
rect 6890 21370 6910 21400
rect 6910 21370 6930 21400
rect 7020 21370 7070 21400
rect 7070 21370 7090 21400
rect 7090 21370 7160 21400
rect 7160 21370 7180 21400
rect 7180 21370 7250 21400
rect 7250 21370 7260 21400
rect 7640 21580 7880 21610
rect 7970 21580 8210 21610
rect 8300 21580 8540 21610
rect 8630 21580 8870 21610
rect 8960 21580 9200 21610
rect 9290 21580 9530 21610
rect 9620 21580 9860 21610
rect 9950 21580 10190 21610
rect 10280 21580 10520 21610
rect 10650 21580 10890 21610
rect 10980 21580 11220 21610
rect 11310 21580 11550 21610
rect 11640 21580 11880 21610
rect 11970 21580 12210 21610
rect 12300 21580 12540 21610
rect 12630 21580 12870 21610
rect 12960 21580 13200 21610
rect 13290 21580 13530 21610
rect 13660 21580 13900 21610
rect 13990 21580 14230 21610
rect 14320 21580 14560 21610
rect 14650 21580 14890 21610
rect 14980 21580 15220 21610
rect 15310 21580 15550 21610
rect 15640 21580 15880 21610
rect 15970 21580 16210 21610
rect 16300 21580 16540 21610
rect 16670 21580 16910 21610
rect 17000 21580 17240 21610
rect 17330 21580 17570 21610
rect 17660 21580 17900 21610
rect 17990 21580 18230 21610
rect 18320 21580 18560 21610
rect 18650 21580 18890 21610
rect 18980 21580 19220 21610
rect 19310 21580 19550 21610
rect 7640 21510 7650 21580
rect 7650 21510 7720 21580
rect 7720 21510 7740 21580
rect 7740 21510 7810 21580
rect 7810 21510 7830 21580
rect 7830 21510 7880 21580
rect 7970 21510 7990 21580
rect 7990 21510 8010 21580
rect 8010 21510 8080 21580
rect 8080 21510 8100 21580
rect 8100 21510 8170 21580
rect 8170 21510 8190 21580
rect 8190 21510 8210 21580
rect 8300 21510 8350 21580
rect 8350 21510 8370 21580
rect 8370 21510 8440 21580
rect 8440 21510 8460 21580
rect 8460 21510 8530 21580
rect 8530 21510 8540 21580
rect 8630 21510 8640 21580
rect 8640 21510 8710 21580
rect 8710 21510 8730 21580
rect 8730 21510 8800 21580
rect 8800 21510 8820 21580
rect 8820 21510 8870 21580
rect 8960 21510 8980 21580
rect 8980 21510 9000 21580
rect 9000 21510 9070 21580
rect 9070 21510 9090 21580
rect 9090 21510 9160 21580
rect 9160 21510 9180 21580
rect 9180 21510 9200 21580
rect 9290 21510 9340 21580
rect 9340 21510 9360 21580
rect 9360 21510 9430 21580
rect 9430 21510 9450 21580
rect 9450 21510 9520 21580
rect 9520 21510 9530 21580
rect 9620 21510 9630 21580
rect 9630 21510 9700 21580
rect 9700 21510 9720 21580
rect 9720 21510 9790 21580
rect 9790 21510 9810 21580
rect 9810 21510 9860 21580
rect 9950 21510 9970 21580
rect 9970 21510 9990 21580
rect 9990 21510 10060 21580
rect 10060 21510 10080 21580
rect 10080 21510 10150 21580
rect 10150 21510 10170 21580
rect 10170 21510 10190 21580
rect 10280 21510 10330 21580
rect 10330 21510 10350 21580
rect 10350 21510 10420 21580
rect 10420 21510 10440 21580
rect 10440 21510 10510 21580
rect 10510 21510 10520 21580
rect 10650 21510 10660 21580
rect 10660 21510 10730 21580
rect 10730 21510 10750 21580
rect 10750 21510 10820 21580
rect 10820 21510 10840 21580
rect 10840 21510 10890 21580
rect 10980 21510 11000 21580
rect 11000 21510 11020 21580
rect 11020 21510 11090 21580
rect 11090 21510 11110 21580
rect 11110 21510 11180 21580
rect 11180 21510 11200 21580
rect 11200 21510 11220 21580
rect 11310 21510 11360 21580
rect 11360 21510 11380 21580
rect 11380 21510 11450 21580
rect 11450 21510 11470 21580
rect 11470 21510 11540 21580
rect 11540 21510 11550 21580
rect 11640 21510 11650 21580
rect 11650 21510 11720 21580
rect 11720 21510 11740 21580
rect 11740 21510 11810 21580
rect 11810 21510 11830 21580
rect 11830 21510 11880 21580
rect 11970 21510 11990 21580
rect 11990 21510 12010 21580
rect 12010 21510 12080 21580
rect 12080 21510 12100 21580
rect 12100 21510 12170 21580
rect 12170 21510 12190 21580
rect 12190 21510 12210 21580
rect 12300 21510 12350 21580
rect 12350 21510 12370 21580
rect 12370 21510 12440 21580
rect 12440 21510 12460 21580
rect 12460 21510 12530 21580
rect 12530 21510 12540 21580
rect 12630 21510 12640 21580
rect 12640 21510 12710 21580
rect 12710 21510 12730 21580
rect 12730 21510 12800 21580
rect 12800 21510 12820 21580
rect 12820 21510 12870 21580
rect 12960 21510 12980 21580
rect 12980 21510 13000 21580
rect 13000 21510 13070 21580
rect 13070 21510 13090 21580
rect 13090 21510 13160 21580
rect 13160 21510 13180 21580
rect 13180 21510 13200 21580
rect 13290 21510 13340 21580
rect 13340 21510 13360 21580
rect 13360 21510 13430 21580
rect 13430 21510 13450 21580
rect 13450 21510 13520 21580
rect 13520 21510 13530 21580
rect 13660 21510 13670 21580
rect 13670 21510 13740 21580
rect 13740 21510 13760 21580
rect 13760 21510 13830 21580
rect 13830 21510 13850 21580
rect 13850 21510 13900 21580
rect 13990 21510 14010 21580
rect 14010 21510 14030 21580
rect 14030 21510 14100 21580
rect 14100 21510 14120 21580
rect 14120 21510 14190 21580
rect 14190 21510 14210 21580
rect 14210 21510 14230 21580
rect 14320 21510 14370 21580
rect 14370 21510 14390 21580
rect 14390 21510 14460 21580
rect 14460 21510 14480 21580
rect 14480 21510 14550 21580
rect 14550 21510 14560 21580
rect 14650 21510 14660 21580
rect 14660 21510 14730 21580
rect 14730 21510 14750 21580
rect 14750 21510 14820 21580
rect 14820 21510 14840 21580
rect 14840 21510 14890 21580
rect 14980 21510 15000 21580
rect 15000 21510 15020 21580
rect 15020 21510 15090 21580
rect 15090 21510 15110 21580
rect 15110 21510 15180 21580
rect 15180 21510 15200 21580
rect 15200 21510 15220 21580
rect 15310 21510 15360 21580
rect 15360 21510 15380 21580
rect 15380 21510 15450 21580
rect 15450 21510 15470 21580
rect 15470 21510 15540 21580
rect 15540 21510 15550 21580
rect 15640 21510 15650 21580
rect 15650 21510 15720 21580
rect 15720 21510 15740 21580
rect 15740 21510 15810 21580
rect 15810 21510 15830 21580
rect 15830 21510 15880 21580
rect 15970 21510 15990 21580
rect 15990 21510 16010 21580
rect 16010 21510 16080 21580
rect 16080 21510 16100 21580
rect 16100 21510 16170 21580
rect 16170 21510 16190 21580
rect 16190 21510 16210 21580
rect 16300 21510 16350 21580
rect 16350 21510 16370 21580
rect 16370 21510 16440 21580
rect 16440 21510 16460 21580
rect 16460 21510 16530 21580
rect 16530 21510 16540 21580
rect 16670 21510 16680 21580
rect 16680 21510 16750 21580
rect 16750 21510 16770 21580
rect 16770 21510 16840 21580
rect 16840 21510 16860 21580
rect 16860 21510 16910 21580
rect 17000 21510 17020 21580
rect 17020 21510 17040 21580
rect 17040 21510 17110 21580
rect 17110 21510 17130 21580
rect 17130 21510 17200 21580
rect 17200 21510 17220 21580
rect 17220 21510 17240 21580
rect 17330 21510 17380 21580
rect 17380 21510 17400 21580
rect 17400 21510 17470 21580
rect 17470 21510 17490 21580
rect 17490 21510 17560 21580
rect 17560 21510 17570 21580
rect 17660 21510 17670 21580
rect 17670 21510 17740 21580
rect 17740 21510 17760 21580
rect 17760 21510 17830 21580
rect 17830 21510 17850 21580
rect 17850 21510 17900 21580
rect 17990 21510 18010 21580
rect 18010 21510 18030 21580
rect 18030 21510 18100 21580
rect 18100 21510 18120 21580
rect 18120 21510 18190 21580
rect 18190 21510 18210 21580
rect 18210 21510 18230 21580
rect 18320 21510 18370 21580
rect 18370 21510 18390 21580
rect 18390 21510 18460 21580
rect 18460 21510 18480 21580
rect 18480 21510 18550 21580
rect 18550 21510 18560 21580
rect 18650 21510 18660 21580
rect 18660 21510 18730 21580
rect 18730 21510 18750 21580
rect 18750 21510 18820 21580
rect 18820 21510 18840 21580
rect 18840 21510 18890 21580
rect 18980 21510 19000 21580
rect 19000 21510 19020 21580
rect 19020 21510 19090 21580
rect 19090 21510 19110 21580
rect 19110 21510 19180 21580
rect 19180 21510 19200 21580
rect 19200 21510 19220 21580
rect 19310 21510 19360 21580
rect 19360 21510 19380 21580
rect 19380 21510 19450 21580
rect 19450 21510 19470 21580
rect 19470 21510 19540 21580
rect 19540 21510 19550 21580
rect 7640 21490 7880 21510
rect 7970 21490 8210 21510
rect 8300 21490 8540 21510
rect 8630 21490 8870 21510
rect 8960 21490 9200 21510
rect 9290 21490 9530 21510
rect 9620 21490 9860 21510
rect 9950 21490 10190 21510
rect 10280 21490 10520 21510
rect 10650 21490 10890 21510
rect 10980 21490 11220 21510
rect 11310 21490 11550 21510
rect 11640 21490 11880 21510
rect 11970 21490 12210 21510
rect 12300 21490 12540 21510
rect 12630 21490 12870 21510
rect 12960 21490 13200 21510
rect 13290 21490 13530 21510
rect 13660 21490 13900 21510
rect 13990 21490 14230 21510
rect 14320 21490 14560 21510
rect 14650 21490 14890 21510
rect 14980 21490 15220 21510
rect 15310 21490 15550 21510
rect 15640 21490 15880 21510
rect 15970 21490 16210 21510
rect 16300 21490 16540 21510
rect 16670 21490 16910 21510
rect 17000 21490 17240 21510
rect 17330 21490 17570 21510
rect 17660 21490 17900 21510
rect 17990 21490 18230 21510
rect 18320 21490 18560 21510
rect 18650 21490 18890 21510
rect 18980 21490 19220 21510
rect 19310 21490 19550 21510
rect 7640 21420 7650 21490
rect 7650 21420 7720 21490
rect 7720 21420 7740 21490
rect 7740 21420 7810 21490
rect 7810 21420 7830 21490
rect 7830 21420 7880 21490
rect 7970 21420 7990 21490
rect 7990 21420 8010 21490
rect 8010 21420 8080 21490
rect 8080 21420 8100 21490
rect 8100 21420 8170 21490
rect 8170 21420 8190 21490
rect 8190 21420 8210 21490
rect 8300 21420 8350 21490
rect 8350 21420 8370 21490
rect 8370 21420 8440 21490
rect 8440 21420 8460 21490
rect 8460 21420 8530 21490
rect 8530 21420 8540 21490
rect 8630 21420 8640 21490
rect 8640 21420 8710 21490
rect 8710 21420 8730 21490
rect 8730 21420 8800 21490
rect 8800 21420 8820 21490
rect 8820 21420 8870 21490
rect 8960 21420 8980 21490
rect 8980 21420 9000 21490
rect 9000 21420 9070 21490
rect 9070 21420 9090 21490
rect 9090 21420 9160 21490
rect 9160 21420 9180 21490
rect 9180 21420 9200 21490
rect 9290 21420 9340 21490
rect 9340 21420 9360 21490
rect 9360 21420 9430 21490
rect 9430 21420 9450 21490
rect 9450 21420 9520 21490
rect 9520 21420 9530 21490
rect 9620 21420 9630 21490
rect 9630 21420 9700 21490
rect 9700 21420 9720 21490
rect 9720 21420 9790 21490
rect 9790 21420 9810 21490
rect 9810 21420 9860 21490
rect 9950 21420 9970 21490
rect 9970 21420 9990 21490
rect 9990 21420 10060 21490
rect 10060 21420 10080 21490
rect 10080 21420 10150 21490
rect 10150 21420 10170 21490
rect 10170 21420 10190 21490
rect 10280 21420 10330 21490
rect 10330 21420 10350 21490
rect 10350 21420 10420 21490
rect 10420 21420 10440 21490
rect 10440 21420 10510 21490
rect 10510 21420 10520 21490
rect 10650 21420 10660 21490
rect 10660 21420 10730 21490
rect 10730 21420 10750 21490
rect 10750 21420 10820 21490
rect 10820 21420 10840 21490
rect 10840 21420 10890 21490
rect 10980 21420 11000 21490
rect 11000 21420 11020 21490
rect 11020 21420 11090 21490
rect 11090 21420 11110 21490
rect 11110 21420 11180 21490
rect 11180 21420 11200 21490
rect 11200 21420 11220 21490
rect 11310 21420 11360 21490
rect 11360 21420 11380 21490
rect 11380 21420 11450 21490
rect 11450 21420 11470 21490
rect 11470 21420 11540 21490
rect 11540 21420 11550 21490
rect 11640 21420 11650 21490
rect 11650 21420 11720 21490
rect 11720 21420 11740 21490
rect 11740 21420 11810 21490
rect 11810 21420 11830 21490
rect 11830 21420 11880 21490
rect 11970 21420 11990 21490
rect 11990 21420 12010 21490
rect 12010 21420 12080 21490
rect 12080 21420 12100 21490
rect 12100 21420 12170 21490
rect 12170 21420 12190 21490
rect 12190 21420 12210 21490
rect 12300 21420 12350 21490
rect 12350 21420 12370 21490
rect 12370 21420 12440 21490
rect 12440 21420 12460 21490
rect 12460 21420 12530 21490
rect 12530 21420 12540 21490
rect 12630 21420 12640 21490
rect 12640 21420 12710 21490
rect 12710 21420 12730 21490
rect 12730 21420 12800 21490
rect 12800 21420 12820 21490
rect 12820 21420 12870 21490
rect 12960 21420 12980 21490
rect 12980 21420 13000 21490
rect 13000 21420 13070 21490
rect 13070 21420 13090 21490
rect 13090 21420 13160 21490
rect 13160 21420 13180 21490
rect 13180 21420 13200 21490
rect 13290 21420 13340 21490
rect 13340 21420 13360 21490
rect 13360 21420 13430 21490
rect 13430 21420 13450 21490
rect 13450 21420 13520 21490
rect 13520 21420 13530 21490
rect 13660 21420 13670 21490
rect 13670 21420 13740 21490
rect 13740 21420 13760 21490
rect 13760 21420 13830 21490
rect 13830 21420 13850 21490
rect 13850 21420 13900 21490
rect 13990 21420 14010 21490
rect 14010 21420 14030 21490
rect 14030 21420 14100 21490
rect 14100 21420 14120 21490
rect 14120 21420 14190 21490
rect 14190 21420 14210 21490
rect 14210 21420 14230 21490
rect 14320 21420 14370 21490
rect 14370 21420 14390 21490
rect 14390 21420 14460 21490
rect 14460 21420 14480 21490
rect 14480 21420 14550 21490
rect 14550 21420 14560 21490
rect 14650 21420 14660 21490
rect 14660 21420 14730 21490
rect 14730 21420 14750 21490
rect 14750 21420 14820 21490
rect 14820 21420 14840 21490
rect 14840 21420 14890 21490
rect 14980 21420 15000 21490
rect 15000 21420 15020 21490
rect 15020 21420 15090 21490
rect 15090 21420 15110 21490
rect 15110 21420 15180 21490
rect 15180 21420 15200 21490
rect 15200 21420 15220 21490
rect 15310 21420 15360 21490
rect 15360 21420 15380 21490
rect 15380 21420 15450 21490
rect 15450 21420 15470 21490
rect 15470 21420 15540 21490
rect 15540 21420 15550 21490
rect 15640 21420 15650 21490
rect 15650 21420 15720 21490
rect 15720 21420 15740 21490
rect 15740 21420 15810 21490
rect 15810 21420 15830 21490
rect 15830 21420 15880 21490
rect 15970 21420 15990 21490
rect 15990 21420 16010 21490
rect 16010 21420 16080 21490
rect 16080 21420 16100 21490
rect 16100 21420 16170 21490
rect 16170 21420 16190 21490
rect 16190 21420 16210 21490
rect 16300 21420 16350 21490
rect 16350 21420 16370 21490
rect 16370 21420 16440 21490
rect 16440 21420 16460 21490
rect 16460 21420 16530 21490
rect 16530 21420 16540 21490
rect 16670 21420 16680 21490
rect 16680 21420 16750 21490
rect 16750 21420 16770 21490
rect 16770 21420 16840 21490
rect 16840 21420 16860 21490
rect 16860 21420 16910 21490
rect 17000 21420 17020 21490
rect 17020 21420 17040 21490
rect 17040 21420 17110 21490
rect 17110 21420 17130 21490
rect 17130 21420 17200 21490
rect 17200 21420 17220 21490
rect 17220 21420 17240 21490
rect 17330 21420 17380 21490
rect 17380 21420 17400 21490
rect 17400 21420 17470 21490
rect 17470 21420 17490 21490
rect 17490 21420 17560 21490
rect 17560 21420 17570 21490
rect 17660 21420 17670 21490
rect 17670 21420 17740 21490
rect 17740 21420 17760 21490
rect 17760 21420 17830 21490
rect 17830 21420 17850 21490
rect 17850 21420 17900 21490
rect 17990 21420 18010 21490
rect 18010 21420 18030 21490
rect 18030 21420 18100 21490
rect 18100 21420 18120 21490
rect 18120 21420 18190 21490
rect 18190 21420 18210 21490
rect 18210 21420 18230 21490
rect 18320 21420 18370 21490
rect 18370 21420 18390 21490
rect 18390 21420 18460 21490
rect 18460 21420 18480 21490
rect 18480 21420 18550 21490
rect 18550 21420 18560 21490
rect 18650 21420 18660 21490
rect 18660 21420 18730 21490
rect 18730 21420 18750 21490
rect 18750 21420 18820 21490
rect 18820 21420 18840 21490
rect 18840 21420 18890 21490
rect 18980 21420 19000 21490
rect 19000 21420 19020 21490
rect 19020 21420 19090 21490
rect 19090 21420 19110 21490
rect 19110 21420 19180 21490
rect 19180 21420 19200 21490
rect 19200 21420 19220 21490
rect 19310 21420 19360 21490
rect 19360 21420 19380 21490
rect 19380 21420 19450 21490
rect 19450 21420 19470 21490
rect 19470 21420 19540 21490
rect 19540 21420 19550 21490
rect 7640 21400 7880 21420
rect 7970 21400 8210 21420
rect 8300 21400 8540 21420
rect 8630 21400 8870 21420
rect 8960 21400 9200 21420
rect 9290 21400 9530 21420
rect 9620 21400 9860 21420
rect 9950 21400 10190 21420
rect 10280 21400 10520 21420
rect 10650 21400 10890 21420
rect 10980 21400 11220 21420
rect 11310 21400 11550 21420
rect 11640 21400 11880 21420
rect 11970 21400 12210 21420
rect 12300 21400 12540 21420
rect 12630 21400 12870 21420
rect 12960 21400 13200 21420
rect 13290 21400 13530 21420
rect 13660 21400 13900 21420
rect 13990 21400 14230 21420
rect 14320 21400 14560 21420
rect 14650 21400 14890 21420
rect 14980 21400 15220 21420
rect 15310 21400 15550 21420
rect 15640 21400 15880 21420
rect 15970 21400 16210 21420
rect 16300 21400 16540 21420
rect 16670 21400 16910 21420
rect 17000 21400 17240 21420
rect 17330 21400 17570 21420
rect 17660 21400 17900 21420
rect 17990 21400 18230 21420
rect 18320 21400 18560 21420
rect 18650 21400 18890 21420
rect 18980 21400 19220 21420
rect 19310 21400 19550 21420
rect 7640 21370 7650 21400
rect 7650 21370 7720 21400
rect 7720 21370 7740 21400
rect 7740 21370 7810 21400
rect 7810 21370 7830 21400
rect 7830 21370 7880 21400
rect 7970 21370 7990 21400
rect 7990 21370 8010 21400
rect 8010 21370 8080 21400
rect 8080 21370 8100 21400
rect 8100 21370 8170 21400
rect 8170 21370 8190 21400
rect 8190 21370 8210 21400
rect 8300 21370 8350 21400
rect 8350 21370 8370 21400
rect 8370 21370 8440 21400
rect 8440 21370 8460 21400
rect 8460 21370 8530 21400
rect 8530 21370 8540 21400
rect 8630 21370 8640 21400
rect 8640 21370 8710 21400
rect 8710 21370 8730 21400
rect 8730 21370 8800 21400
rect 8800 21370 8820 21400
rect 8820 21370 8870 21400
rect 8960 21370 8980 21400
rect 8980 21370 9000 21400
rect 9000 21370 9070 21400
rect 9070 21370 9090 21400
rect 9090 21370 9160 21400
rect 9160 21370 9180 21400
rect 9180 21370 9200 21400
rect 9290 21370 9340 21400
rect 9340 21370 9360 21400
rect 9360 21370 9430 21400
rect 9430 21370 9450 21400
rect 9450 21370 9520 21400
rect 9520 21370 9530 21400
rect 9620 21370 9630 21400
rect 9630 21370 9700 21400
rect 9700 21370 9720 21400
rect 9720 21370 9790 21400
rect 9790 21370 9810 21400
rect 9810 21370 9860 21400
rect 9950 21370 9970 21400
rect 9970 21370 9990 21400
rect 9990 21370 10060 21400
rect 10060 21370 10080 21400
rect 10080 21370 10150 21400
rect 10150 21370 10170 21400
rect 10170 21370 10190 21400
rect 10280 21370 10330 21400
rect 10330 21370 10350 21400
rect 10350 21370 10420 21400
rect 10420 21370 10440 21400
rect 10440 21370 10510 21400
rect 10510 21370 10520 21400
rect 10650 21370 10660 21400
rect 10660 21370 10730 21400
rect 10730 21370 10750 21400
rect 10750 21370 10820 21400
rect 10820 21370 10840 21400
rect 10840 21370 10890 21400
rect 10980 21370 11000 21400
rect 11000 21370 11020 21400
rect 11020 21370 11090 21400
rect 11090 21370 11110 21400
rect 11110 21370 11180 21400
rect 11180 21370 11200 21400
rect 11200 21370 11220 21400
rect 11310 21370 11360 21400
rect 11360 21370 11380 21400
rect 11380 21370 11450 21400
rect 11450 21370 11470 21400
rect 11470 21370 11540 21400
rect 11540 21370 11550 21400
rect 11640 21370 11650 21400
rect 11650 21370 11720 21400
rect 11720 21370 11740 21400
rect 11740 21370 11810 21400
rect 11810 21370 11830 21400
rect 11830 21370 11880 21400
rect 11970 21370 11990 21400
rect 11990 21370 12010 21400
rect 12010 21370 12080 21400
rect 12080 21370 12100 21400
rect 12100 21370 12170 21400
rect 12170 21370 12190 21400
rect 12190 21370 12210 21400
rect 12300 21370 12350 21400
rect 12350 21370 12370 21400
rect 12370 21370 12440 21400
rect 12440 21370 12460 21400
rect 12460 21370 12530 21400
rect 12530 21370 12540 21400
rect 12630 21370 12640 21400
rect 12640 21370 12710 21400
rect 12710 21370 12730 21400
rect 12730 21370 12800 21400
rect 12800 21370 12820 21400
rect 12820 21370 12870 21400
rect 12960 21370 12980 21400
rect 12980 21370 13000 21400
rect 13000 21370 13070 21400
rect 13070 21370 13090 21400
rect 13090 21370 13160 21400
rect 13160 21370 13180 21400
rect 13180 21370 13200 21400
rect 13290 21370 13340 21400
rect 13340 21370 13360 21400
rect 13360 21370 13430 21400
rect 13430 21370 13450 21400
rect 13450 21370 13520 21400
rect 13520 21370 13530 21400
rect 13660 21370 13670 21400
rect 13670 21370 13740 21400
rect 13740 21370 13760 21400
rect 13760 21370 13830 21400
rect 13830 21370 13850 21400
rect 13850 21370 13900 21400
rect 13990 21370 14010 21400
rect 14010 21370 14030 21400
rect 14030 21370 14100 21400
rect 14100 21370 14120 21400
rect 14120 21370 14190 21400
rect 14190 21370 14210 21400
rect 14210 21370 14230 21400
rect 14320 21370 14370 21400
rect 14370 21370 14390 21400
rect 14390 21370 14460 21400
rect 14460 21370 14480 21400
rect 14480 21370 14550 21400
rect 14550 21370 14560 21400
rect 14650 21370 14660 21400
rect 14660 21370 14730 21400
rect 14730 21370 14750 21400
rect 14750 21370 14820 21400
rect 14820 21370 14840 21400
rect 14840 21370 14890 21400
rect 14980 21370 15000 21400
rect 15000 21370 15020 21400
rect 15020 21370 15090 21400
rect 15090 21370 15110 21400
rect 15110 21370 15180 21400
rect 15180 21370 15200 21400
rect 15200 21370 15220 21400
rect 15310 21370 15360 21400
rect 15360 21370 15380 21400
rect 15380 21370 15450 21400
rect 15450 21370 15470 21400
rect 15470 21370 15540 21400
rect 15540 21370 15550 21400
rect 15640 21370 15650 21400
rect 15650 21370 15720 21400
rect 15720 21370 15740 21400
rect 15740 21370 15810 21400
rect 15810 21370 15830 21400
rect 15830 21370 15880 21400
rect 15970 21370 15990 21400
rect 15990 21370 16010 21400
rect 16010 21370 16080 21400
rect 16080 21370 16100 21400
rect 16100 21370 16170 21400
rect 16170 21370 16190 21400
rect 16190 21370 16210 21400
rect 16300 21370 16350 21400
rect 16350 21370 16370 21400
rect 16370 21370 16440 21400
rect 16440 21370 16460 21400
rect 16460 21370 16530 21400
rect 16530 21370 16540 21400
rect 16670 21370 16680 21400
rect 16680 21370 16750 21400
rect 16750 21370 16770 21400
rect 16770 21370 16840 21400
rect 16840 21370 16860 21400
rect 16860 21370 16910 21400
rect 17000 21370 17020 21400
rect 17020 21370 17040 21400
rect 17040 21370 17110 21400
rect 17110 21370 17130 21400
rect 17130 21370 17200 21400
rect 17200 21370 17220 21400
rect 17220 21370 17240 21400
rect 17330 21370 17380 21400
rect 17380 21370 17400 21400
rect 17400 21370 17470 21400
rect 17470 21370 17490 21400
rect 17490 21370 17560 21400
rect 17560 21370 17570 21400
rect 17660 21370 17670 21400
rect 17670 21370 17740 21400
rect 17740 21370 17760 21400
rect 17760 21370 17830 21400
rect 17830 21370 17850 21400
rect 17850 21370 17900 21400
rect 17990 21370 18010 21400
rect 18010 21370 18030 21400
rect 18030 21370 18100 21400
rect 18100 21370 18120 21400
rect 18120 21370 18190 21400
rect 18190 21370 18210 21400
rect 18210 21370 18230 21400
rect 18320 21370 18370 21400
rect 18370 21370 18390 21400
rect 18390 21370 18460 21400
rect 18460 21370 18480 21400
rect 18480 21370 18550 21400
rect 18550 21370 18560 21400
rect 18650 21370 18660 21400
rect 18660 21370 18730 21400
rect 18730 21370 18750 21400
rect 18750 21370 18820 21400
rect 18820 21370 18840 21400
rect 18840 21370 18890 21400
rect 18980 21370 19000 21400
rect 19000 21370 19020 21400
rect 19020 21370 19090 21400
rect 19090 21370 19110 21400
rect 19110 21370 19180 21400
rect 19180 21370 19200 21400
rect 19200 21370 19220 21400
rect 19310 21370 19360 21400
rect 19360 21370 19380 21400
rect 19380 21370 19450 21400
rect 19450 21370 19470 21400
rect 19470 21370 19540 21400
rect 19540 21370 19550 21400
rect 1720 6850 1960 6910
rect 2050 6850 2290 6910
rect 2390 6850 2630 6910
rect 2720 6850 2960 6910
rect 1720 6780 1750 6850
rect 1750 6780 1790 6850
rect 1790 6780 1860 6850
rect 1860 6780 1900 6850
rect 1900 6780 1960 6850
rect 2050 6780 2080 6850
rect 2080 6780 2120 6850
rect 2120 6780 2190 6850
rect 2190 6780 2230 6850
rect 2230 6780 2290 6850
rect 2390 6780 2410 6850
rect 2410 6780 2450 6850
rect 2450 6780 2520 6850
rect 2520 6780 2560 6850
rect 2560 6780 2630 6850
rect 2720 6780 2740 6850
rect 2740 6780 2780 6850
rect 2780 6780 2850 6850
rect 2850 6780 2890 6850
rect 2890 6780 2960 6850
rect 1720 6740 1960 6780
rect 2050 6740 2290 6780
rect 2390 6740 2630 6780
rect 2720 6740 2960 6780
rect 1720 6670 1750 6740
rect 1750 6670 1790 6740
rect 1790 6670 1860 6740
rect 1860 6670 1900 6740
rect 1900 6670 1960 6740
rect 2050 6670 2080 6740
rect 2080 6670 2120 6740
rect 2120 6670 2190 6740
rect 2190 6670 2230 6740
rect 2230 6670 2290 6740
rect 2390 6670 2410 6740
rect 2410 6670 2450 6740
rect 2450 6670 2520 6740
rect 2520 6670 2560 6740
rect 2560 6670 2630 6740
rect 2720 6670 2740 6740
rect 2740 6670 2780 6740
rect 2780 6670 2850 6740
rect 2850 6670 2890 6740
rect 2890 6670 2960 6740
rect 11940 6880 12180 6940
rect 12270 6880 12510 6940
rect 12610 6880 12850 6940
rect 12940 6880 13180 6940
rect 11940 6810 11970 6880
rect 11970 6810 12010 6880
rect 12010 6810 12080 6880
rect 12080 6810 12120 6880
rect 12120 6810 12180 6880
rect 12270 6810 12300 6880
rect 12300 6810 12340 6880
rect 12340 6810 12410 6880
rect 12410 6810 12450 6880
rect 12450 6810 12510 6880
rect 12610 6810 12630 6880
rect 12630 6810 12670 6880
rect 12670 6810 12740 6880
rect 12740 6810 12780 6880
rect 12780 6810 12850 6880
rect 12940 6810 12960 6880
rect 12960 6810 13000 6880
rect 13000 6810 13070 6880
rect 13070 6810 13110 6880
rect 13110 6810 13180 6880
rect 11940 6770 12180 6810
rect 12270 6770 12510 6810
rect 12610 6770 12850 6810
rect 12940 6770 13180 6810
rect 11940 6700 11970 6770
rect 11970 6700 12010 6770
rect 12010 6700 12080 6770
rect 12080 6700 12120 6770
rect 12120 6700 12180 6770
rect 12270 6700 12300 6770
rect 12300 6700 12340 6770
rect 12340 6700 12410 6770
rect 12410 6700 12450 6770
rect 12450 6700 12510 6770
rect 12610 6700 12630 6770
rect 12630 6700 12670 6770
rect 12670 6700 12740 6770
rect 12740 6700 12780 6770
rect 12780 6700 12850 6770
rect 12940 6700 12960 6770
rect 12960 6700 13000 6770
rect 13000 6700 13070 6770
rect 13070 6700 13110 6770
rect 13110 6700 13180 6770
rect 23510 7210 23880 7270
rect 23510 7140 23560 7210
rect 23560 7140 23600 7210
rect 23600 7140 23670 7210
rect 23670 7140 23710 7210
rect 23710 7140 23780 7210
rect 23780 7140 23820 7210
rect 23820 7140 23880 7210
rect 23510 7100 23880 7140
rect 23510 7030 23560 7100
rect 23560 7030 23600 7100
rect 23600 7030 23670 7100
rect 23670 7030 23710 7100
rect 23710 7030 23780 7100
rect 23780 7030 23820 7100
rect 23820 7030 23880 7100
rect 25910 7210 26280 7270
rect 25910 7140 25960 7210
rect 25960 7140 26000 7210
rect 26000 7140 26070 7210
rect 26070 7140 26110 7210
rect 26110 7140 26180 7210
rect 26180 7140 26220 7210
rect 26220 7140 26280 7210
rect 25910 7100 26280 7140
rect 25910 7030 25960 7100
rect 25960 7030 26000 7100
rect 26000 7030 26070 7100
rect 26070 7030 26110 7100
rect 26110 7030 26180 7100
rect 26180 7030 26220 7100
rect 26220 7030 26280 7100
rect 1260 -860 1330 -790
rect 1330 -860 1370 -790
rect 1370 -860 1440 -790
rect 1440 -860 1480 -790
rect 1480 -860 1500 -790
rect 1590 -860 1660 -790
rect 1660 -860 1700 -790
rect 1700 -860 1770 -790
rect 1770 -860 1810 -790
rect 1810 -860 1830 -790
rect 1930 -860 1990 -790
rect 1990 -860 2030 -790
rect 2030 -860 2100 -790
rect 2100 -860 2140 -790
rect 2140 -860 2170 -790
rect 2260 -860 2320 -790
rect 2320 -860 2360 -790
rect 2360 -860 2430 -790
rect 2430 -860 2470 -790
rect 2470 -860 2500 -790
rect 1260 -900 1500 -860
rect 1590 -900 1830 -860
rect 1930 -900 2170 -860
rect 2260 -900 2500 -860
rect 1260 -970 1330 -900
rect 1330 -970 1370 -900
rect 1370 -970 1440 -900
rect 1440 -970 1480 -900
rect 1480 -970 1500 -900
rect 1590 -970 1660 -900
rect 1660 -970 1700 -900
rect 1700 -970 1770 -900
rect 1770 -970 1810 -900
rect 1810 -970 1830 -900
rect 1930 -970 1990 -900
rect 1990 -970 2030 -900
rect 2030 -970 2100 -900
rect 2100 -970 2140 -900
rect 2140 -970 2170 -900
rect 2260 -970 2320 -900
rect 2320 -970 2360 -900
rect 2360 -970 2430 -900
rect 2430 -970 2470 -900
rect 2470 -970 2500 -900
rect 1260 -1030 1500 -970
rect 1590 -1030 1830 -970
rect 1930 -1030 2170 -970
rect 2260 -1030 2500 -970
rect 12400 -860 12430 -790
rect 12430 -860 12470 -790
rect 12470 -860 12540 -790
rect 12540 -860 12580 -790
rect 12580 -860 12640 -790
rect 12730 -860 12760 -790
rect 12760 -860 12800 -790
rect 12800 -860 12870 -790
rect 12870 -860 12910 -790
rect 12910 -860 12970 -790
rect 13070 -860 13090 -790
rect 13090 -860 13130 -790
rect 13130 -860 13200 -790
rect 13200 -860 13240 -790
rect 13240 -860 13310 -790
rect 13400 -860 13420 -790
rect 13420 -860 13460 -790
rect 13460 -860 13530 -790
rect 13530 -860 13570 -790
rect 13570 -860 13640 -790
rect 12400 -900 12640 -860
rect 12730 -900 12970 -860
rect 13070 -900 13310 -860
rect 13400 -900 13640 -860
rect 12400 -970 12430 -900
rect 12430 -970 12470 -900
rect 12470 -970 12540 -900
rect 12540 -970 12580 -900
rect 12580 -970 12640 -900
rect 12730 -970 12760 -900
rect 12760 -970 12800 -900
rect 12800 -970 12870 -900
rect 12870 -970 12910 -900
rect 12910 -970 12970 -900
rect 13070 -970 13090 -900
rect 13090 -970 13130 -900
rect 13130 -970 13200 -900
rect 13200 -970 13240 -900
rect 13240 -970 13310 -900
rect 13400 -970 13420 -900
rect 13420 -970 13460 -900
rect 13460 -970 13530 -900
rect 13530 -970 13570 -900
rect 13570 -970 13640 -900
rect 12400 -1030 12640 -970
rect 12730 -1030 12970 -970
rect 13070 -1030 13310 -970
rect 13400 -1030 13640 -970
rect 1720 -2780 1960 -2720
rect 2050 -2780 2290 -2720
rect 2390 -2780 2630 -2720
rect 2720 -2780 2960 -2720
rect 1720 -2850 1750 -2780
rect 1750 -2850 1790 -2780
rect 1790 -2850 1860 -2780
rect 1860 -2850 1900 -2780
rect 1900 -2850 1960 -2780
rect 2050 -2850 2080 -2780
rect 2080 -2850 2120 -2780
rect 2120 -2850 2190 -2780
rect 2190 -2850 2230 -2780
rect 2230 -2850 2290 -2780
rect 2390 -2850 2410 -2780
rect 2410 -2850 2450 -2780
rect 2450 -2850 2520 -2780
rect 2520 -2850 2560 -2780
rect 2560 -2850 2630 -2780
rect 2720 -2850 2740 -2780
rect 2740 -2850 2780 -2780
rect 2780 -2850 2850 -2780
rect 2850 -2850 2890 -2780
rect 2890 -2850 2960 -2780
rect 1720 -2890 1960 -2850
rect 2050 -2890 2290 -2850
rect 2390 -2890 2630 -2850
rect 2720 -2890 2960 -2850
rect 1720 -2960 1750 -2890
rect 1750 -2960 1790 -2890
rect 1790 -2960 1860 -2890
rect 1860 -2960 1900 -2890
rect 1900 -2960 1960 -2890
rect 2050 -2960 2080 -2890
rect 2080 -2960 2120 -2890
rect 2120 -2960 2190 -2890
rect 2190 -2960 2230 -2890
rect 2230 -2960 2290 -2890
rect 2390 -2960 2410 -2890
rect 2410 -2960 2450 -2890
rect 2450 -2960 2520 -2890
rect 2520 -2960 2560 -2890
rect 2560 -2960 2630 -2890
rect 2720 -2960 2740 -2890
rect 2740 -2960 2780 -2890
rect 2780 -2960 2850 -2890
rect 2850 -2960 2890 -2890
rect 2890 -2960 2960 -2890
rect 11940 -2780 12180 -2720
rect 12270 -2780 12510 -2720
rect 12610 -2780 12850 -2720
rect 12940 -2780 13180 -2720
rect 11940 -2850 11970 -2780
rect 11970 -2850 12010 -2780
rect 12010 -2850 12080 -2780
rect 12080 -2850 12120 -2780
rect 12120 -2850 12180 -2780
rect 12270 -2850 12300 -2780
rect 12300 -2850 12340 -2780
rect 12340 -2850 12410 -2780
rect 12410 -2850 12450 -2780
rect 12450 -2850 12510 -2780
rect 12610 -2850 12630 -2780
rect 12630 -2850 12670 -2780
rect 12670 -2850 12740 -2780
rect 12740 -2850 12780 -2780
rect 12780 -2850 12850 -2780
rect 12940 -2850 12960 -2780
rect 12960 -2850 13000 -2780
rect 13000 -2850 13070 -2780
rect 13070 -2850 13110 -2780
rect 13110 -2850 13180 -2780
rect 11940 -2890 12180 -2850
rect 12270 -2890 12510 -2850
rect 12610 -2890 12850 -2850
rect 12940 -2890 13180 -2850
rect 11940 -2960 11970 -2890
rect 11970 -2960 12010 -2890
rect 12010 -2960 12080 -2890
rect 12080 -2960 12120 -2890
rect 12120 -2960 12180 -2890
rect 12270 -2960 12300 -2890
rect 12300 -2960 12340 -2890
rect 12340 -2960 12410 -2890
rect 12410 -2960 12450 -2890
rect 12450 -2960 12510 -2890
rect 12610 -2960 12630 -2890
rect 12630 -2960 12670 -2890
rect 12670 -2960 12740 -2890
rect 12740 -2960 12780 -2890
rect 12780 -2960 12850 -2890
rect 12940 -2960 12960 -2890
rect 12960 -2960 13000 -2890
rect 13000 -2960 13070 -2890
rect 13070 -2960 13110 -2890
rect 13110 -2960 13180 -2890
rect 22480 2530 22540 2600
rect 22540 2530 22580 2600
rect 22580 2530 22650 2600
rect 22650 2530 22690 2600
rect 22690 2530 22760 2600
rect 22760 2530 22800 2600
rect 22800 2530 22850 2600
rect 22480 2490 22850 2530
rect 22480 2420 22540 2490
rect 22540 2420 22580 2490
rect 22580 2420 22650 2490
rect 22650 2420 22690 2490
rect 22690 2420 22760 2490
rect 22760 2420 22800 2490
rect 22800 2420 22850 2490
rect 22480 2360 22850 2420
rect 26960 2530 27020 2600
rect 27020 2530 27060 2600
rect 27060 2530 27130 2600
rect 27130 2530 27170 2600
rect 27170 2530 27240 2600
rect 27240 2530 27280 2600
rect 27280 2530 27330 2600
rect 26960 2490 27330 2530
rect 26960 2420 27020 2490
rect 27020 2420 27060 2490
rect 27060 2420 27130 2490
rect 27130 2420 27170 2490
rect 27170 2420 27240 2490
rect 27240 2420 27280 2490
rect 27280 2420 27330 2490
rect 26960 2360 27330 2420
rect 23510 920 23880 980
rect 23510 850 23560 920
rect 23560 850 23600 920
rect 23600 850 23670 920
rect 23670 850 23710 920
rect 23710 850 23780 920
rect 23780 850 23820 920
rect 23820 850 23880 920
rect 23510 810 23880 850
rect 23510 740 23560 810
rect 23560 740 23600 810
rect 23600 740 23670 810
rect 23670 740 23710 810
rect 23710 740 23780 810
rect 23780 740 23820 810
rect 23820 740 23880 810
rect 25910 920 26280 980
rect 25910 850 25960 920
rect 25960 850 26000 920
rect 26000 850 26070 920
rect 26070 850 26110 920
rect 26110 850 26180 920
rect 26180 850 26220 920
rect 26220 850 26280 920
rect 25910 810 26280 850
rect 25910 740 25960 810
rect 25960 740 26000 810
rect 26000 740 26070 810
rect 26070 740 26110 810
rect 26110 740 26180 810
rect 26180 740 26220 810
rect 26220 740 26280 810
rect 38230 7750 38260 7770
rect 38260 7750 38280 7770
rect 38280 7750 38350 7770
rect 38350 7750 38370 7770
rect 38370 7750 38440 7770
rect 38440 7750 38470 7770
rect 38230 7730 38470 7750
rect 38230 7660 38260 7730
rect 38260 7660 38280 7730
rect 38280 7660 38350 7730
rect 38350 7660 38370 7730
rect 38370 7660 38440 7730
rect 38440 7660 38470 7730
rect 38230 7640 38470 7660
rect 38230 7570 38260 7640
rect 38260 7570 38280 7640
rect 38280 7570 38350 7640
rect 38350 7570 38370 7640
rect 38370 7570 38440 7640
rect 38440 7570 38470 7640
rect 38230 7550 38470 7570
rect 38230 7530 38260 7550
rect 38260 7530 38280 7550
rect 38280 7530 38350 7550
rect 38350 7530 38370 7550
rect 38370 7530 38440 7550
rect 38440 7530 38470 7550
rect 38230 7390 38260 7440
rect 38260 7390 38280 7440
rect 38280 7390 38350 7440
rect 38350 7390 38370 7440
rect 38370 7390 38440 7440
rect 38440 7390 38470 7440
rect 38230 7370 38470 7390
rect 38230 7300 38260 7370
rect 38260 7300 38280 7370
rect 38280 7300 38350 7370
rect 38350 7300 38370 7370
rect 38370 7300 38440 7370
rect 38440 7300 38470 7370
rect 38230 7280 38470 7300
rect 38230 7210 38260 7280
rect 38260 7210 38280 7280
rect 38280 7210 38350 7280
rect 38350 7210 38370 7280
rect 38370 7210 38440 7280
rect 38440 7210 38470 7280
rect 38230 7200 38470 7210
rect 38230 7060 38470 7070
rect 38230 6990 38260 7060
rect 38260 6990 38280 7060
rect 38280 6990 38350 7060
rect 38350 6990 38370 7060
rect 38370 6990 38440 7060
rect 38440 6990 38470 7060
rect 38230 6970 38470 6990
rect 38230 6900 38260 6970
rect 38260 6900 38280 6970
rect 38280 6900 38350 6970
rect 38350 6900 38370 6970
rect 38370 6900 38440 6970
rect 38440 6900 38470 6970
rect 38230 6880 38470 6900
rect 38230 6830 38260 6880
rect 38260 6830 38280 6880
rect 38280 6830 38350 6880
rect 38350 6830 38370 6880
rect 38370 6830 38440 6880
rect 38440 6830 38470 6880
rect 38230 6720 38260 6740
rect 38260 6720 38280 6740
rect 38280 6720 38350 6740
rect 38350 6720 38370 6740
rect 38370 6720 38440 6740
rect 38440 6720 38470 6740
rect 38230 6700 38470 6720
rect 38230 6630 38260 6700
rect 38260 6630 38280 6700
rect 38280 6630 38350 6700
rect 38350 6630 38370 6700
rect 38370 6630 38440 6700
rect 38440 6630 38470 6700
rect 38230 6610 38470 6630
rect 38230 6540 38260 6610
rect 38260 6540 38280 6610
rect 38280 6540 38350 6610
rect 38350 6540 38370 6610
rect 38370 6540 38440 6610
rect 38440 6540 38470 6610
rect 38230 6520 38470 6540
rect 38230 6500 38260 6520
rect 38260 6500 38280 6520
rect 38280 6500 38350 6520
rect 38350 6500 38370 6520
rect 38370 6500 38440 6520
rect 38440 6500 38470 6520
rect 38230 6360 38260 6410
rect 38260 6360 38280 6410
rect 38280 6360 38350 6410
rect 38350 6360 38370 6410
rect 38370 6360 38440 6410
rect 38440 6360 38470 6410
rect 38230 6340 38470 6360
rect 38230 6270 38260 6340
rect 38260 6270 38280 6340
rect 38280 6270 38350 6340
rect 38350 6270 38370 6340
rect 38370 6270 38440 6340
rect 38440 6270 38470 6340
rect 38230 6250 38470 6270
rect 38230 6180 38260 6250
rect 38260 6180 38280 6250
rect 38280 6180 38350 6250
rect 38350 6180 38370 6250
rect 38370 6180 38440 6250
rect 38440 6180 38470 6250
rect 38230 6170 38470 6180
rect 38230 6070 38470 6080
rect 38230 6000 38260 6070
rect 38260 6000 38280 6070
rect 38280 6000 38350 6070
rect 38350 6000 38370 6070
rect 38370 6000 38440 6070
rect 38440 6000 38470 6070
rect 38230 5980 38470 6000
rect 38230 5910 38260 5980
rect 38260 5910 38280 5980
rect 38280 5910 38350 5980
rect 38350 5910 38370 5980
rect 38370 5910 38440 5980
rect 38440 5910 38470 5980
rect 38230 5890 38470 5910
rect 38230 5840 38260 5890
rect 38260 5840 38280 5890
rect 38280 5840 38350 5890
rect 38350 5840 38370 5890
rect 38370 5840 38440 5890
rect 38440 5840 38470 5890
rect 38230 5730 38260 5750
rect 38260 5730 38280 5750
rect 38280 5730 38350 5750
rect 38350 5730 38370 5750
rect 38370 5730 38440 5750
rect 38440 5730 38470 5750
rect 38230 5710 38470 5730
rect 38230 5640 38260 5710
rect 38260 5640 38280 5710
rect 38280 5640 38350 5710
rect 38350 5640 38370 5710
rect 38370 5640 38440 5710
rect 38440 5640 38470 5710
rect 38230 5620 38470 5640
rect 38230 5550 38260 5620
rect 38260 5550 38280 5620
rect 38280 5550 38350 5620
rect 38350 5550 38370 5620
rect 38370 5550 38440 5620
rect 38440 5550 38470 5620
rect 38230 5530 38470 5550
rect 38230 5510 38260 5530
rect 38260 5510 38280 5530
rect 38280 5510 38350 5530
rect 38350 5510 38370 5530
rect 38370 5510 38440 5530
rect 38440 5510 38470 5530
rect 38230 5370 38260 5420
rect 38260 5370 38280 5420
rect 38280 5370 38350 5420
rect 38350 5370 38370 5420
rect 38370 5370 38440 5420
rect 38440 5370 38470 5420
rect 38230 5350 38470 5370
rect 38230 5280 38260 5350
rect 38260 5280 38280 5350
rect 38280 5280 38350 5350
rect 38350 5280 38370 5350
rect 38370 5280 38440 5350
rect 38440 5280 38470 5350
rect 38230 5260 38470 5280
rect 38230 5190 38260 5260
rect 38260 5190 38280 5260
rect 38280 5190 38350 5260
rect 38350 5190 38370 5260
rect 38370 5190 38440 5260
rect 38440 5190 38470 5260
rect 38230 5180 38470 5190
rect 38230 5080 38470 5090
rect 38230 5010 38260 5080
rect 38260 5010 38280 5080
rect 38280 5010 38350 5080
rect 38350 5010 38370 5080
rect 38370 5010 38440 5080
rect 38440 5010 38470 5080
rect 38230 4990 38470 5010
rect 38230 4920 38260 4990
rect 38260 4920 38280 4990
rect 38280 4920 38350 4990
rect 38350 4920 38370 4990
rect 38370 4920 38440 4990
rect 38440 4920 38470 4990
rect 38230 4900 38470 4920
rect 38230 4850 38260 4900
rect 38260 4850 38280 4900
rect 38280 4850 38350 4900
rect 38350 4850 38370 4900
rect 38370 4850 38440 4900
rect 38440 4850 38470 4900
rect 38230 4740 38260 4760
rect 38260 4740 38280 4760
rect 38280 4740 38350 4760
rect 38350 4740 38370 4760
rect 38370 4740 38440 4760
rect 38440 4740 38470 4760
rect 38230 4720 38470 4740
rect 38230 4650 38260 4720
rect 38260 4650 38280 4720
rect 38280 4650 38350 4720
rect 38350 4650 38370 4720
rect 38370 4650 38440 4720
rect 38440 4650 38470 4720
rect 38230 4630 38470 4650
rect 38230 4560 38260 4630
rect 38260 4560 38280 4630
rect 38280 4560 38350 4630
rect 38350 4560 38370 4630
rect 38370 4560 38440 4630
rect 38440 4560 38470 4630
rect 38230 4540 38470 4560
rect 38230 4520 38260 4540
rect 38260 4520 38280 4540
rect 38280 4520 38350 4540
rect 38350 4520 38370 4540
rect 38370 4520 38440 4540
rect 38440 4520 38470 4540
rect 38230 4380 38260 4430
rect 38260 4380 38280 4430
rect 38280 4380 38350 4430
rect 38350 4380 38370 4430
rect 38370 4380 38440 4430
rect 38440 4380 38470 4430
rect 38230 4360 38470 4380
rect 38230 4290 38260 4360
rect 38260 4290 38280 4360
rect 38280 4290 38350 4360
rect 38350 4290 38370 4360
rect 38370 4290 38440 4360
rect 38440 4290 38470 4360
rect 38230 4270 38470 4290
rect 38230 4200 38260 4270
rect 38260 4200 38280 4270
rect 38280 4200 38350 4270
rect 38350 4200 38370 4270
rect 38370 4200 38440 4270
rect 38440 4200 38470 4270
rect 38230 4190 38470 4200
rect 38230 4050 38470 4060
rect 38230 3980 38260 4050
rect 38260 3980 38280 4050
rect 38280 3980 38350 4050
rect 38350 3980 38370 4050
rect 38370 3980 38440 4050
rect 38440 3980 38470 4050
rect 38230 3960 38470 3980
rect 38230 3890 38260 3960
rect 38260 3890 38280 3960
rect 38280 3890 38350 3960
rect 38350 3890 38370 3960
rect 38370 3890 38440 3960
rect 38440 3890 38470 3960
rect 38230 3870 38470 3890
rect 38230 3820 38260 3870
rect 38260 3820 38280 3870
rect 38280 3820 38350 3870
rect 38350 3820 38370 3870
rect 38370 3820 38440 3870
rect 38440 3820 38470 3870
rect 38230 3710 38260 3730
rect 38260 3710 38280 3730
rect 38280 3710 38350 3730
rect 38350 3710 38370 3730
rect 38370 3710 38440 3730
rect 38440 3710 38470 3730
rect 38230 3690 38470 3710
rect 38230 3620 38260 3690
rect 38260 3620 38280 3690
rect 38280 3620 38350 3690
rect 38350 3620 38370 3690
rect 38370 3620 38440 3690
rect 38440 3620 38470 3690
rect 38230 3600 38470 3620
rect 38230 3530 38260 3600
rect 38260 3530 38280 3600
rect 38280 3530 38350 3600
rect 38350 3530 38370 3600
rect 38370 3530 38440 3600
rect 38440 3530 38470 3600
rect 38230 3510 38470 3530
rect 38230 3490 38260 3510
rect 38260 3490 38280 3510
rect 38280 3490 38350 3510
rect 38350 3490 38370 3510
rect 38370 3490 38440 3510
rect 38440 3490 38470 3510
rect 38230 3350 38260 3400
rect 38260 3350 38280 3400
rect 38280 3350 38350 3400
rect 38350 3350 38370 3400
rect 38370 3350 38440 3400
rect 38440 3350 38470 3400
rect 38230 3330 38470 3350
rect 38230 3260 38260 3330
rect 38260 3260 38280 3330
rect 38280 3260 38350 3330
rect 38350 3260 38370 3330
rect 38370 3260 38440 3330
rect 38440 3260 38470 3330
rect 38230 3240 38470 3260
rect 38230 3170 38260 3240
rect 38260 3170 38280 3240
rect 38280 3170 38350 3240
rect 38350 3170 38370 3240
rect 38370 3170 38440 3240
rect 38440 3170 38470 3240
rect 38230 3160 38470 3170
rect 38230 3060 38470 3070
rect 38230 2990 38260 3060
rect 38260 2990 38280 3060
rect 38280 2990 38350 3060
rect 38350 2990 38370 3060
rect 38370 2990 38440 3060
rect 38440 2990 38470 3060
rect 38230 2970 38470 2990
rect 38230 2900 38260 2970
rect 38260 2900 38280 2970
rect 38280 2900 38350 2970
rect 38350 2900 38370 2970
rect 38370 2900 38440 2970
rect 38440 2900 38470 2970
rect 38230 2880 38470 2900
rect 38230 2830 38260 2880
rect 38260 2830 38280 2880
rect 38280 2830 38350 2880
rect 38350 2830 38370 2880
rect 38370 2830 38440 2880
rect 38440 2830 38470 2880
rect 38230 2720 38260 2740
rect 38260 2720 38280 2740
rect 38280 2720 38350 2740
rect 38350 2720 38370 2740
rect 38370 2720 38440 2740
rect 38440 2720 38470 2740
rect 38230 2700 38470 2720
rect 38230 2630 38260 2700
rect 38260 2630 38280 2700
rect 38280 2630 38350 2700
rect 38350 2630 38370 2700
rect 38370 2630 38440 2700
rect 38440 2630 38470 2700
rect 38230 2610 38470 2630
rect 38230 2540 38260 2610
rect 38260 2540 38280 2610
rect 38280 2540 38350 2610
rect 38350 2540 38370 2610
rect 38370 2540 38440 2610
rect 38440 2540 38470 2610
rect 38230 2520 38470 2540
rect 38230 2500 38260 2520
rect 38260 2500 38280 2520
rect 38280 2500 38350 2520
rect 38350 2500 38370 2520
rect 38370 2500 38440 2520
rect 38440 2500 38470 2520
rect 38230 2360 38260 2410
rect 38260 2360 38280 2410
rect 38280 2360 38350 2410
rect 38350 2360 38370 2410
rect 38370 2360 38440 2410
rect 38440 2360 38470 2410
rect 38230 2340 38470 2360
rect 38230 2270 38260 2340
rect 38260 2270 38280 2340
rect 38280 2270 38350 2340
rect 38350 2270 38370 2340
rect 38370 2270 38440 2340
rect 38440 2270 38470 2340
rect 38230 2250 38470 2270
rect 38230 2180 38260 2250
rect 38260 2180 38280 2250
rect 38280 2180 38350 2250
rect 38350 2180 38370 2250
rect 38370 2180 38440 2250
rect 38440 2180 38470 2250
rect 38230 2170 38470 2180
rect 38230 2070 38470 2080
rect 38230 2000 38260 2070
rect 38260 2000 38280 2070
rect 38280 2000 38350 2070
rect 38350 2000 38370 2070
rect 38370 2000 38440 2070
rect 38440 2000 38470 2070
rect 38230 1980 38470 2000
rect 38230 1910 38260 1980
rect 38260 1910 38280 1980
rect 38280 1910 38350 1980
rect 38350 1910 38370 1980
rect 38370 1910 38440 1980
rect 38440 1910 38470 1980
rect 38230 1890 38470 1910
rect 38230 1840 38260 1890
rect 38260 1840 38280 1890
rect 38280 1840 38350 1890
rect 38350 1840 38370 1890
rect 38370 1840 38440 1890
rect 38440 1840 38470 1890
rect 38230 1730 38260 1750
rect 38260 1730 38280 1750
rect 38280 1730 38350 1750
rect 38350 1730 38370 1750
rect 38370 1730 38440 1750
rect 38440 1730 38470 1750
rect 38230 1710 38470 1730
rect 38230 1640 38260 1710
rect 38260 1640 38280 1710
rect 38280 1640 38350 1710
rect 38350 1640 38370 1710
rect 38370 1640 38440 1710
rect 38440 1640 38470 1710
rect 38230 1620 38470 1640
rect 38230 1550 38260 1620
rect 38260 1550 38280 1620
rect 38280 1550 38350 1620
rect 38350 1550 38370 1620
rect 38370 1550 38440 1620
rect 38440 1550 38470 1620
rect 38230 1530 38470 1550
rect 38230 1510 38260 1530
rect 38260 1510 38280 1530
rect 38280 1510 38350 1530
rect 38350 1510 38370 1530
rect 38370 1510 38440 1530
rect 38440 1510 38470 1530
rect 38230 1370 38260 1420
rect 38260 1370 38280 1420
rect 38280 1370 38350 1420
rect 38350 1370 38370 1420
rect 38370 1370 38440 1420
rect 38440 1370 38470 1420
rect 38230 1350 38470 1370
rect 38230 1280 38260 1350
rect 38260 1280 38280 1350
rect 38280 1280 38350 1350
rect 38350 1280 38370 1350
rect 38370 1280 38440 1350
rect 38440 1280 38470 1350
rect 38230 1260 38470 1280
rect 38230 1190 38260 1260
rect 38260 1190 38280 1260
rect 38280 1190 38350 1260
rect 38350 1190 38370 1260
rect 38370 1190 38440 1260
rect 38440 1190 38470 1260
rect 38230 1180 38470 1190
rect 22480 -3760 22540 -3690
rect 22540 -3760 22580 -3690
rect 22580 -3760 22650 -3690
rect 22650 -3760 22690 -3690
rect 22690 -3760 22760 -3690
rect 22760 -3760 22800 -3690
rect 22800 -3760 22850 -3690
rect 22480 -3800 22850 -3760
rect 22480 -3870 22540 -3800
rect 22540 -3870 22580 -3800
rect 22580 -3870 22650 -3800
rect 22650 -3870 22690 -3800
rect 22690 -3870 22760 -3800
rect 22760 -3870 22800 -3800
rect 22800 -3870 22850 -3800
rect 22480 -3930 22850 -3870
rect 26960 -3760 27020 -3690
rect 27020 -3760 27060 -3690
rect 27060 -3760 27130 -3690
rect 27130 -3760 27170 -3690
rect 27170 -3760 27240 -3690
rect 27240 -3760 27280 -3690
rect 27280 -3760 27330 -3690
rect 26960 -3800 27330 -3760
rect 26960 -3870 27020 -3800
rect 27020 -3870 27060 -3800
rect 27060 -3870 27130 -3800
rect 27130 -3870 27170 -3800
rect 27170 -3870 27240 -3800
rect 27240 -3870 27280 -3800
rect 27280 -3870 27330 -3800
rect 26960 -3930 27330 -3870
rect -1170 -6400 -1160 -6370
rect -1160 -6400 -1090 -6370
rect -1090 -6400 -1070 -6370
rect -1070 -6400 -1000 -6370
rect -1000 -6400 -980 -6370
rect -980 -6400 -930 -6370
rect -840 -6400 -820 -6370
rect -820 -6400 -800 -6370
rect -800 -6400 -730 -6370
rect -730 -6400 -710 -6370
rect -710 -6400 -640 -6370
rect -640 -6400 -620 -6370
rect -620 -6400 -600 -6370
rect -510 -6400 -460 -6370
rect -460 -6400 -440 -6370
rect -440 -6400 -370 -6370
rect -370 -6400 -350 -6370
rect -350 -6400 -280 -6370
rect -280 -6400 -270 -6370
rect -180 -6400 -170 -6370
rect -170 -6400 -100 -6370
rect -100 -6400 -80 -6370
rect -80 -6400 -10 -6370
rect -10 -6400 10 -6370
rect 10 -6400 60 -6370
rect -1170 -6420 -930 -6400
rect -840 -6420 -600 -6400
rect -510 -6420 -270 -6400
rect -180 -6420 60 -6400
rect -1170 -6490 -1160 -6420
rect -1160 -6490 -1090 -6420
rect -1090 -6490 -1070 -6420
rect -1070 -6490 -1000 -6420
rect -1000 -6490 -980 -6420
rect -980 -6490 -930 -6420
rect -840 -6490 -820 -6420
rect -820 -6490 -800 -6420
rect -800 -6490 -730 -6420
rect -730 -6490 -710 -6420
rect -710 -6490 -640 -6420
rect -640 -6490 -620 -6420
rect -620 -6490 -600 -6420
rect -510 -6490 -460 -6420
rect -460 -6490 -440 -6420
rect -440 -6490 -370 -6420
rect -370 -6490 -350 -6420
rect -350 -6490 -280 -6420
rect -280 -6490 -270 -6420
rect -180 -6490 -170 -6420
rect -170 -6490 -100 -6420
rect -100 -6490 -80 -6420
rect -80 -6490 -10 -6420
rect -10 -6490 10 -6420
rect 10 -6490 60 -6420
rect -1170 -6510 -930 -6490
rect -840 -6510 -600 -6490
rect -510 -6510 -270 -6490
rect -180 -6510 60 -6490
rect -1170 -6580 -1160 -6510
rect -1160 -6580 -1090 -6510
rect -1090 -6580 -1070 -6510
rect -1070 -6580 -1000 -6510
rect -1000 -6580 -980 -6510
rect -980 -6580 -930 -6510
rect -840 -6580 -820 -6510
rect -820 -6580 -800 -6510
rect -800 -6580 -730 -6510
rect -730 -6580 -710 -6510
rect -710 -6580 -640 -6510
rect -640 -6580 -620 -6510
rect -620 -6580 -600 -6510
rect -510 -6580 -460 -6510
rect -460 -6580 -440 -6510
rect -440 -6580 -370 -6510
rect -370 -6580 -350 -6510
rect -350 -6580 -280 -6510
rect -280 -6580 -270 -6510
rect -180 -6580 -170 -6510
rect -170 -6580 -100 -6510
rect -100 -6580 -80 -6510
rect -80 -6580 -10 -6510
rect -10 -6580 10 -6510
rect 10 -6580 60 -6510
rect -1170 -6610 -930 -6580
rect -840 -6610 -600 -6580
rect -510 -6610 -270 -6580
rect -180 -6610 60 -6580
rect 14720 -6400 14770 -6370
rect 14770 -6400 14790 -6370
rect 14790 -6400 14860 -6370
rect 14860 -6400 14880 -6370
rect 14880 -6400 14950 -6370
rect 14950 -6400 14960 -6370
rect 15050 -6400 15060 -6370
rect 15060 -6400 15130 -6370
rect 15130 -6400 15150 -6370
rect 15150 -6400 15220 -6370
rect 15220 -6400 15240 -6370
rect 15240 -6400 15290 -6370
rect 15380 -6400 15400 -6370
rect 15400 -6400 15420 -6370
rect 15420 -6400 15490 -6370
rect 15490 -6400 15510 -6370
rect 15510 -6400 15580 -6370
rect 15580 -6400 15600 -6370
rect 15600 -6400 15620 -6370
rect 15710 -6400 15760 -6370
rect 15760 -6400 15780 -6370
rect 15780 -6400 15850 -6370
rect 15850 -6400 15870 -6370
rect 15870 -6400 15940 -6370
rect 15940 -6400 15950 -6370
rect 14720 -6420 14960 -6400
rect 15050 -6420 15290 -6400
rect 15380 -6420 15620 -6400
rect 15710 -6420 15950 -6400
rect 14720 -6490 14770 -6420
rect 14770 -6490 14790 -6420
rect 14790 -6490 14860 -6420
rect 14860 -6490 14880 -6420
rect 14880 -6490 14950 -6420
rect 14950 -6490 14960 -6420
rect 15050 -6490 15060 -6420
rect 15060 -6490 15130 -6420
rect 15130 -6490 15150 -6420
rect 15150 -6490 15220 -6420
rect 15220 -6490 15240 -6420
rect 15240 -6490 15290 -6420
rect 15380 -6490 15400 -6420
rect 15400 -6490 15420 -6420
rect 15420 -6490 15490 -6420
rect 15490 -6490 15510 -6420
rect 15510 -6490 15580 -6420
rect 15580 -6490 15600 -6420
rect 15600 -6490 15620 -6420
rect 15710 -6490 15760 -6420
rect 15760 -6490 15780 -6420
rect 15780 -6490 15850 -6420
rect 15850 -6490 15870 -6420
rect 15870 -6490 15940 -6420
rect 15940 -6490 15950 -6420
rect 14720 -6510 14960 -6490
rect 15050 -6510 15290 -6490
rect 15380 -6510 15620 -6490
rect 15710 -6510 15950 -6490
rect 14720 -6580 14770 -6510
rect 14770 -6580 14790 -6510
rect 14790 -6580 14860 -6510
rect 14860 -6580 14880 -6510
rect 14880 -6580 14950 -6510
rect 14950 -6580 14960 -6510
rect 15050 -6580 15060 -6510
rect 15060 -6580 15130 -6510
rect 15130 -6580 15150 -6510
rect 15150 -6580 15220 -6510
rect 15220 -6580 15240 -6510
rect 15240 -6580 15290 -6510
rect 15380 -6580 15400 -6510
rect 15400 -6580 15420 -6510
rect 15420 -6580 15490 -6510
rect 15490 -6580 15510 -6510
rect 15510 -6580 15580 -6510
rect 15580 -6580 15600 -6510
rect 15600 -6580 15620 -6510
rect 15710 -6580 15760 -6510
rect 15760 -6580 15780 -6510
rect 15780 -6580 15850 -6510
rect 15850 -6580 15870 -6510
rect 15870 -6580 15940 -6510
rect 15940 -6580 15950 -6510
rect 14720 -6610 14960 -6580
rect 15050 -6610 15290 -6580
rect 15380 -6610 15620 -6580
rect 15710 -6610 15950 -6580
rect 21650 -8430 21700 -8370
rect 21700 -8430 21730 -8370
rect 21730 -8430 21800 -8370
rect 21800 -8430 21830 -8370
rect 21830 -8430 21890 -8370
rect 21650 -8460 21890 -8430
rect 21650 -8530 21700 -8460
rect 21700 -8530 21730 -8460
rect 21730 -8530 21800 -8460
rect 21800 -8530 21830 -8460
rect 21830 -8530 21890 -8460
rect 21650 -8560 21890 -8530
rect 21650 -8610 21700 -8560
rect 21700 -8610 21730 -8560
rect 21730 -8610 21800 -8560
rect 21800 -8610 21830 -8560
rect 21830 -8610 21890 -8560
rect 1260 -10410 1330 -10340
rect 1330 -10410 1370 -10340
rect 1370 -10410 1440 -10340
rect 1440 -10410 1480 -10340
rect 1480 -10410 1500 -10340
rect 1590 -10410 1660 -10340
rect 1660 -10410 1700 -10340
rect 1700 -10410 1770 -10340
rect 1770 -10410 1810 -10340
rect 1810 -10410 1830 -10340
rect 1930 -10410 1990 -10340
rect 1990 -10410 2030 -10340
rect 2030 -10410 2100 -10340
rect 2100 -10410 2140 -10340
rect 2140 -10410 2170 -10340
rect 2260 -10410 2320 -10340
rect 2320 -10410 2360 -10340
rect 2360 -10410 2430 -10340
rect 2430 -10410 2470 -10340
rect 2470 -10410 2500 -10340
rect 1260 -10450 1500 -10410
rect 1590 -10450 1830 -10410
rect 1930 -10450 2170 -10410
rect 2260 -10450 2500 -10410
rect 1260 -10520 1330 -10450
rect 1330 -10520 1370 -10450
rect 1370 -10520 1440 -10450
rect 1440 -10520 1480 -10450
rect 1480 -10520 1500 -10450
rect 1590 -10520 1660 -10450
rect 1660 -10520 1700 -10450
rect 1700 -10520 1770 -10450
rect 1770 -10520 1810 -10450
rect 1810 -10520 1830 -10450
rect 1930 -10520 1990 -10450
rect 1990 -10520 2030 -10450
rect 2030 -10520 2100 -10450
rect 2100 -10520 2140 -10450
rect 2140 -10520 2170 -10450
rect 2260 -10520 2320 -10450
rect 2320 -10520 2360 -10450
rect 2360 -10520 2430 -10450
rect 2430 -10520 2470 -10450
rect 2470 -10520 2500 -10450
rect 1260 -10580 1500 -10520
rect 1590 -10580 1830 -10520
rect 1930 -10580 2170 -10520
rect 2260 -10580 2500 -10520
rect 12400 -10440 12470 -10370
rect 12470 -10440 12510 -10370
rect 12510 -10440 12580 -10370
rect 12580 -10440 12620 -10370
rect 12620 -10440 12640 -10370
rect 12730 -10440 12800 -10370
rect 12800 -10440 12840 -10370
rect 12840 -10440 12910 -10370
rect 12910 -10440 12950 -10370
rect 12950 -10440 12970 -10370
rect 13070 -10440 13130 -10370
rect 13130 -10440 13170 -10370
rect 13170 -10440 13240 -10370
rect 13240 -10440 13280 -10370
rect 13280 -10440 13310 -10370
rect 13400 -10440 13460 -10370
rect 13460 -10440 13500 -10370
rect 13500 -10440 13570 -10370
rect 13570 -10440 13610 -10370
rect 13610 -10440 13640 -10370
rect 12400 -10480 12640 -10440
rect 12730 -10480 12970 -10440
rect 13070 -10480 13310 -10440
rect 13400 -10480 13640 -10440
rect 12400 -10550 12470 -10480
rect 12470 -10550 12510 -10480
rect 12510 -10550 12580 -10480
rect 12580 -10550 12620 -10480
rect 12620 -10550 12640 -10480
rect 12730 -10550 12800 -10480
rect 12800 -10550 12840 -10480
rect 12840 -10550 12910 -10480
rect 12910 -10550 12950 -10480
rect 12950 -10550 12970 -10480
rect 13070 -10550 13130 -10480
rect 13130 -10550 13170 -10480
rect 13170 -10550 13240 -10480
rect 13240 -10550 13280 -10480
rect 13280 -10550 13310 -10480
rect 13400 -10550 13460 -10480
rect 13460 -10550 13500 -10480
rect 13500 -10550 13570 -10480
rect 13570 -10550 13610 -10480
rect 13610 -10550 13640 -10480
rect 12400 -10610 12640 -10550
rect 12730 -10610 12970 -10550
rect 13070 -10610 13310 -10550
rect 13400 -10610 13640 -10550
rect 38230 150 38260 170
rect 38260 150 38280 170
rect 38280 150 38350 170
rect 38350 150 38370 170
rect 38370 150 38440 170
rect 38440 150 38470 170
rect 38230 130 38470 150
rect 38230 60 38260 130
rect 38260 60 38280 130
rect 38280 60 38350 130
rect 38350 60 38370 130
rect 38370 60 38440 130
rect 38440 60 38470 130
rect 38230 40 38470 60
rect 38230 -30 38260 40
rect 38260 -30 38280 40
rect 38280 -30 38350 40
rect 38350 -30 38370 40
rect 38370 -30 38440 40
rect 38440 -30 38470 40
rect 38230 -50 38470 -30
rect 38230 -70 38260 -50
rect 38260 -70 38280 -50
rect 38280 -70 38350 -50
rect 38350 -70 38370 -50
rect 38370 -70 38440 -50
rect 38440 -70 38470 -50
rect 38230 -210 38260 -160
rect 38260 -210 38280 -160
rect 38280 -210 38350 -160
rect 38350 -210 38370 -160
rect 38370 -210 38440 -160
rect 38440 -210 38470 -160
rect 38230 -230 38470 -210
rect 38230 -300 38260 -230
rect 38260 -300 38280 -230
rect 38280 -300 38350 -230
rect 38350 -300 38370 -230
rect 38370 -300 38440 -230
rect 38440 -300 38470 -230
rect 38230 -320 38470 -300
rect 38230 -390 38260 -320
rect 38260 -390 38280 -320
rect 38280 -390 38350 -320
rect 38350 -390 38370 -320
rect 38370 -390 38440 -320
rect 38440 -390 38470 -320
rect 38230 -400 38470 -390
rect 38230 -540 38470 -530
rect 38230 -610 38260 -540
rect 38260 -610 38280 -540
rect 38280 -610 38350 -540
rect 38350 -610 38370 -540
rect 38370 -610 38440 -540
rect 38440 -610 38470 -540
rect 38230 -630 38470 -610
rect 38230 -700 38260 -630
rect 38260 -700 38280 -630
rect 38280 -700 38350 -630
rect 38350 -700 38370 -630
rect 38370 -700 38440 -630
rect 38440 -700 38470 -630
rect 38230 -720 38470 -700
rect 38230 -770 38260 -720
rect 38260 -770 38280 -720
rect 38280 -770 38350 -720
rect 38350 -770 38370 -720
rect 38370 -770 38440 -720
rect 38440 -770 38470 -720
rect 38230 -880 38260 -860
rect 38260 -880 38280 -860
rect 38280 -880 38350 -860
rect 38350 -880 38370 -860
rect 38370 -880 38440 -860
rect 38440 -880 38470 -860
rect 38230 -900 38470 -880
rect 38230 -970 38260 -900
rect 38260 -970 38280 -900
rect 38280 -970 38350 -900
rect 38350 -970 38370 -900
rect 38370 -970 38440 -900
rect 38440 -970 38470 -900
rect 38230 -990 38470 -970
rect 38230 -1060 38260 -990
rect 38260 -1060 38280 -990
rect 38280 -1060 38350 -990
rect 38350 -1060 38370 -990
rect 38370 -1060 38440 -990
rect 38440 -1060 38470 -990
rect 38230 -1080 38470 -1060
rect 38230 -1100 38260 -1080
rect 38260 -1100 38280 -1080
rect 38280 -1100 38350 -1080
rect 38350 -1100 38370 -1080
rect 38370 -1100 38440 -1080
rect 38440 -1100 38470 -1080
rect 38230 -1240 38260 -1190
rect 38260 -1240 38280 -1190
rect 38280 -1240 38350 -1190
rect 38350 -1240 38370 -1190
rect 38370 -1240 38440 -1190
rect 38440 -1240 38470 -1190
rect 38230 -1260 38470 -1240
rect 38230 -1330 38260 -1260
rect 38260 -1330 38280 -1260
rect 38280 -1330 38350 -1260
rect 38350 -1330 38370 -1260
rect 38370 -1330 38440 -1260
rect 38440 -1330 38470 -1260
rect 38230 -1350 38470 -1330
rect 38230 -1420 38260 -1350
rect 38260 -1420 38280 -1350
rect 38280 -1420 38350 -1350
rect 38350 -1420 38370 -1350
rect 38370 -1420 38440 -1350
rect 38440 -1420 38470 -1350
rect 38230 -1430 38470 -1420
rect 38230 -1530 38470 -1520
rect 38230 -1600 38260 -1530
rect 38260 -1600 38280 -1530
rect 38280 -1600 38350 -1530
rect 38350 -1600 38370 -1530
rect 38370 -1600 38440 -1530
rect 38440 -1600 38470 -1530
rect 38230 -1620 38470 -1600
rect 38230 -1690 38260 -1620
rect 38260 -1690 38280 -1620
rect 38280 -1690 38350 -1620
rect 38350 -1690 38370 -1620
rect 38370 -1690 38440 -1620
rect 38440 -1690 38470 -1620
rect 38230 -1710 38470 -1690
rect 38230 -1760 38260 -1710
rect 38260 -1760 38280 -1710
rect 38280 -1760 38350 -1710
rect 38350 -1760 38370 -1710
rect 38370 -1760 38440 -1710
rect 38440 -1760 38470 -1710
rect 38230 -1870 38260 -1850
rect 38260 -1870 38280 -1850
rect 38280 -1870 38350 -1850
rect 38350 -1870 38370 -1850
rect 38370 -1870 38440 -1850
rect 38440 -1870 38470 -1850
rect 38230 -1890 38470 -1870
rect 38230 -1960 38260 -1890
rect 38260 -1960 38280 -1890
rect 38280 -1960 38350 -1890
rect 38350 -1960 38370 -1890
rect 38370 -1960 38440 -1890
rect 38440 -1960 38470 -1890
rect 38230 -1980 38470 -1960
rect 38230 -2050 38260 -1980
rect 38260 -2050 38280 -1980
rect 38280 -2050 38350 -1980
rect 38350 -2050 38370 -1980
rect 38370 -2050 38440 -1980
rect 38440 -2050 38470 -1980
rect 38230 -2070 38470 -2050
rect 38230 -2090 38260 -2070
rect 38260 -2090 38280 -2070
rect 38280 -2090 38350 -2070
rect 38350 -2090 38370 -2070
rect 38370 -2090 38440 -2070
rect 38440 -2090 38470 -2070
rect 38230 -2230 38260 -2180
rect 38260 -2230 38280 -2180
rect 38280 -2230 38350 -2180
rect 38350 -2230 38370 -2180
rect 38370 -2230 38440 -2180
rect 38440 -2230 38470 -2180
rect 38230 -2250 38470 -2230
rect 38230 -2320 38260 -2250
rect 38260 -2320 38280 -2250
rect 38280 -2320 38350 -2250
rect 38350 -2320 38370 -2250
rect 38370 -2320 38440 -2250
rect 38440 -2320 38470 -2250
rect 38230 -2340 38470 -2320
rect 38230 -2410 38260 -2340
rect 38260 -2410 38280 -2340
rect 38280 -2410 38350 -2340
rect 38350 -2410 38370 -2340
rect 38370 -2410 38440 -2340
rect 38440 -2410 38470 -2340
rect 38230 -2420 38470 -2410
rect 38230 -2520 38470 -2510
rect 38230 -2590 38260 -2520
rect 38260 -2590 38280 -2520
rect 38280 -2590 38350 -2520
rect 38350 -2590 38370 -2520
rect 38370 -2590 38440 -2520
rect 38440 -2590 38470 -2520
rect 38230 -2610 38470 -2590
rect 38230 -2680 38260 -2610
rect 38260 -2680 38280 -2610
rect 38280 -2680 38350 -2610
rect 38350 -2680 38370 -2610
rect 38370 -2680 38440 -2610
rect 38440 -2680 38470 -2610
rect 38230 -2700 38470 -2680
rect 38230 -2750 38260 -2700
rect 38260 -2750 38280 -2700
rect 38280 -2750 38350 -2700
rect 38350 -2750 38370 -2700
rect 38370 -2750 38440 -2700
rect 38440 -2750 38470 -2700
rect 38230 -2860 38260 -2840
rect 38260 -2860 38280 -2840
rect 38280 -2860 38350 -2840
rect 38350 -2860 38370 -2840
rect 38370 -2860 38440 -2840
rect 38440 -2860 38470 -2840
rect 38230 -2880 38470 -2860
rect 38230 -2950 38260 -2880
rect 38260 -2950 38280 -2880
rect 38280 -2950 38350 -2880
rect 38350 -2950 38370 -2880
rect 38370 -2950 38440 -2880
rect 38440 -2950 38470 -2880
rect 38230 -2970 38470 -2950
rect 38230 -3040 38260 -2970
rect 38260 -3040 38280 -2970
rect 38280 -3040 38350 -2970
rect 38350 -3040 38370 -2970
rect 38370 -3040 38440 -2970
rect 38440 -3040 38470 -2970
rect 38230 -3060 38470 -3040
rect 38230 -3080 38260 -3060
rect 38260 -3080 38280 -3060
rect 38280 -3080 38350 -3060
rect 38350 -3080 38370 -3060
rect 38370 -3080 38440 -3060
rect 38440 -3080 38470 -3060
rect 38230 -3220 38260 -3170
rect 38260 -3220 38280 -3170
rect 38280 -3220 38350 -3170
rect 38350 -3220 38370 -3170
rect 38370 -3220 38440 -3170
rect 38440 -3220 38470 -3170
rect 38230 -3240 38470 -3220
rect 38230 -3310 38260 -3240
rect 38260 -3310 38280 -3240
rect 38280 -3310 38350 -3240
rect 38350 -3310 38370 -3240
rect 38370 -3310 38440 -3240
rect 38440 -3310 38470 -3240
rect 38230 -3330 38470 -3310
rect 38230 -3400 38260 -3330
rect 38260 -3400 38280 -3330
rect 38280 -3400 38350 -3330
rect 38350 -3400 38370 -3330
rect 38370 -3400 38440 -3330
rect 38440 -3400 38470 -3330
rect 38230 -3410 38470 -3400
rect 38230 -3550 38470 -3540
rect 38230 -3620 38260 -3550
rect 38260 -3620 38280 -3550
rect 38280 -3620 38350 -3550
rect 38350 -3620 38370 -3550
rect 38370 -3620 38440 -3550
rect 38440 -3620 38470 -3550
rect 38230 -3640 38470 -3620
rect 38230 -3710 38260 -3640
rect 38260 -3710 38280 -3640
rect 38280 -3710 38350 -3640
rect 38350 -3710 38370 -3640
rect 38370 -3710 38440 -3640
rect 38440 -3710 38470 -3640
rect 38230 -3730 38470 -3710
rect 38230 -3780 38260 -3730
rect 38260 -3780 38280 -3730
rect 38280 -3780 38350 -3730
rect 38350 -3780 38370 -3730
rect 38370 -3780 38440 -3730
rect 38440 -3780 38470 -3730
rect 38230 -3890 38260 -3870
rect 38260 -3890 38280 -3870
rect 38280 -3890 38350 -3870
rect 38350 -3890 38370 -3870
rect 38370 -3890 38440 -3870
rect 38440 -3890 38470 -3870
rect 38230 -3910 38470 -3890
rect 38230 -3980 38260 -3910
rect 38260 -3980 38280 -3910
rect 38280 -3980 38350 -3910
rect 38350 -3980 38370 -3910
rect 38370 -3980 38440 -3910
rect 38440 -3980 38470 -3910
rect 38230 -4000 38470 -3980
rect 38230 -4070 38260 -4000
rect 38260 -4070 38280 -4000
rect 38280 -4070 38350 -4000
rect 38350 -4070 38370 -4000
rect 38370 -4070 38440 -4000
rect 38440 -4070 38470 -4000
rect 38230 -4090 38470 -4070
rect 38230 -4110 38260 -4090
rect 38260 -4110 38280 -4090
rect 38280 -4110 38350 -4090
rect 38350 -4110 38370 -4090
rect 38370 -4110 38440 -4090
rect 38440 -4110 38470 -4090
rect 38230 -4250 38260 -4200
rect 38260 -4250 38280 -4200
rect 38280 -4250 38350 -4200
rect 38350 -4250 38370 -4200
rect 38370 -4250 38440 -4200
rect 38440 -4250 38470 -4200
rect 38230 -4270 38470 -4250
rect 38230 -4340 38260 -4270
rect 38260 -4340 38280 -4270
rect 38280 -4340 38350 -4270
rect 38350 -4340 38370 -4270
rect 38370 -4340 38440 -4270
rect 38440 -4340 38470 -4270
rect 38230 -4360 38470 -4340
rect 38230 -4430 38260 -4360
rect 38260 -4430 38280 -4360
rect 38280 -4430 38350 -4360
rect 38350 -4430 38370 -4360
rect 38370 -4430 38440 -4360
rect 38440 -4430 38470 -4360
rect 38230 -4440 38470 -4430
rect 38230 -4540 38470 -4530
rect 38230 -4610 38260 -4540
rect 38260 -4610 38280 -4540
rect 38280 -4610 38350 -4540
rect 38350 -4610 38370 -4540
rect 38370 -4610 38440 -4540
rect 38440 -4610 38470 -4540
rect 38230 -4630 38470 -4610
rect 38230 -4700 38260 -4630
rect 38260 -4700 38280 -4630
rect 38280 -4700 38350 -4630
rect 38350 -4700 38370 -4630
rect 38370 -4700 38440 -4630
rect 38440 -4700 38470 -4630
rect 38230 -4720 38470 -4700
rect 38230 -4770 38260 -4720
rect 38260 -4770 38280 -4720
rect 38280 -4770 38350 -4720
rect 38350 -4770 38370 -4720
rect 38370 -4770 38440 -4720
rect 38440 -4770 38470 -4720
rect 38230 -4880 38260 -4860
rect 38260 -4880 38280 -4860
rect 38280 -4880 38350 -4860
rect 38350 -4880 38370 -4860
rect 38370 -4880 38440 -4860
rect 38440 -4880 38470 -4860
rect 38230 -4900 38470 -4880
rect 38230 -4970 38260 -4900
rect 38260 -4970 38280 -4900
rect 38280 -4970 38350 -4900
rect 38350 -4970 38370 -4900
rect 38370 -4970 38440 -4900
rect 38440 -4970 38470 -4900
rect 38230 -4990 38470 -4970
rect 38230 -5060 38260 -4990
rect 38260 -5060 38280 -4990
rect 38280 -5060 38350 -4990
rect 38350 -5060 38370 -4990
rect 38370 -5060 38440 -4990
rect 38440 -5060 38470 -4990
rect 38230 -5080 38470 -5060
rect 38230 -5100 38260 -5080
rect 38260 -5100 38280 -5080
rect 38280 -5100 38350 -5080
rect 38350 -5100 38370 -5080
rect 38370 -5100 38440 -5080
rect 38440 -5100 38470 -5080
rect 38230 -5240 38260 -5190
rect 38260 -5240 38280 -5190
rect 38280 -5240 38350 -5190
rect 38350 -5240 38370 -5190
rect 38370 -5240 38440 -5190
rect 38440 -5240 38470 -5190
rect 38230 -5260 38470 -5240
rect 38230 -5330 38260 -5260
rect 38260 -5330 38280 -5260
rect 38280 -5330 38350 -5260
rect 38350 -5330 38370 -5260
rect 38370 -5330 38440 -5260
rect 38440 -5330 38470 -5260
rect 38230 -5350 38470 -5330
rect 38230 -5420 38260 -5350
rect 38260 -5420 38280 -5350
rect 38280 -5420 38350 -5350
rect 38350 -5420 38370 -5350
rect 38370 -5420 38440 -5350
rect 38440 -5420 38470 -5350
rect 38230 -5430 38470 -5420
rect 38230 -5530 38470 -5520
rect 38230 -5600 38260 -5530
rect 38260 -5600 38280 -5530
rect 38280 -5600 38350 -5530
rect 38350 -5600 38370 -5530
rect 38370 -5600 38440 -5530
rect 38440 -5600 38470 -5530
rect 38230 -5620 38470 -5600
rect 38230 -5690 38260 -5620
rect 38260 -5690 38280 -5620
rect 38280 -5690 38350 -5620
rect 38350 -5690 38370 -5620
rect 38370 -5690 38440 -5620
rect 38440 -5690 38470 -5620
rect 38230 -5710 38470 -5690
rect 38230 -5760 38260 -5710
rect 38260 -5760 38280 -5710
rect 38280 -5760 38350 -5710
rect 38350 -5760 38370 -5710
rect 38370 -5760 38440 -5710
rect 38440 -5760 38470 -5710
rect 38230 -5870 38260 -5850
rect 38260 -5870 38280 -5850
rect 38280 -5870 38350 -5850
rect 38350 -5870 38370 -5850
rect 38370 -5870 38440 -5850
rect 38440 -5870 38470 -5850
rect 38230 -5890 38470 -5870
rect 38230 -5960 38260 -5890
rect 38260 -5960 38280 -5890
rect 38280 -5960 38350 -5890
rect 38350 -5960 38370 -5890
rect 38370 -5960 38440 -5890
rect 38440 -5960 38470 -5890
rect 38230 -5980 38470 -5960
rect 38230 -6050 38260 -5980
rect 38260 -6050 38280 -5980
rect 38280 -6050 38350 -5980
rect 38350 -6050 38370 -5980
rect 38370 -6050 38440 -5980
rect 38440 -6050 38470 -5980
rect 38230 -6070 38470 -6050
rect 38230 -6090 38260 -6070
rect 38260 -6090 38280 -6070
rect 38280 -6090 38350 -6070
rect 38350 -6090 38370 -6070
rect 38370 -6090 38440 -6070
rect 38440 -6090 38470 -6070
rect 38230 -6230 38260 -6180
rect 38260 -6230 38280 -6180
rect 38280 -6230 38350 -6180
rect 38350 -6230 38370 -6180
rect 38370 -6230 38440 -6180
rect 38440 -6230 38470 -6180
rect 38230 -6250 38470 -6230
rect 38230 -6320 38260 -6250
rect 38260 -6320 38280 -6250
rect 38280 -6320 38350 -6250
rect 38350 -6320 38370 -6250
rect 38370 -6320 38440 -6250
rect 38440 -6320 38470 -6250
rect 38230 -6340 38470 -6320
rect 38230 -6410 38260 -6340
rect 38260 -6410 38280 -6340
rect 38280 -6410 38350 -6340
rect 38350 -6410 38370 -6340
rect 38370 -6410 38440 -6340
rect 38440 -6410 38470 -6340
rect 38230 -6420 38470 -6410
rect 2390 -12300 2630 -12240
rect 2720 -12300 2960 -12240
rect 3060 -12300 3300 -12240
rect 3390 -12300 3630 -12240
rect 2390 -12370 2420 -12300
rect 2420 -12370 2460 -12300
rect 2460 -12370 2530 -12300
rect 2530 -12370 2570 -12300
rect 2570 -12370 2630 -12300
rect 2720 -12370 2750 -12300
rect 2750 -12370 2790 -12300
rect 2790 -12370 2860 -12300
rect 2860 -12370 2900 -12300
rect 2900 -12370 2960 -12300
rect 3060 -12370 3080 -12300
rect 3080 -12370 3120 -12300
rect 3120 -12370 3190 -12300
rect 3190 -12370 3230 -12300
rect 3230 -12370 3300 -12300
rect 3390 -12370 3410 -12300
rect 3410 -12370 3450 -12300
rect 3450 -12370 3520 -12300
rect 3520 -12370 3560 -12300
rect 3560 -12370 3630 -12300
rect 2390 -12410 2630 -12370
rect 2720 -12410 2960 -12370
rect 3060 -12410 3300 -12370
rect 3390 -12410 3630 -12370
rect 2390 -12480 2420 -12410
rect 2420 -12480 2460 -12410
rect 2460 -12480 2530 -12410
rect 2530 -12480 2570 -12410
rect 2570 -12480 2630 -12410
rect 2720 -12480 2750 -12410
rect 2750 -12480 2790 -12410
rect 2790 -12480 2860 -12410
rect 2860 -12480 2900 -12410
rect 2900 -12480 2960 -12410
rect 3060 -12480 3080 -12410
rect 3080 -12480 3120 -12410
rect 3120 -12480 3190 -12410
rect 3190 -12480 3230 -12410
rect 3230 -12480 3300 -12410
rect 3390 -12480 3410 -12410
rect 3410 -12480 3450 -12410
rect 3450 -12480 3520 -12410
rect 3520 -12480 3560 -12410
rect 3560 -12480 3630 -12410
rect 11270 -12300 11510 -12240
rect 11600 -12300 11840 -12240
rect 11940 -12300 12180 -12240
rect 12270 -12300 12510 -12240
rect 11270 -12370 11300 -12300
rect 11300 -12370 11340 -12300
rect 11340 -12370 11410 -12300
rect 11410 -12370 11450 -12300
rect 11450 -12370 11510 -12300
rect 11600 -12370 11630 -12300
rect 11630 -12370 11670 -12300
rect 11670 -12370 11740 -12300
rect 11740 -12370 11780 -12300
rect 11780 -12370 11840 -12300
rect 11940 -12370 11960 -12300
rect 11960 -12370 12000 -12300
rect 12000 -12370 12070 -12300
rect 12070 -12370 12110 -12300
rect 12110 -12370 12180 -12300
rect 12270 -12370 12290 -12300
rect 12290 -12370 12330 -12300
rect 12330 -12370 12400 -12300
rect 12400 -12370 12440 -12300
rect 12440 -12370 12510 -12300
rect 11270 -12410 11510 -12370
rect 11600 -12410 11840 -12370
rect 11940 -12410 12180 -12370
rect 12270 -12410 12510 -12370
rect 11270 -12480 11300 -12410
rect 11300 -12480 11340 -12410
rect 11340 -12480 11410 -12410
rect 11410 -12480 11450 -12410
rect 11450 -12480 11510 -12410
rect 11600 -12480 11630 -12410
rect 11630 -12480 11670 -12410
rect 11670 -12480 11740 -12410
rect 11740 -12480 11780 -12410
rect 11780 -12480 11840 -12410
rect 11940 -12480 11960 -12410
rect 11960 -12480 12000 -12410
rect 12000 -12480 12070 -12410
rect 12070 -12480 12110 -12410
rect 12110 -12480 12180 -12410
rect 12270 -12480 12290 -12410
rect 12290 -12480 12330 -12410
rect 12330 -12480 12400 -12410
rect 12400 -12480 12440 -12410
rect 12440 -12480 12510 -12410
rect 21650 -14090 21700 -14030
rect 21700 -14090 21730 -14030
rect 21730 -14090 21800 -14030
rect 21800 -14090 21830 -14030
rect 21830 -14090 21890 -14030
rect 21650 -14120 21890 -14090
rect 21650 -14190 21700 -14120
rect 21700 -14190 21730 -14120
rect 21730 -14190 21800 -14120
rect 21800 -14190 21830 -14120
rect 21830 -14190 21890 -14120
rect 21650 -14220 21890 -14190
rect 21650 -14270 21700 -14220
rect 21700 -14270 21730 -14220
rect 21730 -14270 21800 -14220
rect 21800 -14270 21830 -14220
rect 21830 -14270 21890 -14220
rect 21650 -20170 21700 -20110
rect 21700 -20170 21730 -20110
rect 21730 -20170 21800 -20110
rect 21800 -20170 21830 -20110
rect 21830 -20170 21890 -20110
rect 21650 -20200 21890 -20170
rect 21650 -20270 21700 -20200
rect 21700 -20270 21730 -20200
rect 21730 -20270 21800 -20200
rect 21800 -20270 21830 -20200
rect 21830 -20270 21890 -20200
rect 21650 -20300 21890 -20270
rect 21650 -20350 21700 -20300
rect 21700 -20350 21730 -20300
rect 21730 -20350 21800 -20300
rect 21800 -20350 21830 -20300
rect 21830 -20350 21890 -20300
rect 2390 -22730 2460 -22660
rect 2460 -22730 2500 -22660
rect 2500 -22730 2570 -22660
rect 2570 -22730 2610 -22660
rect 2610 -22730 2630 -22660
rect 2720 -22730 2790 -22660
rect 2790 -22730 2830 -22660
rect 2830 -22730 2900 -22660
rect 2900 -22730 2940 -22660
rect 2940 -22730 2960 -22660
rect 3060 -22730 3120 -22660
rect 3120 -22730 3160 -22660
rect 3160 -22730 3230 -22660
rect 3230 -22730 3270 -22660
rect 3270 -22730 3300 -22660
rect 3390 -22730 3450 -22660
rect 3450 -22730 3490 -22660
rect 3490 -22730 3560 -22660
rect 3560 -22730 3600 -22660
rect 3600 -22730 3630 -22660
rect 2390 -22770 2630 -22730
rect 2720 -22770 2960 -22730
rect 3060 -22770 3300 -22730
rect 3390 -22770 3630 -22730
rect 2390 -22840 2460 -22770
rect 2460 -22840 2500 -22770
rect 2500 -22840 2570 -22770
rect 2570 -22840 2610 -22770
rect 2610 -22840 2630 -22770
rect 2720 -22840 2790 -22770
rect 2790 -22840 2830 -22770
rect 2830 -22840 2900 -22770
rect 2900 -22840 2940 -22770
rect 2940 -22840 2960 -22770
rect 3060 -22840 3120 -22770
rect 3120 -22840 3160 -22770
rect 3160 -22840 3230 -22770
rect 3230 -22840 3270 -22770
rect 3270 -22840 3300 -22770
rect 3390 -22840 3450 -22770
rect 3450 -22840 3490 -22770
rect 3490 -22840 3560 -22770
rect 3560 -22840 3600 -22770
rect 3600 -22840 3630 -22770
rect 2390 -22900 2630 -22840
rect 2720 -22900 2960 -22840
rect 3060 -22900 3300 -22840
rect 3390 -22900 3630 -22840
rect 11270 -22730 11340 -22660
rect 11340 -22730 11380 -22660
rect 11380 -22730 11450 -22660
rect 11450 -22730 11490 -22660
rect 11490 -22730 11510 -22660
rect 11600 -22730 11670 -22660
rect 11670 -22730 11710 -22660
rect 11710 -22730 11780 -22660
rect 11780 -22730 11820 -22660
rect 11820 -22730 11840 -22660
rect 11940 -22730 12000 -22660
rect 12000 -22730 12040 -22660
rect 12040 -22730 12110 -22660
rect 12110 -22730 12150 -22660
rect 12150 -22730 12180 -22660
rect 12270 -22730 12330 -22660
rect 12330 -22730 12370 -22660
rect 12370 -22730 12440 -22660
rect 12440 -22730 12480 -22660
rect 12480 -22730 12510 -22660
rect 11270 -22770 11510 -22730
rect 11600 -22770 11840 -22730
rect 11940 -22770 12180 -22730
rect 12270 -22770 12510 -22730
rect 11270 -22840 11340 -22770
rect 11340 -22840 11380 -22770
rect 11380 -22840 11450 -22770
rect 11450 -22840 11490 -22770
rect 11490 -22840 11510 -22770
rect 11600 -22840 11670 -22770
rect 11670 -22840 11710 -22770
rect 11710 -22840 11780 -22770
rect 11780 -22840 11820 -22770
rect 11820 -22840 11840 -22770
rect 11940 -22840 12000 -22770
rect 12000 -22840 12040 -22770
rect 12040 -22840 12110 -22770
rect 12110 -22840 12150 -22770
rect 12150 -22840 12180 -22770
rect 12270 -22840 12330 -22770
rect 12330 -22840 12370 -22770
rect 12370 -22840 12440 -22770
rect 12440 -22840 12480 -22770
rect 12480 -22840 12510 -22770
rect 11270 -22900 11510 -22840
rect 11600 -22900 11840 -22840
rect 11940 -22900 12180 -22840
rect 12270 -22900 12510 -22840
<< mimcap2 >>
rect -4980 20830 7260 20960
rect -4980 20590 -4670 20830
rect -4430 20590 -4340 20830
rect -4100 20590 -4010 20830
rect -3770 20590 -3680 20830
rect -3440 20590 -3350 20830
rect -3110 20590 -3020 20830
rect -2780 20590 -2690 20830
rect -2450 20590 -2360 20830
rect -2120 20590 -2030 20830
rect -1790 20590 -1700 20830
rect -1460 20590 -1370 20830
rect -1130 20590 -1040 20830
rect -800 20590 -710 20830
rect -470 20590 -380 20830
rect -140 20590 -50 20830
rect 190 20590 280 20830
rect 520 20590 610 20830
rect 850 20590 940 20830
rect 1180 20590 1270 20830
rect 1510 20590 1600 20830
rect 1840 20590 1930 20830
rect 2170 20590 2260 20830
rect 2500 20590 2590 20830
rect 2830 20590 2920 20830
rect 3160 20590 3250 20830
rect 3490 20590 3580 20830
rect 3820 20590 3910 20830
rect 4150 20590 4240 20830
rect 4480 20590 4570 20830
rect 4810 20590 4900 20830
rect 5140 20590 5230 20830
rect 5470 20590 5560 20830
rect 5800 20590 5890 20830
rect 6130 20590 6220 20830
rect 6460 20590 6550 20830
rect 6790 20590 6880 20830
rect 7120 20590 7260 20830
rect -4980 20500 7260 20590
rect -4980 20260 -4670 20500
rect -4430 20260 -4340 20500
rect -4100 20260 -4010 20500
rect -3770 20260 -3680 20500
rect -3440 20260 -3350 20500
rect -3110 20260 -3020 20500
rect -2780 20260 -2690 20500
rect -2450 20260 -2360 20500
rect -2120 20260 -2030 20500
rect -1790 20260 -1700 20500
rect -1460 20260 -1370 20500
rect -1130 20260 -1040 20500
rect -800 20260 -710 20500
rect -470 20260 -380 20500
rect -140 20260 -50 20500
rect 190 20260 280 20500
rect 520 20260 610 20500
rect 850 20260 940 20500
rect 1180 20260 1270 20500
rect 1510 20260 1600 20500
rect 1840 20260 1930 20500
rect 2170 20260 2260 20500
rect 2500 20260 2590 20500
rect 2830 20260 2920 20500
rect 3160 20260 3250 20500
rect 3490 20260 3580 20500
rect 3820 20260 3910 20500
rect 4150 20260 4240 20500
rect 4480 20260 4570 20500
rect 4810 20260 4900 20500
rect 5140 20260 5230 20500
rect 5470 20260 5560 20500
rect 5800 20260 5890 20500
rect 6130 20260 6220 20500
rect 6460 20260 6550 20500
rect 6790 20260 6880 20500
rect 7120 20260 7260 20500
rect -4980 20170 7260 20260
rect -4980 19930 -4670 20170
rect -4430 19930 -4340 20170
rect -4100 19930 -4010 20170
rect -3770 19930 -3680 20170
rect -3440 19930 -3350 20170
rect -3110 19930 -3020 20170
rect -2780 19930 -2690 20170
rect -2450 19930 -2360 20170
rect -2120 19930 -2030 20170
rect -1790 19930 -1700 20170
rect -1460 19930 -1370 20170
rect -1130 19930 -1040 20170
rect -800 19930 -710 20170
rect -470 19930 -380 20170
rect -140 19930 -50 20170
rect 190 19930 280 20170
rect 520 19930 610 20170
rect 850 19930 940 20170
rect 1180 19930 1270 20170
rect 1510 19930 1600 20170
rect 1840 19930 1930 20170
rect 2170 19930 2260 20170
rect 2500 19930 2590 20170
rect 2830 19930 2920 20170
rect 3160 19930 3250 20170
rect 3490 19930 3580 20170
rect 3820 19930 3910 20170
rect 4150 19930 4240 20170
rect 4480 19930 4570 20170
rect 4810 19930 4900 20170
rect 5140 19930 5230 20170
rect 5470 19930 5560 20170
rect 5800 19930 5890 20170
rect 6130 19930 6220 20170
rect 6460 19930 6550 20170
rect 6790 19930 6880 20170
rect 7120 19930 7260 20170
rect -4980 19840 7260 19930
rect -4980 19600 -4670 19840
rect -4430 19600 -4340 19840
rect -4100 19600 -4010 19840
rect -3770 19600 -3680 19840
rect -3440 19600 -3350 19840
rect -3110 19600 -3020 19840
rect -2780 19600 -2690 19840
rect -2450 19600 -2360 19840
rect -2120 19600 -2030 19840
rect -1790 19600 -1700 19840
rect -1460 19600 -1370 19840
rect -1130 19600 -1040 19840
rect -800 19600 -710 19840
rect -470 19600 -380 19840
rect -140 19600 -50 19840
rect 190 19600 280 19840
rect 520 19600 610 19840
rect 850 19600 940 19840
rect 1180 19600 1270 19840
rect 1510 19600 1600 19840
rect 1840 19600 1930 19840
rect 2170 19600 2260 19840
rect 2500 19600 2590 19840
rect 2830 19600 2920 19840
rect 3160 19600 3250 19840
rect 3490 19600 3580 19840
rect 3820 19600 3910 19840
rect 4150 19600 4240 19840
rect 4480 19600 4570 19840
rect 4810 19600 4900 19840
rect 5140 19600 5230 19840
rect 5470 19600 5560 19840
rect 5800 19600 5890 19840
rect 6130 19600 6220 19840
rect 6460 19600 6550 19840
rect 6790 19600 6880 19840
rect 7120 19600 7260 19840
rect -4980 19510 7260 19600
rect -4980 19270 -4670 19510
rect -4430 19270 -4340 19510
rect -4100 19270 -4010 19510
rect -3770 19270 -3680 19510
rect -3440 19270 -3350 19510
rect -3110 19270 -3020 19510
rect -2780 19270 -2690 19510
rect -2450 19270 -2360 19510
rect -2120 19270 -2030 19510
rect -1790 19270 -1700 19510
rect -1460 19270 -1370 19510
rect -1130 19270 -1040 19510
rect -800 19270 -710 19510
rect -470 19270 -380 19510
rect -140 19270 -50 19510
rect 190 19270 280 19510
rect 520 19270 610 19510
rect 850 19270 940 19510
rect 1180 19270 1270 19510
rect 1510 19270 1600 19510
rect 1840 19270 1930 19510
rect 2170 19270 2260 19510
rect 2500 19270 2590 19510
rect 2830 19270 2920 19510
rect 3160 19270 3250 19510
rect 3490 19270 3580 19510
rect 3820 19270 3910 19510
rect 4150 19270 4240 19510
rect 4480 19270 4570 19510
rect 4810 19270 4900 19510
rect 5140 19270 5230 19510
rect 5470 19270 5560 19510
rect 5800 19270 5890 19510
rect 6130 19270 6220 19510
rect 6460 19270 6550 19510
rect 6790 19270 6880 19510
rect 7120 19270 7260 19510
rect -4980 19180 7260 19270
rect -4980 18940 -4670 19180
rect -4430 18940 -4340 19180
rect -4100 18940 -4010 19180
rect -3770 18940 -3680 19180
rect -3440 18940 -3350 19180
rect -3110 18940 -3020 19180
rect -2780 18940 -2690 19180
rect -2450 18940 -2360 19180
rect -2120 18940 -2030 19180
rect -1790 18940 -1700 19180
rect -1460 18940 -1370 19180
rect -1130 18940 -1040 19180
rect -800 18940 -710 19180
rect -470 18940 -380 19180
rect -140 18940 -50 19180
rect 190 18940 280 19180
rect 520 18940 610 19180
rect 850 18940 940 19180
rect 1180 18940 1270 19180
rect 1510 18940 1600 19180
rect 1840 18940 1930 19180
rect 2170 18940 2260 19180
rect 2500 18940 2590 19180
rect 2830 18940 2920 19180
rect 3160 18940 3250 19180
rect 3490 18940 3580 19180
rect 3820 18940 3910 19180
rect 4150 18940 4240 19180
rect 4480 18940 4570 19180
rect 4810 18940 4900 19180
rect 5140 18940 5230 19180
rect 5470 18940 5560 19180
rect 5800 18940 5890 19180
rect 6130 18940 6220 19180
rect 6460 18940 6550 19180
rect 6790 18940 6880 19180
rect 7120 18940 7260 19180
rect -4980 18850 7260 18940
rect -4980 18610 -4670 18850
rect -4430 18610 -4340 18850
rect -4100 18610 -4010 18850
rect -3770 18610 -3680 18850
rect -3440 18610 -3350 18850
rect -3110 18610 -3020 18850
rect -2780 18610 -2690 18850
rect -2450 18610 -2360 18850
rect -2120 18610 -2030 18850
rect -1790 18610 -1700 18850
rect -1460 18610 -1370 18850
rect -1130 18610 -1040 18850
rect -800 18610 -710 18850
rect -470 18610 -380 18850
rect -140 18610 -50 18850
rect 190 18610 280 18850
rect 520 18610 610 18850
rect 850 18610 940 18850
rect 1180 18610 1270 18850
rect 1510 18610 1600 18850
rect 1840 18610 1930 18850
rect 2170 18610 2260 18850
rect 2500 18610 2590 18850
rect 2830 18610 2920 18850
rect 3160 18610 3250 18850
rect 3490 18610 3580 18850
rect 3820 18610 3910 18850
rect 4150 18610 4240 18850
rect 4480 18610 4570 18850
rect 4810 18610 4900 18850
rect 5140 18610 5230 18850
rect 5470 18610 5560 18850
rect 5800 18610 5890 18850
rect 6130 18610 6220 18850
rect 6460 18610 6550 18850
rect 6790 18610 6880 18850
rect 7120 18610 7260 18850
rect -4980 18520 7260 18610
rect -4980 18280 -4670 18520
rect -4430 18280 -4340 18520
rect -4100 18280 -4010 18520
rect -3770 18280 -3680 18520
rect -3440 18280 -3350 18520
rect -3110 18280 -3020 18520
rect -2780 18280 -2690 18520
rect -2450 18280 -2360 18520
rect -2120 18280 -2030 18520
rect -1790 18280 -1700 18520
rect -1460 18280 -1370 18520
rect -1130 18280 -1040 18520
rect -800 18280 -710 18520
rect -470 18280 -380 18520
rect -140 18280 -50 18520
rect 190 18280 280 18520
rect 520 18280 610 18520
rect 850 18280 940 18520
rect 1180 18280 1270 18520
rect 1510 18280 1600 18520
rect 1840 18280 1930 18520
rect 2170 18280 2260 18520
rect 2500 18280 2590 18520
rect 2830 18280 2920 18520
rect 3160 18280 3250 18520
rect 3490 18280 3580 18520
rect 3820 18280 3910 18520
rect 4150 18280 4240 18520
rect 4480 18280 4570 18520
rect 4810 18280 4900 18520
rect 5140 18280 5230 18520
rect 5470 18280 5560 18520
rect 5800 18280 5890 18520
rect 6130 18280 6220 18520
rect 6460 18280 6550 18520
rect 6790 18280 6880 18520
rect 7120 18280 7260 18520
rect -4980 18190 7260 18280
rect -4980 17950 -4670 18190
rect -4430 17950 -4340 18190
rect -4100 17950 -4010 18190
rect -3770 17950 -3680 18190
rect -3440 17950 -3350 18190
rect -3110 17950 -3020 18190
rect -2780 17950 -2690 18190
rect -2450 17950 -2360 18190
rect -2120 17950 -2030 18190
rect -1790 17950 -1700 18190
rect -1460 17950 -1370 18190
rect -1130 17950 -1040 18190
rect -800 17950 -710 18190
rect -470 17950 -380 18190
rect -140 17950 -50 18190
rect 190 17950 280 18190
rect 520 17950 610 18190
rect 850 17950 940 18190
rect 1180 17950 1270 18190
rect 1510 17950 1600 18190
rect 1840 17950 1930 18190
rect 2170 17950 2260 18190
rect 2500 17950 2590 18190
rect 2830 17950 2920 18190
rect 3160 17950 3250 18190
rect 3490 17950 3580 18190
rect 3820 17950 3910 18190
rect 4150 17950 4240 18190
rect 4480 17950 4570 18190
rect 4810 17950 4900 18190
rect 5140 17950 5230 18190
rect 5470 17950 5560 18190
rect 5800 17950 5890 18190
rect 6130 17950 6220 18190
rect 6460 17950 6550 18190
rect 6790 17950 6880 18190
rect 7120 17950 7260 18190
rect -4980 17860 7260 17950
rect -4980 17620 -4670 17860
rect -4430 17620 -4340 17860
rect -4100 17620 -4010 17860
rect -3770 17620 -3680 17860
rect -3440 17620 -3350 17860
rect -3110 17620 -3020 17860
rect -2780 17620 -2690 17860
rect -2450 17620 -2360 17860
rect -2120 17620 -2030 17860
rect -1790 17620 -1700 17860
rect -1460 17620 -1370 17860
rect -1130 17620 -1040 17860
rect -800 17620 -710 17860
rect -470 17620 -380 17860
rect -140 17620 -50 17860
rect 190 17620 280 17860
rect 520 17620 610 17860
rect 850 17620 940 17860
rect 1180 17620 1270 17860
rect 1510 17620 1600 17860
rect 1840 17620 1930 17860
rect 2170 17620 2260 17860
rect 2500 17620 2590 17860
rect 2830 17620 2920 17860
rect 3160 17620 3250 17860
rect 3490 17620 3580 17860
rect 3820 17620 3910 17860
rect 4150 17620 4240 17860
rect 4480 17620 4570 17860
rect 4810 17620 4900 17860
rect 5140 17620 5230 17860
rect 5470 17620 5560 17860
rect 5800 17620 5890 17860
rect 6130 17620 6220 17860
rect 6460 17620 6550 17860
rect 6790 17620 6880 17860
rect 7120 17620 7260 17860
rect -4980 17530 7260 17620
rect -4980 17290 -4670 17530
rect -4430 17290 -4340 17530
rect -4100 17290 -4010 17530
rect -3770 17290 -3680 17530
rect -3440 17290 -3350 17530
rect -3110 17290 -3020 17530
rect -2780 17290 -2690 17530
rect -2450 17290 -2360 17530
rect -2120 17290 -2030 17530
rect -1790 17290 -1700 17530
rect -1460 17290 -1370 17530
rect -1130 17290 -1040 17530
rect -800 17290 -710 17530
rect -470 17290 -380 17530
rect -140 17290 -50 17530
rect 190 17290 280 17530
rect 520 17290 610 17530
rect 850 17290 940 17530
rect 1180 17290 1270 17530
rect 1510 17290 1600 17530
rect 1840 17290 1930 17530
rect 2170 17290 2260 17530
rect 2500 17290 2590 17530
rect 2830 17290 2920 17530
rect 3160 17290 3250 17530
rect 3490 17290 3580 17530
rect 3820 17290 3910 17530
rect 4150 17290 4240 17530
rect 4480 17290 4570 17530
rect 4810 17290 4900 17530
rect 5140 17290 5230 17530
rect 5470 17290 5560 17530
rect 5800 17290 5890 17530
rect 6130 17290 6220 17530
rect 6460 17290 6550 17530
rect 6790 17290 6880 17530
rect 7120 17290 7260 17530
rect -4980 17200 7260 17290
rect -4980 16960 -4670 17200
rect -4430 16960 -4340 17200
rect -4100 16960 -4010 17200
rect -3770 16960 -3680 17200
rect -3440 16960 -3350 17200
rect -3110 16960 -3020 17200
rect -2780 16960 -2690 17200
rect -2450 16960 -2360 17200
rect -2120 16960 -2030 17200
rect -1790 16960 -1700 17200
rect -1460 16960 -1370 17200
rect -1130 16960 -1040 17200
rect -800 16960 -710 17200
rect -470 16960 -380 17200
rect -140 16960 -50 17200
rect 190 16960 280 17200
rect 520 16960 610 17200
rect 850 16960 940 17200
rect 1180 16960 1270 17200
rect 1510 16960 1600 17200
rect 1840 16960 1930 17200
rect 2170 16960 2260 17200
rect 2500 16960 2590 17200
rect 2830 16960 2920 17200
rect 3160 16960 3250 17200
rect 3490 16960 3580 17200
rect 3820 16960 3910 17200
rect 4150 16960 4240 17200
rect 4480 16960 4570 17200
rect 4810 16960 4900 17200
rect 5140 16960 5230 17200
rect 5470 16960 5560 17200
rect 5800 16960 5890 17200
rect 6130 16960 6220 17200
rect 6460 16960 6550 17200
rect 6790 16960 6880 17200
rect 7120 16960 7260 17200
rect -4980 16870 7260 16960
rect -4980 16630 -4670 16870
rect -4430 16630 -4340 16870
rect -4100 16630 -4010 16870
rect -3770 16630 -3680 16870
rect -3440 16630 -3350 16870
rect -3110 16630 -3020 16870
rect -2780 16630 -2690 16870
rect -2450 16630 -2360 16870
rect -2120 16630 -2030 16870
rect -1790 16630 -1700 16870
rect -1460 16630 -1370 16870
rect -1130 16630 -1040 16870
rect -800 16630 -710 16870
rect -470 16630 -380 16870
rect -140 16630 -50 16870
rect 190 16630 280 16870
rect 520 16630 610 16870
rect 850 16630 940 16870
rect 1180 16630 1270 16870
rect 1510 16630 1600 16870
rect 1840 16630 1930 16870
rect 2170 16630 2260 16870
rect 2500 16630 2590 16870
rect 2830 16630 2920 16870
rect 3160 16630 3250 16870
rect 3490 16630 3580 16870
rect 3820 16630 3910 16870
rect 4150 16630 4240 16870
rect 4480 16630 4570 16870
rect 4810 16630 4900 16870
rect 5140 16630 5230 16870
rect 5470 16630 5560 16870
rect 5800 16630 5890 16870
rect 6130 16630 6220 16870
rect 6460 16630 6550 16870
rect 6790 16630 6880 16870
rect 7120 16630 7260 16870
rect -4980 16540 7260 16630
rect -4980 16300 -4670 16540
rect -4430 16300 -4340 16540
rect -4100 16300 -4010 16540
rect -3770 16300 -3680 16540
rect -3440 16300 -3350 16540
rect -3110 16300 -3020 16540
rect -2780 16300 -2690 16540
rect -2450 16300 -2360 16540
rect -2120 16300 -2030 16540
rect -1790 16300 -1700 16540
rect -1460 16300 -1370 16540
rect -1130 16300 -1040 16540
rect -800 16300 -710 16540
rect -470 16300 -380 16540
rect -140 16300 -50 16540
rect 190 16300 280 16540
rect 520 16300 610 16540
rect 850 16300 940 16540
rect 1180 16300 1270 16540
rect 1510 16300 1600 16540
rect 1840 16300 1930 16540
rect 2170 16300 2260 16540
rect 2500 16300 2590 16540
rect 2830 16300 2920 16540
rect 3160 16300 3250 16540
rect 3490 16300 3580 16540
rect 3820 16300 3910 16540
rect 4150 16300 4240 16540
rect 4480 16300 4570 16540
rect 4810 16300 4900 16540
rect 5140 16300 5230 16540
rect 5470 16300 5560 16540
rect 5800 16300 5890 16540
rect 6130 16300 6220 16540
rect 6460 16300 6550 16540
rect 6790 16300 6880 16540
rect 7120 16300 7260 16540
rect -4980 16210 7260 16300
rect -4980 15970 -4670 16210
rect -4430 15970 -4340 16210
rect -4100 15970 -4010 16210
rect -3770 15970 -3680 16210
rect -3440 15970 -3350 16210
rect -3110 15970 -3020 16210
rect -2780 15970 -2690 16210
rect -2450 15970 -2360 16210
rect -2120 15970 -2030 16210
rect -1790 15970 -1700 16210
rect -1460 15970 -1370 16210
rect -1130 15970 -1040 16210
rect -800 15970 -710 16210
rect -470 15970 -380 16210
rect -140 15970 -50 16210
rect 190 15970 280 16210
rect 520 15970 610 16210
rect 850 15970 940 16210
rect 1180 15970 1270 16210
rect 1510 15970 1600 16210
rect 1840 15970 1930 16210
rect 2170 15970 2260 16210
rect 2500 15970 2590 16210
rect 2830 15970 2920 16210
rect 3160 15970 3250 16210
rect 3490 15970 3580 16210
rect 3820 15970 3910 16210
rect 4150 15970 4240 16210
rect 4480 15970 4570 16210
rect 4810 15970 4900 16210
rect 5140 15970 5230 16210
rect 5470 15970 5560 16210
rect 5800 15970 5890 16210
rect 6130 15970 6220 16210
rect 6460 15970 6550 16210
rect 6790 15970 6880 16210
rect 7120 15970 7260 16210
rect -4980 15880 7260 15970
rect -4980 15640 -4670 15880
rect -4430 15640 -4340 15880
rect -4100 15640 -4010 15880
rect -3770 15640 -3680 15880
rect -3440 15640 -3350 15880
rect -3110 15640 -3020 15880
rect -2780 15640 -2690 15880
rect -2450 15640 -2360 15880
rect -2120 15640 -2030 15880
rect -1790 15640 -1700 15880
rect -1460 15640 -1370 15880
rect -1130 15640 -1040 15880
rect -800 15640 -710 15880
rect -470 15640 -380 15880
rect -140 15640 -50 15880
rect 190 15640 280 15880
rect 520 15640 610 15880
rect 850 15640 940 15880
rect 1180 15640 1270 15880
rect 1510 15640 1600 15880
rect 1840 15640 1930 15880
rect 2170 15640 2260 15880
rect 2500 15640 2590 15880
rect 2830 15640 2920 15880
rect 3160 15640 3250 15880
rect 3490 15640 3580 15880
rect 3820 15640 3910 15880
rect 4150 15640 4240 15880
rect 4480 15640 4570 15880
rect 4810 15640 4900 15880
rect 5140 15640 5230 15880
rect 5470 15640 5560 15880
rect 5800 15640 5890 15880
rect 6130 15640 6220 15880
rect 6460 15640 6550 15880
rect 6790 15640 6880 15880
rect 7120 15640 7260 15880
rect -4980 15550 7260 15640
rect -4980 15310 -4670 15550
rect -4430 15310 -4340 15550
rect -4100 15310 -4010 15550
rect -3770 15310 -3680 15550
rect -3440 15310 -3350 15550
rect -3110 15310 -3020 15550
rect -2780 15310 -2690 15550
rect -2450 15310 -2360 15550
rect -2120 15310 -2030 15550
rect -1790 15310 -1700 15550
rect -1460 15310 -1370 15550
rect -1130 15310 -1040 15550
rect -800 15310 -710 15550
rect -470 15310 -380 15550
rect -140 15310 -50 15550
rect 190 15310 280 15550
rect 520 15310 610 15550
rect 850 15310 940 15550
rect 1180 15310 1270 15550
rect 1510 15310 1600 15550
rect 1840 15310 1930 15550
rect 2170 15310 2260 15550
rect 2500 15310 2590 15550
rect 2830 15310 2920 15550
rect 3160 15310 3250 15550
rect 3490 15310 3580 15550
rect 3820 15310 3910 15550
rect 4150 15310 4240 15550
rect 4480 15310 4570 15550
rect 4810 15310 4900 15550
rect 5140 15310 5230 15550
rect 5470 15310 5560 15550
rect 5800 15310 5890 15550
rect 6130 15310 6220 15550
rect 6460 15310 6550 15550
rect 6790 15310 6880 15550
rect 7120 15310 7260 15550
rect -4980 15220 7260 15310
rect -4980 14980 -4670 15220
rect -4430 14980 -4340 15220
rect -4100 14980 -4010 15220
rect -3770 14980 -3680 15220
rect -3440 14980 -3350 15220
rect -3110 14980 -3020 15220
rect -2780 14980 -2690 15220
rect -2450 14980 -2360 15220
rect -2120 14980 -2030 15220
rect -1790 14980 -1700 15220
rect -1460 14980 -1370 15220
rect -1130 14980 -1040 15220
rect -800 14980 -710 15220
rect -470 14980 -380 15220
rect -140 14980 -50 15220
rect 190 14980 280 15220
rect 520 14980 610 15220
rect 850 14980 940 15220
rect 1180 14980 1270 15220
rect 1510 14980 1600 15220
rect 1840 14980 1930 15220
rect 2170 14980 2260 15220
rect 2500 14980 2590 15220
rect 2830 14980 2920 15220
rect 3160 14980 3250 15220
rect 3490 14980 3580 15220
rect 3820 14980 3910 15220
rect 4150 14980 4240 15220
rect 4480 14980 4570 15220
rect 4810 14980 4900 15220
rect 5140 14980 5230 15220
rect 5470 14980 5560 15220
rect 5800 14980 5890 15220
rect 6130 14980 6220 15220
rect 6460 14980 6550 15220
rect 6790 14980 6880 15220
rect 7120 14980 7260 15220
rect -4980 14890 7260 14980
rect -4980 14650 -4670 14890
rect -4430 14650 -4340 14890
rect -4100 14650 -4010 14890
rect -3770 14650 -3680 14890
rect -3440 14650 -3350 14890
rect -3110 14650 -3020 14890
rect -2780 14650 -2690 14890
rect -2450 14650 -2360 14890
rect -2120 14650 -2030 14890
rect -1790 14650 -1700 14890
rect -1460 14650 -1370 14890
rect -1130 14650 -1040 14890
rect -800 14650 -710 14890
rect -470 14650 -380 14890
rect -140 14650 -50 14890
rect 190 14650 280 14890
rect 520 14650 610 14890
rect 850 14650 940 14890
rect 1180 14650 1270 14890
rect 1510 14650 1600 14890
rect 1840 14650 1930 14890
rect 2170 14650 2260 14890
rect 2500 14650 2590 14890
rect 2830 14650 2920 14890
rect 3160 14650 3250 14890
rect 3490 14650 3580 14890
rect 3820 14650 3910 14890
rect 4150 14650 4240 14890
rect 4480 14650 4570 14890
rect 4810 14650 4900 14890
rect 5140 14650 5230 14890
rect 5470 14650 5560 14890
rect 5800 14650 5890 14890
rect 6130 14650 6220 14890
rect 6460 14650 6550 14890
rect 6790 14650 6880 14890
rect 7120 14650 7260 14890
rect -4980 14560 7260 14650
rect -4980 14320 -4670 14560
rect -4430 14320 -4340 14560
rect -4100 14320 -4010 14560
rect -3770 14320 -3680 14560
rect -3440 14320 -3350 14560
rect -3110 14320 -3020 14560
rect -2780 14320 -2690 14560
rect -2450 14320 -2360 14560
rect -2120 14320 -2030 14560
rect -1790 14320 -1700 14560
rect -1460 14320 -1370 14560
rect -1130 14320 -1040 14560
rect -800 14320 -710 14560
rect -470 14320 -380 14560
rect -140 14320 -50 14560
rect 190 14320 280 14560
rect 520 14320 610 14560
rect 850 14320 940 14560
rect 1180 14320 1270 14560
rect 1510 14320 1600 14560
rect 1840 14320 1930 14560
rect 2170 14320 2260 14560
rect 2500 14320 2590 14560
rect 2830 14320 2920 14560
rect 3160 14320 3250 14560
rect 3490 14320 3580 14560
rect 3820 14320 3910 14560
rect 4150 14320 4240 14560
rect 4480 14320 4570 14560
rect 4810 14320 4900 14560
rect 5140 14320 5230 14560
rect 5470 14320 5560 14560
rect 5800 14320 5890 14560
rect 6130 14320 6220 14560
rect 6460 14320 6550 14560
rect 6790 14320 6880 14560
rect 7120 14320 7260 14560
rect -4980 14230 7260 14320
rect -4980 13990 -4670 14230
rect -4430 13990 -4340 14230
rect -4100 13990 -4010 14230
rect -3770 13990 -3680 14230
rect -3440 13990 -3350 14230
rect -3110 13990 -3020 14230
rect -2780 13990 -2690 14230
rect -2450 13990 -2360 14230
rect -2120 13990 -2030 14230
rect -1790 13990 -1700 14230
rect -1460 13990 -1370 14230
rect -1130 13990 -1040 14230
rect -800 13990 -710 14230
rect -470 13990 -380 14230
rect -140 13990 -50 14230
rect 190 13990 280 14230
rect 520 13990 610 14230
rect 850 13990 940 14230
rect 1180 13990 1270 14230
rect 1510 13990 1600 14230
rect 1840 13990 1930 14230
rect 2170 13990 2260 14230
rect 2500 13990 2590 14230
rect 2830 13990 2920 14230
rect 3160 13990 3250 14230
rect 3490 13990 3580 14230
rect 3820 13990 3910 14230
rect 4150 13990 4240 14230
rect 4480 13990 4570 14230
rect 4810 13990 4900 14230
rect 5140 13990 5230 14230
rect 5470 13990 5560 14230
rect 5800 13990 5890 14230
rect 6130 13990 6220 14230
rect 6460 13990 6550 14230
rect 6790 13990 6880 14230
rect 7120 13990 7260 14230
rect -4980 13900 7260 13990
rect -4980 13660 -4670 13900
rect -4430 13660 -4340 13900
rect -4100 13660 -4010 13900
rect -3770 13660 -3680 13900
rect -3440 13660 -3350 13900
rect -3110 13660 -3020 13900
rect -2780 13660 -2690 13900
rect -2450 13660 -2360 13900
rect -2120 13660 -2030 13900
rect -1790 13660 -1700 13900
rect -1460 13660 -1370 13900
rect -1130 13660 -1040 13900
rect -800 13660 -710 13900
rect -470 13660 -380 13900
rect -140 13660 -50 13900
rect 190 13660 280 13900
rect 520 13660 610 13900
rect 850 13660 940 13900
rect 1180 13660 1270 13900
rect 1510 13660 1600 13900
rect 1840 13660 1930 13900
rect 2170 13660 2260 13900
rect 2500 13660 2590 13900
rect 2830 13660 2920 13900
rect 3160 13660 3250 13900
rect 3490 13660 3580 13900
rect 3820 13660 3910 13900
rect 4150 13660 4240 13900
rect 4480 13660 4570 13900
rect 4810 13660 4900 13900
rect 5140 13660 5230 13900
rect 5470 13660 5560 13900
rect 5800 13660 5890 13900
rect 6130 13660 6220 13900
rect 6460 13660 6550 13900
rect 6790 13660 6880 13900
rect 7120 13660 7260 13900
rect -4980 13570 7260 13660
rect -4980 13330 -4670 13570
rect -4430 13330 -4340 13570
rect -4100 13330 -4010 13570
rect -3770 13330 -3680 13570
rect -3440 13330 -3350 13570
rect -3110 13330 -3020 13570
rect -2780 13330 -2690 13570
rect -2450 13330 -2360 13570
rect -2120 13330 -2030 13570
rect -1790 13330 -1700 13570
rect -1460 13330 -1370 13570
rect -1130 13330 -1040 13570
rect -800 13330 -710 13570
rect -470 13330 -380 13570
rect -140 13330 -50 13570
rect 190 13330 280 13570
rect 520 13330 610 13570
rect 850 13330 940 13570
rect 1180 13330 1270 13570
rect 1510 13330 1600 13570
rect 1840 13330 1930 13570
rect 2170 13330 2260 13570
rect 2500 13330 2590 13570
rect 2830 13330 2920 13570
rect 3160 13330 3250 13570
rect 3490 13330 3580 13570
rect 3820 13330 3910 13570
rect 4150 13330 4240 13570
rect 4480 13330 4570 13570
rect 4810 13330 4900 13570
rect 5140 13330 5230 13570
rect 5470 13330 5560 13570
rect 5800 13330 5890 13570
rect 6130 13330 6220 13570
rect 6460 13330 6550 13570
rect 6790 13330 6880 13570
rect 7120 13330 7260 13570
rect -4980 13240 7260 13330
rect -4980 13000 -4670 13240
rect -4430 13000 -4340 13240
rect -4100 13000 -4010 13240
rect -3770 13000 -3680 13240
rect -3440 13000 -3350 13240
rect -3110 13000 -3020 13240
rect -2780 13000 -2690 13240
rect -2450 13000 -2360 13240
rect -2120 13000 -2030 13240
rect -1790 13000 -1700 13240
rect -1460 13000 -1370 13240
rect -1130 13000 -1040 13240
rect -800 13000 -710 13240
rect -470 13000 -380 13240
rect -140 13000 -50 13240
rect 190 13000 280 13240
rect 520 13000 610 13240
rect 850 13000 940 13240
rect 1180 13000 1270 13240
rect 1510 13000 1600 13240
rect 1840 13000 1930 13240
rect 2170 13000 2260 13240
rect 2500 13000 2590 13240
rect 2830 13000 2920 13240
rect 3160 13000 3250 13240
rect 3490 13000 3580 13240
rect 3820 13000 3910 13240
rect 4150 13000 4240 13240
rect 4480 13000 4570 13240
rect 4810 13000 4900 13240
rect 5140 13000 5230 13240
rect 5470 13000 5560 13240
rect 5800 13000 5890 13240
rect 6130 13000 6220 13240
rect 6460 13000 6550 13240
rect 6790 13000 6880 13240
rect 7120 13000 7260 13240
rect -4980 12910 7260 13000
rect -4980 12670 -4670 12910
rect -4430 12670 -4340 12910
rect -4100 12670 -4010 12910
rect -3770 12670 -3680 12910
rect -3440 12670 -3350 12910
rect -3110 12670 -3020 12910
rect -2780 12670 -2690 12910
rect -2450 12670 -2360 12910
rect -2120 12670 -2030 12910
rect -1790 12670 -1700 12910
rect -1460 12670 -1370 12910
rect -1130 12670 -1040 12910
rect -800 12670 -710 12910
rect -470 12670 -380 12910
rect -140 12670 -50 12910
rect 190 12670 280 12910
rect 520 12670 610 12910
rect 850 12670 940 12910
rect 1180 12670 1270 12910
rect 1510 12670 1600 12910
rect 1840 12670 1930 12910
rect 2170 12670 2260 12910
rect 2500 12670 2590 12910
rect 2830 12670 2920 12910
rect 3160 12670 3250 12910
rect 3490 12670 3580 12910
rect 3820 12670 3910 12910
rect 4150 12670 4240 12910
rect 4480 12670 4570 12910
rect 4810 12670 4900 12910
rect 5140 12670 5230 12910
rect 5470 12670 5560 12910
rect 5800 12670 5890 12910
rect 6130 12670 6220 12910
rect 6460 12670 6550 12910
rect 6790 12670 6880 12910
rect 7120 12670 7260 12910
rect -4980 12580 7260 12670
rect -4980 12340 -4670 12580
rect -4430 12340 -4340 12580
rect -4100 12340 -4010 12580
rect -3770 12340 -3680 12580
rect -3440 12340 -3350 12580
rect -3110 12340 -3020 12580
rect -2780 12340 -2690 12580
rect -2450 12340 -2360 12580
rect -2120 12340 -2030 12580
rect -1790 12340 -1700 12580
rect -1460 12340 -1370 12580
rect -1130 12340 -1040 12580
rect -800 12340 -710 12580
rect -470 12340 -380 12580
rect -140 12340 -50 12580
rect 190 12340 280 12580
rect 520 12340 610 12580
rect 850 12340 940 12580
rect 1180 12340 1270 12580
rect 1510 12340 1600 12580
rect 1840 12340 1930 12580
rect 2170 12340 2260 12580
rect 2500 12340 2590 12580
rect 2830 12340 2920 12580
rect 3160 12340 3250 12580
rect 3490 12340 3580 12580
rect 3820 12340 3910 12580
rect 4150 12340 4240 12580
rect 4480 12340 4570 12580
rect 4810 12340 4900 12580
rect 5140 12340 5230 12580
rect 5470 12340 5560 12580
rect 5800 12340 5890 12580
rect 6130 12340 6220 12580
rect 6460 12340 6550 12580
rect 6790 12340 6880 12580
rect 7120 12340 7260 12580
rect -4980 12250 7260 12340
rect -4980 12010 -4670 12250
rect -4430 12010 -4340 12250
rect -4100 12010 -4010 12250
rect -3770 12010 -3680 12250
rect -3440 12010 -3350 12250
rect -3110 12010 -3020 12250
rect -2780 12010 -2690 12250
rect -2450 12010 -2360 12250
rect -2120 12010 -2030 12250
rect -1790 12010 -1700 12250
rect -1460 12010 -1370 12250
rect -1130 12010 -1040 12250
rect -800 12010 -710 12250
rect -470 12010 -380 12250
rect -140 12010 -50 12250
rect 190 12010 280 12250
rect 520 12010 610 12250
rect 850 12010 940 12250
rect 1180 12010 1270 12250
rect 1510 12010 1600 12250
rect 1840 12010 1930 12250
rect 2170 12010 2260 12250
rect 2500 12010 2590 12250
rect 2830 12010 2920 12250
rect 3160 12010 3250 12250
rect 3490 12010 3580 12250
rect 3820 12010 3910 12250
rect 4150 12010 4240 12250
rect 4480 12010 4570 12250
rect 4810 12010 4900 12250
rect 5140 12010 5230 12250
rect 5470 12010 5560 12250
rect 5800 12010 5890 12250
rect 6130 12010 6220 12250
rect 6460 12010 6550 12250
rect 6790 12010 6880 12250
rect 7120 12010 7260 12250
rect -4980 11920 7260 12010
rect -4980 11680 -4670 11920
rect -4430 11680 -4340 11920
rect -4100 11680 -4010 11920
rect -3770 11680 -3680 11920
rect -3440 11680 -3350 11920
rect -3110 11680 -3020 11920
rect -2780 11680 -2690 11920
rect -2450 11680 -2360 11920
rect -2120 11680 -2030 11920
rect -1790 11680 -1700 11920
rect -1460 11680 -1370 11920
rect -1130 11680 -1040 11920
rect -800 11680 -710 11920
rect -470 11680 -380 11920
rect -140 11680 -50 11920
rect 190 11680 280 11920
rect 520 11680 610 11920
rect 850 11680 940 11920
rect 1180 11680 1270 11920
rect 1510 11680 1600 11920
rect 1840 11680 1930 11920
rect 2170 11680 2260 11920
rect 2500 11680 2590 11920
rect 2830 11680 2920 11920
rect 3160 11680 3250 11920
rect 3490 11680 3580 11920
rect 3820 11680 3910 11920
rect 4150 11680 4240 11920
rect 4480 11680 4570 11920
rect 4810 11680 4900 11920
rect 5140 11680 5230 11920
rect 5470 11680 5560 11920
rect 5800 11680 5890 11920
rect 6130 11680 6220 11920
rect 6460 11680 6550 11920
rect 6790 11680 6880 11920
rect 7120 11680 7260 11920
rect -4980 11590 7260 11680
rect -4980 11350 -4670 11590
rect -4430 11350 -4340 11590
rect -4100 11350 -4010 11590
rect -3770 11350 -3680 11590
rect -3440 11350 -3350 11590
rect -3110 11350 -3020 11590
rect -2780 11350 -2690 11590
rect -2450 11350 -2360 11590
rect -2120 11350 -2030 11590
rect -1790 11350 -1700 11590
rect -1460 11350 -1370 11590
rect -1130 11350 -1040 11590
rect -800 11350 -710 11590
rect -470 11350 -380 11590
rect -140 11350 -50 11590
rect 190 11350 280 11590
rect 520 11350 610 11590
rect 850 11350 940 11590
rect 1180 11350 1270 11590
rect 1510 11350 1600 11590
rect 1840 11350 1930 11590
rect 2170 11350 2260 11590
rect 2500 11350 2590 11590
rect 2830 11350 2920 11590
rect 3160 11350 3250 11590
rect 3490 11350 3580 11590
rect 3820 11350 3910 11590
rect 4150 11350 4240 11590
rect 4480 11350 4570 11590
rect 4810 11350 4900 11590
rect 5140 11350 5230 11590
rect 5470 11350 5560 11590
rect 5800 11350 5890 11590
rect 6130 11350 6220 11590
rect 6460 11350 6550 11590
rect 6790 11350 6880 11590
rect 7120 11350 7260 11590
rect -4980 11260 7260 11350
rect -4980 11020 -4670 11260
rect -4430 11020 -4340 11260
rect -4100 11020 -4010 11260
rect -3770 11020 -3680 11260
rect -3440 11020 -3350 11260
rect -3110 11020 -3020 11260
rect -2780 11020 -2690 11260
rect -2450 11020 -2360 11260
rect -2120 11020 -2030 11260
rect -1790 11020 -1700 11260
rect -1460 11020 -1370 11260
rect -1130 11020 -1040 11260
rect -800 11020 -710 11260
rect -470 11020 -380 11260
rect -140 11020 -50 11260
rect 190 11020 280 11260
rect 520 11020 610 11260
rect 850 11020 940 11260
rect 1180 11020 1270 11260
rect 1510 11020 1600 11260
rect 1840 11020 1930 11260
rect 2170 11020 2260 11260
rect 2500 11020 2590 11260
rect 2830 11020 2920 11260
rect 3160 11020 3250 11260
rect 3490 11020 3580 11260
rect 3820 11020 3910 11260
rect 4150 11020 4240 11260
rect 4480 11020 4570 11260
rect 4810 11020 4900 11260
rect 5140 11020 5230 11260
rect 5470 11020 5560 11260
rect 5800 11020 5890 11260
rect 6130 11020 6220 11260
rect 6460 11020 6550 11260
rect 6790 11020 6880 11260
rect 7120 11020 7260 11260
rect -4980 10930 7260 11020
rect -4980 10690 -4670 10930
rect -4430 10690 -4340 10930
rect -4100 10690 -4010 10930
rect -3770 10690 -3680 10930
rect -3440 10690 -3350 10930
rect -3110 10690 -3020 10930
rect -2780 10690 -2690 10930
rect -2450 10690 -2360 10930
rect -2120 10690 -2030 10930
rect -1790 10690 -1700 10930
rect -1460 10690 -1370 10930
rect -1130 10690 -1040 10930
rect -800 10690 -710 10930
rect -470 10690 -380 10930
rect -140 10690 -50 10930
rect 190 10690 280 10930
rect 520 10690 610 10930
rect 850 10690 940 10930
rect 1180 10690 1270 10930
rect 1510 10690 1600 10930
rect 1840 10690 1930 10930
rect 2170 10690 2260 10930
rect 2500 10690 2590 10930
rect 2830 10690 2920 10930
rect 3160 10690 3250 10930
rect 3490 10690 3580 10930
rect 3820 10690 3910 10930
rect 4150 10690 4240 10930
rect 4480 10690 4570 10930
rect 4810 10690 4900 10930
rect 5140 10690 5230 10930
rect 5470 10690 5560 10930
rect 5800 10690 5890 10930
rect 6130 10690 6220 10930
rect 6460 10690 6550 10930
rect 6790 10690 6880 10930
rect 7120 10690 7260 10930
rect -4980 10600 7260 10690
rect -4980 10360 -4670 10600
rect -4430 10360 -4340 10600
rect -4100 10360 -4010 10600
rect -3770 10360 -3680 10600
rect -3440 10360 -3350 10600
rect -3110 10360 -3020 10600
rect -2780 10360 -2690 10600
rect -2450 10360 -2360 10600
rect -2120 10360 -2030 10600
rect -1790 10360 -1700 10600
rect -1460 10360 -1370 10600
rect -1130 10360 -1040 10600
rect -800 10360 -710 10600
rect -470 10360 -380 10600
rect -140 10360 -50 10600
rect 190 10360 280 10600
rect 520 10360 610 10600
rect 850 10360 940 10600
rect 1180 10360 1270 10600
rect 1510 10360 1600 10600
rect 1840 10360 1930 10600
rect 2170 10360 2260 10600
rect 2500 10360 2590 10600
rect 2830 10360 2920 10600
rect 3160 10360 3250 10600
rect 3490 10360 3580 10600
rect 3820 10360 3910 10600
rect 4150 10360 4240 10600
rect 4480 10360 4570 10600
rect 4810 10360 4900 10600
rect 5140 10360 5230 10600
rect 5470 10360 5560 10600
rect 5800 10360 5890 10600
rect 6130 10360 6220 10600
rect 6460 10360 6550 10600
rect 6790 10360 6880 10600
rect 7120 10360 7260 10600
rect -4980 10270 7260 10360
rect -4980 10030 -4670 10270
rect -4430 10030 -4340 10270
rect -4100 10030 -4010 10270
rect -3770 10030 -3680 10270
rect -3440 10030 -3350 10270
rect -3110 10030 -3020 10270
rect -2780 10030 -2690 10270
rect -2450 10030 -2360 10270
rect -2120 10030 -2030 10270
rect -1790 10030 -1700 10270
rect -1460 10030 -1370 10270
rect -1130 10030 -1040 10270
rect -800 10030 -710 10270
rect -470 10030 -380 10270
rect -140 10030 -50 10270
rect 190 10030 280 10270
rect 520 10030 610 10270
rect 850 10030 940 10270
rect 1180 10030 1270 10270
rect 1510 10030 1600 10270
rect 1840 10030 1930 10270
rect 2170 10030 2260 10270
rect 2500 10030 2590 10270
rect 2830 10030 2920 10270
rect 3160 10030 3250 10270
rect 3490 10030 3580 10270
rect 3820 10030 3910 10270
rect 4150 10030 4240 10270
rect 4480 10030 4570 10270
rect 4810 10030 4900 10270
rect 5140 10030 5230 10270
rect 5470 10030 5560 10270
rect 5800 10030 5890 10270
rect 6130 10030 6220 10270
rect 6460 10030 6550 10270
rect 6790 10030 6880 10270
rect 7120 10030 7260 10270
rect -4980 9940 7260 10030
rect -4980 9700 -4670 9940
rect -4430 9700 -4340 9940
rect -4100 9700 -4010 9940
rect -3770 9700 -3680 9940
rect -3440 9700 -3350 9940
rect -3110 9700 -3020 9940
rect -2780 9700 -2690 9940
rect -2450 9700 -2360 9940
rect -2120 9700 -2030 9940
rect -1790 9700 -1700 9940
rect -1460 9700 -1370 9940
rect -1130 9700 -1040 9940
rect -800 9700 -710 9940
rect -470 9700 -380 9940
rect -140 9700 -50 9940
rect 190 9700 280 9940
rect 520 9700 610 9940
rect 850 9700 940 9940
rect 1180 9700 1270 9940
rect 1510 9700 1600 9940
rect 1840 9700 1930 9940
rect 2170 9700 2260 9940
rect 2500 9700 2590 9940
rect 2830 9700 2920 9940
rect 3160 9700 3250 9940
rect 3490 9700 3580 9940
rect 3820 9700 3910 9940
rect 4150 9700 4240 9940
rect 4480 9700 4570 9940
rect 4810 9700 4900 9940
rect 5140 9700 5230 9940
rect 5470 9700 5560 9940
rect 5800 9700 5890 9940
rect 6130 9700 6220 9940
rect 6460 9700 6550 9940
rect 6790 9700 6880 9940
rect 7120 9700 7260 9940
rect -4980 9610 7260 9700
rect -4980 9370 -4670 9610
rect -4430 9370 -4340 9610
rect -4100 9370 -4010 9610
rect -3770 9370 -3680 9610
rect -3440 9370 -3350 9610
rect -3110 9370 -3020 9610
rect -2780 9370 -2690 9610
rect -2450 9370 -2360 9610
rect -2120 9370 -2030 9610
rect -1790 9370 -1700 9610
rect -1460 9370 -1370 9610
rect -1130 9370 -1040 9610
rect -800 9370 -710 9610
rect -470 9370 -380 9610
rect -140 9370 -50 9610
rect 190 9370 280 9610
rect 520 9370 610 9610
rect 850 9370 940 9610
rect 1180 9370 1270 9610
rect 1510 9370 1600 9610
rect 1840 9370 1930 9610
rect 2170 9370 2260 9610
rect 2500 9370 2590 9610
rect 2830 9370 2920 9610
rect 3160 9370 3250 9610
rect 3490 9370 3580 9610
rect 3820 9370 3910 9610
rect 4150 9370 4240 9610
rect 4480 9370 4570 9610
rect 4810 9370 4900 9610
rect 5140 9370 5230 9610
rect 5470 9370 5560 9610
rect 5800 9370 5890 9610
rect 6130 9370 6220 9610
rect 6460 9370 6550 9610
rect 6790 9370 6880 9610
rect 7120 9370 7260 9610
rect -4980 9280 7260 9370
rect -4980 9040 -4670 9280
rect -4430 9040 -4340 9280
rect -4100 9040 -4010 9280
rect -3770 9040 -3680 9280
rect -3440 9040 -3350 9280
rect -3110 9040 -3020 9280
rect -2780 9040 -2690 9280
rect -2450 9040 -2360 9280
rect -2120 9040 -2030 9280
rect -1790 9040 -1700 9280
rect -1460 9040 -1370 9280
rect -1130 9040 -1040 9280
rect -800 9040 -710 9280
rect -470 9040 -380 9280
rect -140 9040 -50 9280
rect 190 9040 280 9280
rect 520 9040 610 9280
rect 850 9040 940 9280
rect 1180 9040 1270 9280
rect 1510 9040 1600 9280
rect 1840 9040 1930 9280
rect 2170 9040 2260 9280
rect 2500 9040 2590 9280
rect 2830 9040 2920 9280
rect 3160 9040 3250 9280
rect 3490 9040 3580 9280
rect 3820 9040 3910 9280
rect 4150 9040 4240 9280
rect 4480 9040 4570 9280
rect 4810 9040 4900 9280
rect 5140 9040 5230 9280
rect 5470 9040 5560 9280
rect 5800 9040 5890 9280
rect 6130 9040 6220 9280
rect 6460 9040 6550 9280
rect 6790 9040 6880 9280
rect 7120 9040 7260 9280
rect -4980 8720 7260 9040
rect 7640 20830 19880 20960
rect 7640 20590 7780 20830
rect 8020 20590 8110 20830
rect 8350 20590 8440 20830
rect 8680 20590 8770 20830
rect 9010 20590 9100 20830
rect 9340 20590 9430 20830
rect 9670 20590 9760 20830
rect 10000 20590 10090 20830
rect 10330 20590 10420 20830
rect 10660 20590 10750 20830
rect 10990 20590 11080 20830
rect 11320 20590 11410 20830
rect 11650 20590 11740 20830
rect 11980 20590 12070 20830
rect 12310 20590 12400 20830
rect 12640 20590 12730 20830
rect 12970 20590 13060 20830
rect 13300 20590 13390 20830
rect 13630 20590 13720 20830
rect 13960 20590 14050 20830
rect 14290 20590 14380 20830
rect 14620 20590 14710 20830
rect 14950 20590 15040 20830
rect 15280 20590 15370 20830
rect 15610 20590 15700 20830
rect 15940 20590 16030 20830
rect 16270 20590 16360 20830
rect 16600 20590 16690 20830
rect 16930 20590 17020 20830
rect 17260 20590 17350 20830
rect 17590 20590 17680 20830
rect 17920 20590 18010 20830
rect 18250 20590 18340 20830
rect 18580 20590 18670 20830
rect 18910 20590 19000 20830
rect 19240 20590 19330 20830
rect 19570 20590 19880 20830
rect 7640 20500 19880 20590
rect 7640 20260 7780 20500
rect 8020 20260 8110 20500
rect 8350 20260 8440 20500
rect 8680 20260 8770 20500
rect 9010 20260 9100 20500
rect 9340 20260 9430 20500
rect 9670 20260 9760 20500
rect 10000 20260 10090 20500
rect 10330 20260 10420 20500
rect 10660 20260 10750 20500
rect 10990 20260 11080 20500
rect 11320 20260 11410 20500
rect 11650 20260 11740 20500
rect 11980 20260 12070 20500
rect 12310 20260 12400 20500
rect 12640 20260 12730 20500
rect 12970 20260 13060 20500
rect 13300 20260 13390 20500
rect 13630 20260 13720 20500
rect 13960 20260 14050 20500
rect 14290 20260 14380 20500
rect 14620 20260 14710 20500
rect 14950 20260 15040 20500
rect 15280 20260 15370 20500
rect 15610 20260 15700 20500
rect 15940 20260 16030 20500
rect 16270 20260 16360 20500
rect 16600 20260 16690 20500
rect 16930 20260 17020 20500
rect 17260 20260 17350 20500
rect 17590 20260 17680 20500
rect 17920 20260 18010 20500
rect 18250 20260 18340 20500
rect 18580 20260 18670 20500
rect 18910 20260 19000 20500
rect 19240 20260 19330 20500
rect 19570 20260 19880 20500
rect 7640 20170 19880 20260
rect 7640 19930 7780 20170
rect 8020 19930 8110 20170
rect 8350 19930 8440 20170
rect 8680 19930 8770 20170
rect 9010 19930 9100 20170
rect 9340 19930 9430 20170
rect 9670 19930 9760 20170
rect 10000 19930 10090 20170
rect 10330 19930 10420 20170
rect 10660 19930 10750 20170
rect 10990 19930 11080 20170
rect 11320 19930 11410 20170
rect 11650 19930 11740 20170
rect 11980 19930 12070 20170
rect 12310 19930 12400 20170
rect 12640 19930 12730 20170
rect 12970 19930 13060 20170
rect 13300 19930 13390 20170
rect 13630 19930 13720 20170
rect 13960 19930 14050 20170
rect 14290 19930 14380 20170
rect 14620 19930 14710 20170
rect 14950 19930 15040 20170
rect 15280 19930 15370 20170
rect 15610 19930 15700 20170
rect 15940 19930 16030 20170
rect 16270 19930 16360 20170
rect 16600 19930 16690 20170
rect 16930 19930 17020 20170
rect 17260 19930 17350 20170
rect 17590 19930 17680 20170
rect 17920 19930 18010 20170
rect 18250 19930 18340 20170
rect 18580 19930 18670 20170
rect 18910 19930 19000 20170
rect 19240 19930 19330 20170
rect 19570 19930 19880 20170
rect 7640 19840 19880 19930
rect 7640 19600 7780 19840
rect 8020 19600 8110 19840
rect 8350 19600 8440 19840
rect 8680 19600 8770 19840
rect 9010 19600 9100 19840
rect 9340 19600 9430 19840
rect 9670 19600 9760 19840
rect 10000 19600 10090 19840
rect 10330 19600 10420 19840
rect 10660 19600 10750 19840
rect 10990 19600 11080 19840
rect 11320 19600 11410 19840
rect 11650 19600 11740 19840
rect 11980 19600 12070 19840
rect 12310 19600 12400 19840
rect 12640 19600 12730 19840
rect 12970 19600 13060 19840
rect 13300 19600 13390 19840
rect 13630 19600 13720 19840
rect 13960 19600 14050 19840
rect 14290 19600 14380 19840
rect 14620 19600 14710 19840
rect 14950 19600 15040 19840
rect 15280 19600 15370 19840
rect 15610 19600 15700 19840
rect 15940 19600 16030 19840
rect 16270 19600 16360 19840
rect 16600 19600 16690 19840
rect 16930 19600 17020 19840
rect 17260 19600 17350 19840
rect 17590 19600 17680 19840
rect 17920 19600 18010 19840
rect 18250 19600 18340 19840
rect 18580 19600 18670 19840
rect 18910 19600 19000 19840
rect 19240 19600 19330 19840
rect 19570 19600 19880 19840
rect 7640 19510 19880 19600
rect 7640 19270 7780 19510
rect 8020 19270 8110 19510
rect 8350 19270 8440 19510
rect 8680 19270 8770 19510
rect 9010 19270 9100 19510
rect 9340 19270 9430 19510
rect 9670 19270 9760 19510
rect 10000 19270 10090 19510
rect 10330 19270 10420 19510
rect 10660 19270 10750 19510
rect 10990 19270 11080 19510
rect 11320 19270 11410 19510
rect 11650 19270 11740 19510
rect 11980 19270 12070 19510
rect 12310 19270 12400 19510
rect 12640 19270 12730 19510
rect 12970 19270 13060 19510
rect 13300 19270 13390 19510
rect 13630 19270 13720 19510
rect 13960 19270 14050 19510
rect 14290 19270 14380 19510
rect 14620 19270 14710 19510
rect 14950 19270 15040 19510
rect 15280 19270 15370 19510
rect 15610 19270 15700 19510
rect 15940 19270 16030 19510
rect 16270 19270 16360 19510
rect 16600 19270 16690 19510
rect 16930 19270 17020 19510
rect 17260 19270 17350 19510
rect 17590 19270 17680 19510
rect 17920 19270 18010 19510
rect 18250 19270 18340 19510
rect 18580 19270 18670 19510
rect 18910 19270 19000 19510
rect 19240 19270 19330 19510
rect 19570 19270 19880 19510
rect 7640 19180 19880 19270
rect 7640 18940 7780 19180
rect 8020 18940 8110 19180
rect 8350 18940 8440 19180
rect 8680 18940 8770 19180
rect 9010 18940 9100 19180
rect 9340 18940 9430 19180
rect 9670 18940 9760 19180
rect 10000 18940 10090 19180
rect 10330 18940 10420 19180
rect 10660 18940 10750 19180
rect 10990 18940 11080 19180
rect 11320 18940 11410 19180
rect 11650 18940 11740 19180
rect 11980 18940 12070 19180
rect 12310 18940 12400 19180
rect 12640 18940 12730 19180
rect 12970 18940 13060 19180
rect 13300 18940 13390 19180
rect 13630 18940 13720 19180
rect 13960 18940 14050 19180
rect 14290 18940 14380 19180
rect 14620 18940 14710 19180
rect 14950 18940 15040 19180
rect 15280 18940 15370 19180
rect 15610 18940 15700 19180
rect 15940 18940 16030 19180
rect 16270 18940 16360 19180
rect 16600 18940 16690 19180
rect 16930 18940 17020 19180
rect 17260 18940 17350 19180
rect 17590 18940 17680 19180
rect 17920 18940 18010 19180
rect 18250 18940 18340 19180
rect 18580 18940 18670 19180
rect 18910 18940 19000 19180
rect 19240 18940 19330 19180
rect 19570 18940 19880 19180
rect 7640 18850 19880 18940
rect 7640 18610 7780 18850
rect 8020 18610 8110 18850
rect 8350 18610 8440 18850
rect 8680 18610 8770 18850
rect 9010 18610 9100 18850
rect 9340 18610 9430 18850
rect 9670 18610 9760 18850
rect 10000 18610 10090 18850
rect 10330 18610 10420 18850
rect 10660 18610 10750 18850
rect 10990 18610 11080 18850
rect 11320 18610 11410 18850
rect 11650 18610 11740 18850
rect 11980 18610 12070 18850
rect 12310 18610 12400 18850
rect 12640 18610 12730 18850
rect 12970 18610 13060 18850
rect 13300 18610 13390 18850
rect 13630 18610 13720 18850
rect 13960 18610 14050 18850
rect 14290 18610 14380 18850
rect 14620 18610 14710 18850
rect 14950 18610 15040 18850
rect 15280 18610 15370 18850
rect 15610 18610 15700 18850
rect 15940 18610 16030 18850
rect 16270 18610 16360 18850
rect 16600 18610 16690 18850
rect 16930 18610 17020 18850
rect 17260 18610 17350 18850
rect 17590 18610 17680 18850
rect 17920 18610 18010 18850
rect 18250 18610 18340 18850
rect 18580 18610 18670 18850
rect 18910 18610 19000 18850
rect 19240 18610 19330 18850
rect 19570 18610 19880 18850
rect 7640 18520 19880 18610
rect 7640 18280 7780 18520
rect 8020 18280 8110 18520
rect 8350 18280 8440 18520
rect 8680 18280 8770 18520
rect 9010 18280 9100 18520
rect 9340 18280 9430 18520
rect 9670 18280 9760 18520
rect 10000 18280 10090 18520
rect 10330 18280 10420 18520
rect 10660 18280 10750 18520
rect 10990 18280 11080 18520
rect 11320 18280 11410 18520
rect 11650 18280 11740 18520
rect 11980 18280 12070 18520
rect 12310 18280 12400 18520
rect 12640 18280 12730 18520
rect 12970 18280 13060 18520
rect 13300 18280 13390 18520
rect 13630 18280 13720 18520
rect 13960 18280 14050 18520
rect 14290 18280 14380 18520
rect 14620 18280 14710 18520
rect 14950 18280 15040 18520
rect 15280 18280 15370 18520
rect 15610 18280 15700 18520
rect 15940 18280 16030 18520
rect 16270 18280 16360 18520
rect 16600 18280 16690 18520
rect 16930 18280 17020 18520
rect 17260 18280 17350 18520
rect 17590 18280 17680 18520
rect 17920 18280 18010 18520
rect 18250 18280 18340 18520
rect 18580 18280 18670 18520
rect 18910 18280 19000 18520
rect 19240 18280 19330 18520
rect 19570 18280 19880 18520
rect 7640 18190 19880 18280
rect 7640 17950 7780 18190
rect 8020 17950 8110 18190
rect 8350 17950 8440 18190
rect 8680 17950 8770 18190
rect 9010 17950 9100 18190
rect 9340 17950 9430 18190
rect 9670 17950 9760 18190
rect 10000 17950 10090 18190
rect 10330 17950 10420 18190
rect 10660 17950 10750 18190
rect 10990 17950 11080 18190
rect 11320 17950 11410 18190
rect 11650 17950 11740 18190
rect 11980 17950 12070 18190
rect 12310 17950 12400 18190
rect 12640 17950 12730 18190
rect 12970 17950 13060 18190
rect 13300 17950 13390 18190
rect 13630 17950 13720 18190
rect 13960 17950 14050 18190
rect 14290 17950 14380 18190
rect 14620 17950 14710 18190
rect 14950 17950 15040 18190
rect 15280 17950 15370 18190
rect 15610 17950 15700 18190
rect 15940 17950 16030 18190
rect 16270 17950 16360 18190
rect 16600 17950 16690 18190
rect 16930 17950 17020 18190
rect 17260 17950 17350 18190
rect 17590 17950 17680 18190
rect 17920 17950 18010 18190
rect 18250 17950 18340 18190
rect 18580 17950 18670 18190
rect 18910 17950 19000 18190
rect 19240 17950 19330 18190
rect 19570 17950 19880 18190
rect 7640 17860 19880 17950
rect 7640 17620 7780 17860
rect 8020 17620 8110 17860
rect 8350 17620 8440 17860
rect 8680 17620 8770 17860
rect 9010 17620 9100 17860
rect 9340 17620 9430 17860
rect 9670 17620 9760 17860
rect 10000 17620 10090 17860
rect 10330 17620 10420 17860
rect 10660 17620 10750 17860
rect 10990 17620 11080 17860
rect 11320 17620 11410 17860
rect 11650 17620 11740 17860
rect 11980 17620 12070 17860
rect 12310 17620 12400 17860
rect 12640 17620 12730 17860
rect 12970 17620 13060 17860
rect 13300 17620 13390 17860
rect 13630 17620 13720 17860
rect 13960 17620 14050 17860
rect 14290 17620 14380 17860
rect 14620 17620 14710 17860
rect 14950 17620 15040 17860
rect 15280 17620 15370 17860
rect 15610 17620 15700 17860
rect 15940 17620 16030 17860
rect 16270 17620 16360 17860
rect 16600 17620 16690 17860
rect 16930 17620 17020 17860
rect 17260 17620 17350 17860
rect 17590 17620 17680 17860
rect 17920 17620 18010 17860
rect 18250 17620 18340 17860
rect 18580 17620 18670 17860
rect 18910 17620 19000 17860
rect 19240 17620 19330 17860
rect 19570 17620 19880 17860
rect 7640 17530 19880 17620
rect 7640 17290 7780 17530
rect 8020 17290 8110 17530
rect 8350 17290 8440 17530
rect 8680 17290 8770 17530
rect 9010 17290 9100 17530
rect 9340 17290 9430 17530
rect 9670 17290 9760 17530
rect 10000 17290 10090 17530
rect 10330 17290 10420 17530
rect 10660 17290 10750 17530
rect 10990 17290 11080 17530
rect 11320 17290 11410 17530
rect 11650 17290 11740 17530
rect 11980 17290 12070 17530
rect 12310 17290 12400 17530
rect 12640 17290 12730 17530
rect 12970 17290 13060 17530
rect 13300 17290 13390 17530
rect 13630 17290 13720 17530
rect 13960 17290 14050 17530
rect 14290 17290 14380 17530
rect 14620 17290 14710 17530
rect 14950 17290 15040 17530
rect 15280 17290 15370 17530
rect 15610 17290 15700 17530
rect 15940 17290 16030 17530
rect 16270 17290 16360 17530
rect 16600 17290 16690 17530
rect 16930 17290 17020 17530
rect 17260 17290 17350 17530
rect 17590 17290 17680 17530
rect 17920 17290 18010 17530
rect 18250 17290 18340 17530
rect 18580 17290 18670 17530
rect 18910 17290 19000 17530
rect 19240 17290 19330 17530
rect 19570 17290 19880 17530
rect 7640 17200 19880 17290
rect 7640 16960 7780 17200
rect 8020 16960 8110 17200
rect 8350 16960 8440 17200
rect 8680 16960 8770 17200
rect 9010 16960 9100 17200
rect 9340 16960 9430 17200
rect 9670 16960 9760 17200
rect 10000 16960 10090 17200
rect 10330 16960 10420 17200
rect 10660 16960 10750 17200
rect 10990 16960 11080 17200
rect 11320 16960 11410 17200
rect 11650 16960 11740 17200
rect 11980 16960 12070 17200
rect 12310 16960 12400 17200
rect 12640 16960 12730 17200
rect 12970 16960 13060 17200
rect 13300 16960 13390 17200
rect 13630 16960 13720 17200
rect 13960 16960 14050 17200
rect 14290 16960 14380 17200
rect 14620 16960 14710 17200
rect 14950 16960 15040 17200
rect 15280 16960 15370 17200
rect 15610 16960 15700 17200
rect 15940 16960 16030 17200
rect 16270 16960 16360 17200
rect 16600 16960 16690 17200
rect 16930 16960 17020 17200
rect 17260 16960 17350 17200
rect 17590 16960 17680 17200
rect 17920 16960 18010 17200
rect 18250 16960 18340 17200
rect 18580 16960 18670 17200
rect 18910 16960 19000 17200
rect 19240 16960 19330 17200
rect 19570 16960 19880 17200
rect 7640 16870 19880 16960
rect 7640 16630 7780 16870
rect 8020 16630 8110 16870
rect 8350 16630 8440 16870
rect 8680 16630 8770 16870
rect 9010 16630 9100 16870
rect 9340 16630 9430 16870
rect 9670 16630 9760 16870
rect 10000 16630 10090 16870
rect 10330 16630 10420 16870
rect 10660 16630 10750 16870
rect 10990 16630 11080 16870
rect 11320 16630 11410 16870
rect 11650 16630 11740 16870
rect 11980 16630 12070 16870
rect 12310 16630 12400 16870
rect 12640 16630 12730 16870
rect 12970 16630 13060 16870
rect 13300 16630 13390 16870
rect 13630 16630 13720 16870
rect 13960 16630 14050 16870
rect 14290 16630 14380 16870
rect 14620 16630 14710 16870
rect 14950 16630 15040 16870
rect 15280 16630 15370 16870
rect 15610 16630 15700 16870
rect 15940 16630 16030 16870
rect 16270 16630 16360 16870
rect 16600 16630 16690 16870
rect 16930 16630 17020 16870
rect 17260 16630 17350 16870
rect 17590 16630 17680 16870
rect 17920 16630 18010 16870
rect 18250 16630 18340 16870
rect 18580 16630 18670 16870
rect 18910 16630 19000 16870
rect 19240 16630 19330 16870
rect 19570 16630 19880 16870
rect 7640 16540 19880 16630
rect 7640 16300 7780 16540
rect 8020 16300 8110 16540
rect 8350 16300 8440 16540
rect 8680 16300 8770 16540
rect 9010 16300 9100 16540
rect 9340 16300 9430 16540
rect 9670 16300 9760 16540
rect 10000 16300 10090 16540
rect 10330 16300 10420 16540
rect 10660 16300 10750 16540
rect 10990 16300 11080 16540
rect 11320 16300 11410 16540
rect 11650 16300 11740 16540
rect 11980 16300 12070 16540
rect 12310 16300 12400 16540
rect 12640 16300 12730 16540
rect 12970 16300 13060 16540
rect 13300 16300 13390 16540
rect 13630 16300 13720 16540
rect 13960 16300 14050 16540
rect 14290 16300 14380 16540
rect 14620 16300 14710 16540
rect 14950 16300 15040 16540
rect 15280 16300 15370 16540
rect 15610 16300 15700 16540
rect 15940 16300 16030 16540
rect 16270 16300 16360 16540
rect 16600 16300 16690 16540
rect 16930 16300 17020 16540
rect 17260 16300 17350 16540
rect 17590 16300 17680 16540
rect 17920 16300 18010 16540
rect 18250 16300 18340 16540
rect 18580 16300 18670 16540
rect 18910 16300 19000 16540
rect 19240 16300 19330 16540
rect 19570 16300 19880 16540
rect 7640 16210 19880 16300
rect 7640 15970 7780 16210
rect 8020 15970 8110 16210
rect 8350 15970 8440 16210
rect 8680 15970 8770 16210
rect 9010 15970 9100 16210
rect 9340 15970 9430 16210
rect 9670 15970 9760 16210
rect 10000 15970 10090 16210
rect 10330 15970 10420 16210
rect 10660 15970 10750 16210
rect 10990 15970 11080 16210
rect 11320 15970 11410 16210
rect 11650 15970 11740 16210
rect 11980 15970 12070 16210
rect 12310 15970 12400 16210
rect 12640 15970 12730 16210
rect 12970 15970 13060 16210
rect 13300 15970 13390 16210
rect 13630 15970 13720 16210
rect 13960 15970 14050 16210
rect 14290 15970 14380 16210
rect 14620 15970 14710 16210
rect 14950 15970 15040 16210
rect 15280 15970 15370 16210
rect 15610 15970 15700 16210
rect 15940 15970 16030 16210
rect 16270 15970 16360 16210
rect 16600 15970 16690 16210
rect 16930 15970 17020 16210
rect 17260 15970 17350 16210
rect 17590 15970 17680 16210
rect 17920 15970 18010 16210
rect 18250 15970 18340 16210
rect 18580 15970 18670 16210
rect 18910 15970 19000 16210
rect 19240 15970 19330 16210
rect 19570 15970 19880 16210
rect 7640 15880 19880 15970
rect 7640 15640 7780 15880
rect 8020 15640 8110 15880
rect 8350 15640 8440 15880
rect 8680 15640 8770 15880
rect 9010 15640 9100 15880
rect 9340 15640 9430 15880
rect 9670 15640 9760 15880
rect 10000 15640 10090 15880
rect 10330 15640 10420 15880
rect 10660 15640 10750 15880
rect 10990 15640 11080 15880
rect 11320 15640 11410 15880
rect 11650 15640 11740 15880
rect 11980 15640 12070 15880
rect 12310 15640 12400 15880
rect 12640 15640 12730 15880
rect 12970 15640 13060 15880
rect 13300 15640 13390 15880
rect 13630 15640 13720 15880
rect 13960 15640 14050 15880
rect 14290 15640 14380 15880
rect 14620 15640 14710 15880
rect 14950 15640 15040 15880
rect 15280 15640 15370 15880
rect 15610 15640 15700 15880
rect 15940 15640 16030 15880
rect 16270 15640 16360 15880
rect 16600 15640 16690 15880
rect 16930 15640 17020 15880
rect 17260 15640 17350 15880
rect 17590 15640 17680 15880
rect 17920 15640 18010 15880
rect 18250 15640 18340 15880
rect 18580 15640 18670 15880
rect 18910 15640 19000 15880
rect 19240 15640 19330 15880
rect 19570 15640 19880 15880
rect 7640 15550 19880 15640
rect 7640 15310 7780 15550
rect 8020 15310 8110 15550
rect 8350 15310 8440 15550
rect 8680 15310 8770 15550
rect 9010 15310 9100 15550
rect 9340 15310 9430 15550
rect 9670 15310 9760 15550
rect 10000 15310 10090 15550
rect 10330 15310 10420 15550
rect 10660 15310 10750 15550
rect 10990 15310 11080 15550
rect 11320 15310 11410 15550
rect 11650 15310 11740 15550
rect 11980 15310 12070 15550
rect 12310 15310 12400 15550
rect 12640 15310 12730 15550
rect 12970 15310 13060 15550
rect 13300 15310 13390 15550
rect 13630 15310 13720 15550
rect 13960 15310 14050 15550
rect 14290 15310 14380 15550
rect 14620 15310 14710 15550
rect 14950 15310 15040 15550
rect 15280 15310 15370 15550
rect 15610 15310 15700 15550
rect 15940 15310 16030 15550
rect 16270 15310 16360 15550
rect 16600 15310 16690 15550
rect 16930 15310 17020 15550
rect 17260 15310 17350 15550
rect 17590 15310 17680 15550
rect 17920 15310 18010 15550
rect 18250 15310 18340 15550
rect 18580 15310 18670 15550
rect 18910 15310 19000 15550
rect 19240 15310 19330 15550
rect 19570 15310 19880 15550
rect 7640 15220 19880 15310
rect 7640 14980 7780 15220
rect 8020 14980 8110 15220
rect 8350 14980 8440 15220
rect 8680 14980 8770 15220
rect 9010 14980 9100 15220
rect 9340 14980 9430 15220
rect 9670 14980 9760 15220
rect 10000 14980 10090 15220
rect 10330 14980 10420 15220
rect 10660 14980 10750 15220
rect 10990 14980 11080 15220
rect 11320 14980 11410 15220
rect 11650 14980 11740 15220
rect 11980 14980 12070 15220
rect 12310 14980 12400 15220
rect 12640 14980 12730 15220
rect 12970 14980 13060 15220
rect 13300 14980 13390 15220
rect 13630 14980 13720 15220
rect 13960 14980 14050 15220
rect 14290 14980 14380 15220
rect 14620 14980 14710 15220
rect 14950 14980 15040 15220
rect 15280 14980 15370 15220
rect 15610 14980 15700 15220
rect 15940 14980 16030 15220
rect 16270 14980 16360 15220
rect 16600 14980 16690 15220
rect 16930 14980 17020 15220
rect 17260 14980 17350 15220
rect 17590 14980 17680 15220
rect 17920 14980 18010 15220
rect 18250 14980 18340 15220
rect 18580 14980 18670 15220
rect 18910 14980 19000 15220
rect 19240 14980 19330 15220
rect 19570 14980 19880 15220
rect 7640 14890 19880 14980
rect 7640 14650 7780 14890
rect 8020 14650 8110 14890
rect 8350 14650 8440 14890
rect 8680 14650 8770 14890
rect 9010 14650 9100 14890
rect 9340 14650 9430 14890
rect 9670 14650 9760 14890
rect 10000 14650 10090 14890
rect 10330 14650 10420 14890
rect 10660 14650 10750 14890
rect 10990 14650 11080 14890
rect 11320 14650 11410 14890
rect 11650 14650 11740 14890
rect 11980 14650 12070 14890
rect 12310 14650 12400 14890
rect 12640 14650 12730 14890
rect 12970 14650 13060 14890
rect 13300 14650 13390 14890
rect 13630 14650 13720 14890
rect 13960 14650 14050 14890
rect 14290 14650 14380 14890
rect 14620 14650 14710 14890
rect 14950 14650 15040 14890
rect 15280 14650 15370 14890
rect 15610 14650 15700 14890
rect 15940 14650 16030 14890
rect 16270 14650 16360 14890
rect 16600 14650 16690 14890
rect 16930 14650 17020 14890
rect 17260 14650 17350 14890
rect 17590 14650 17680 14890
rect 17920 14650 18010 14890
rect 18250 14650 18340 14890
rect 18580 14650 18670 14890
rect 18910 14650 19000 14890
rect 19240 14650 19330 14890
rect 19570 14650 19880 14890
rect 7640 14560 19880 14650
rect 7640 14320 7780 14560
rect 8020 14320 8110 14560
rect 8350 14320 8440 14560
rect 8680 14320 8770 14560
rect 9010 14320 9100 14560
rect 9340 14320 9430 14560
rect 9670 14320 9760 14560
rect 10000 14320 10090 14560
rect 10330 14320 10420 14560
rect 10660 14320 10750 14560
rect 10990 14320 11080 14560
rect 11320 14320 11410 14560
rect 11650 14320 11740 14560
rect 11980 14320 12070 14560
rect 12310 14320 12400 14560
rect 12640 14320 12730 14560
rect 12970 14320 13060 14560
rect 13300 14320 13390 14560
rect 13630 14320 13720 14560
rect 13960 14320 14050 14560
rect 14290 14320 14380 14560
rect 14620 14320 14710 14560
rect 14950 14320 15040 14560
rect 15280 14320 15370 14560
rect 15610 14320 15700 14560
rect 15940 14320 16030 14560
rect 16270 14320 16360 14560
rect 16600 14320 16690 14560
rect 16930 14320 17020 14560
rect 17260 14320 17350 14560
rect 17590 14320 17680 14560
rect 17920 14320 18010 14560
rect 18250 14320 18340 14560
rect 18580 14320 18670 14560
rect 18910 14320 19000 14560
rect 19240 14320 19330 14560
rect 19570 14320 19880 14560
rect 7640 14230 19880 14320
rect 7640 13990 7780 14230
rect 8020 13990 8110 14230
rect 8350 13990 8440 14230
rect 8680 13990 8770 14230
rect 9010 13990 9100 14230
rect 9340 13990 9430 14230
rect 9670 13990 9760 14230
rect 10000 13990 10090 14230
rect 10330 13990 10420 14230
rect 10660 13990 10750 14230
rect 10990 13990 11080 14230
rect 11320 13990 11410 14230
rect 11650 13990 11740 14230
rect 11980 13990 12070 14230
rect 12310 13990 12400 14230
rect 12640 13990 12730 14230
rect 12970 13990 13060 14230
rect 13300 13990 13390 14230
rect 13630 13990 13720 14230
rect 13960 13990 14050 14230
rect 14290 13990 14380 14230
rect 14620 13990 14710 14230
rect 14950 13990 15040 14230
rect 15280 13990 15370 14230
rect 15610 13990 15700 14230
rect 15940 13990 16030 14230
rect 16270 13990 16360 14230
rect 16600 13990 16690 14230
rect 16930 13990 17020 14230
rect 17260 13990 17350 14230
rect 17590 13990 17680 14230
rect 17920 13990 18010 14230
rect 18250 13990 18340 14230
rect 18580 13990 18670 14230
rect 18910 13990 19000 14230
rect 19240 13990 19330 14230
rect 19570 13990 19880 14230
rect 7640 13900 19880 13990
rect 7640 13660 7780 13900
rect 8020 13660 8110 13900
rect 8350 13660 8440 13900
rect 8680 13660 8770 13900
rect 9010 13660 9100 13900
rect 9340 13660 9430 13900
rect 9670 13660 9760 13900
rect 10000 13660 10090 13900
rect 10330 13660 10420 13900
rect 10660 13660 10750 13900
rect 10990 13660 11080 13900
rect 11320 13660 11410 13900
rect 11650 13660 11740 13900
rect 11980 13660 12070 13900
rect 12310 13660 12400 13900
rect 12640 13660 12730 13900
rect 12970 13660 13060 13900
rect 13300 13660 13390 13900
rect 13630 13660 13720 13900
rect 13960 13660 14050 13900
rect 14290 13660 14380 13900
rect 14620 13660 14710 13900
rect 14950 13660 15040 13900
rect 15280 13660 15370 13900
rect 15610 13660 15700 13900
rect 15940 13660 16030 13900
rect 16270 13660 16360 13900
rect 16600 13660 16690 13900
rect 16930 13660 17020 13900
rect 17260 13660 17350 13900
rect 17590 13660 17680 13900
rect 17920 13660 18010 13900
rect 18250 13660 18340 13900
rect 18580 13660 18670 13900
rect 18910 13660 19000 13900
rect 19240 13660 19330 13900
rect 19570 13660 19880 13900
rect 7640 13570 19880 13660
rect 7640 13330 7780 13570
rect 8020 13330 8110 13570
rect 8350 13330 8440 13570
rect 8680 13330 8770 13570
rect 9010 13330 9100 13570
rect 9340 13330 9430 13570
rect 9670 13330 9760 13570
rect 10000 13330 10090 13570
rect 10330 13330 10420 13570
rect 10660 13330 10750 13570
rect 10990 13330 11080 13570
rect 11320 13330 11410 13570
rect 11650 13330 11740 13570
rect 11980 13330 12070 13570
rect 12310 13330 12400 13570
rect 12640 13330 12730 13570
rect 12970 13330 13060 13570
rect 13300 13330 13390 13570
rect 13630 13330 13720 13570
rect 13960 13330 14050 13570
rect 14290 13330 14380 13570
rect 14620 13330 14710 13570
rect 14950 13330 15040 13570
rect 15280 13330 15370 13570
rect 15610 13330 15700 13570
rect 15940 13330 16030 13570
rect 16270 13330 16360 13570
rect 16600 13330 16690 13570
rect 16930 13330 17020 13570
rect 17260 13330 17350 13570
rect 17590 13330 17680 13570
rect 17920 13330 18010 13570
rect 18250 13330 18340 13570
rect 18580 13330 18670 13570
rect 18910 13330 19000 13570
rect 19240 13330 19330 13570
rect 19570 13330 19880 13570
rect 7640 13240 19880 13330
rect 7640 13000 7780 13240
rect 8020 13000 8110 13240
rect 8350 13000 8440 13240
rect 8680 13000 8770 13240
rect 9010 13000 9100 13240
rect 9340 13000 9430 13240
rect 9670 13000 9760 13240
rect 10000 13000 10090 13240
rect 10330 13000 10420 13240
rect 10660 13000 10750 13240
rect 10990 13000 11080 13240
rect 11320 13000 11410 13240
rect 11650 13000 11740 13240
rect 11980 13000 12070 13240
rect 12310 13000 12400 13240
rect 12640 13000 12730 13240
rect 12970 13000 13060 13240
rect 13300 13000 13390 13240
rect 13630 13000 13720 13240
rect 13960 13000 14050 13240
rect 14290 13000 14380 13240
rect 14620 13000 14710 13240
rect 14950 13000 15040 13240
rect 15280 13000 15370 13240
rect 15610 13000 15700 13240
rect 15940 13000 16030 13240
rect 16270 13000 16360 13240
rect 16600 13000 16690 13240
rect 16930 13000 17020 13240
rect 17260 13000 17350 13240
rect 17590 13000 17680 13240
rect 17920 13000 18010 13240
rect 18250 13000 18340 13240
rect 18580 13000 18670 13240
rect 18910 13000 19000 13240
rect 19240 13000 19330 13240
rect 19570 13000 19880 13240
rect 7640 12910 19880 13000
rect 7640 12670 7780 12910
rect 8020 12670 8110 12910
rect 8350 12670 8440 12910
rect 8680 12670 8770 12910
rect 9010 12670 9100 12910
rect 9340 12670 9430 12910
rect 9670 12670 9760 12910
rect 10000 12670 10090 12910
rect 10330 12670 10420 12910
rect 10660 12670 10750 12910
rect 10990 12670 11080 12910
rect 11320 12670 11410 12910
rect 11650 12670 11740 12910
rect 11980 12670 12070 12910
rect 12310 12670 12400 12910
rect 12640 12670 12730 12910
rect 12970 12670 13060 12910
rect 13300 12670 13390 12910
rect 13630 12670 13720 12910
rect 13960 12670 14050 12910
rect 14290 12670 14380 12910
rect 14620 12670 14710 12910
rect 14950 12670 15040 12910
rect 15280 12670 15370 12910
rect 15610 12670 15700 12910
rect 15940 12670 16030 12910
rect 16270 12670 16360 12910
rect 16600 12670 16690 12910
rect 16930 12670 17020 12910
rect 17260 12670 17350 12910
rect 17590 12670 17680 12910
rect 17920 12670 18010 12910
rect 18250 12670 18340 12910
rect 18580 12670 18670 12910
rect 18910 12670 19000 12910
rect 19240 12670 19330 12910
rect 19570 12670 19880 12910
rect 7640 12580 19880 12670
rect 7640 12340 7780 12580
rect 8020 12340 8110 12580
rect 8350 12340 8440 12580
rect 8680 12340 8770 12580
rect 9010 12340 9100 12580
rect 9340 12340 9430 12580
rect 9670 12340 9760 12580
rect 10000 12340 10090 12580
rect 10330 12340 10420 12580
rect 10660 12340 10750 12580
rect 10990 12340 11080 12580
rect 11320 12340 11410 12580
rect 11650 12340 11740 12580
rect 11980 12340 12070 12580
rect 12310 12340 12400 12580
rect 12640 12340 12730 12580
rect 12970 12340 13060 12580
rect 13300 12340 13390 12580
rect 13630 12340 13720 12580
rect 13960 12340 14050 12580
rect 14290 12340 14380 12580
rect 14620 12340 14710 12580
rect 14950 12340 15040 12580
rect 15280 12340 15370 12580
rect 15610 12340 15700 12580
rect 15940 12340 16030 12580
rect 16270 12340 16360 12580
rect 16600 12340 16690 12580
rect 16930 12340 17020 12580
rect 17260 12340 17350 12580
rect 17590 12340 17680 12580
rect 17920 12340 18010 12580
rect 18250 12340 18340 12580
rect 18580 12340 18670 12580
rect 18910 12340 19000 12580
rect 19240 12340 19330 12580
rect 19570 12340 19880 12580
rect 7640 12250 19880 12340
rect 7640 12010 7780 12250
rect 8020 12010 8110 12250
rect 8350 12010 8440 12250
rect 8680 12010 8770 12250
rect 9010 12010 9100 12250
rect 9340 12010 9430 12250
rect 9670 12010 9760 12250
rect 10000 12010 10090 12250
rect 10330 12010 10420 12250
rect 10660 12010 10750 12250
rect 10990 12010 11080 12250
rect 11320 12010 11410 12250
rect 11650 12010 11740 12250
rect 11980 12010 12070 12250
rect 12310 12010 12400 12250
rect 12640 12010 12730 12250
rect 12970 12010 13060 12250
rect 13300 12010 13390 12250
rect 13630 12010 13720 12250
rect 13960 12010 14050 12250
rect 14290 12010 14380 12250
rect 14620 12010 14710 12250
rect 14950 12010 15040 12250
rect 15280 12010 15370 12250
rect 15610 12010 15700 12250
rect 15940 12010 16030 12250
rect 16270 12010 16360 12250
rect 16600 12010 16690 12250
rect 16930 12010 17020 12250
rect 17260 12010 17350 12250
rect 17590 12010 17680 12250
rect 17920 12010 18010 12250
rect 18250 12010 18340 12250
rect 18580 12010 18670 12250
rect 18910 12010 19000 12250
rect 19240 12010 19330 12250
rect 19570 12010 19880 12250
rect 7640 11920 19880 12010
rect 7640 11680 7780 11920
rect 8020 11680 8110 11920
rect 8350 11680 8440 11920
rect 8680 11680 8770 11920
rect 9010 11680 9100 11920
rect 9340 11680 9430 11920
rect 9670 11680 9760 11920
rect 10000 11680 10090 11920
rect 10330 11680 10420 11920
rect 10660 11680 10750 11920
rect 10990 11680 11080 11920
rect 11320 11680 11410 11920
rect 11650 11680 11740 11920
rect 11980 11680 12070 11920
rect 12310 11680 12400 11920
rect 12640 11680 12730 11920
rect 12970 11680 13060 11920
rect 13300 11680 13390 11920
rect 13630 11680 13720 11920
rect 13960 11680 14050 11920
rect 14290 11680 14380 11920
rect 14620 11680 14710 11920
rect 14950 11680 15040 11920
rect 15280 11680 15370 11920
rect 15610 11680 15700 11920
rect 15940 11680 16030 11920
rect 16270 11680 16360 11920
rect 16600 11680 16690 11920
rect 16930 11680 17020 11920
rect 17260 11680 17350 11920
rect 17590 11680 17680 11920
rect 17920 11680 18010 11920
rect 18250 11680 18340 11920
rect 18580 11680 18670 11920
rect 18910 11680 19000 11920
rect 19240 11680 19330 11920
rect 19570 11680 19880 11920
rect 7640 11590 19880 11680
rect 7640 11350 7780 11590
rect 8020 11350 8110 11590
rect 8350 11350 8440 11590
rect 8680 11350 8770 11590
rect 9010 11350 9100 11590
rect 9340 11350 9430 11590
rect 9670 11350 9760 11590
rect 10000 11350 10090 11590
rect 10330 11350 10420 11590
rect 10660 11350 10750 11590
rect 10990 11350 11080 11590
rect 11320 11350 11410 11590
rect 11650 11350 11740 11590
rect 11980 11350 12070 11590
rect 12310 11350 12400 11590
rect 12640 11350 12730 11590
rect 12970 11350 13060 11590
rect 13300 11350 13390 11590
rect 13630 11350 13720 11590
rect 13960 11350 14050 11590
rect 14290 11350 14380 11590
rect 14620 11350 14710 11590
rect 14950 11350 15040 11590
rect 15280 11350 15370 11590
rect 15610 11350 15700 11590
rect 15940 11350 16030 11590
rect 16270 11350 16360 11590
rect 16600 11350 16690 11590
rect 16930 11350 17020 11590
rect 17260 11350 17350 11590
rect 17590 11350 17680 11590
rect 17920 11350 18010 11590
rect 18250 11350 18340 11590
rect 18580 11350 18670 11590
rect 18910 11350 19000 11590
rect 19240 11350 19330 11590
rect 19570 11350 19880 11590
rect 7640 11260 19880 11350
rect 7640 11020 7780 11260
rect 8020 11020 8110 11260
rect 8350 11020 8440 11260
rect 8680 11020 8770 11260
rect 9010 11020 9100 11260
rect 9340 11020 9430 11260
rect 9670 11020 9760 11260
rect 10000 11020 10090 11260
rect 10330 11020 10420 11260
rect 10660 11020 10750 11260
rect 10990 11020 11080 11260
rect 11320 11020 11410 11260
rect 11650 11020 11740 11260
rect 11980 11020 12070 11260
rect 12310 11020 12400 11260
rect 12640 11020 12730 11260
rect 12970 11020 13060 11260
rect 13300 11020 13390 11260
rect 13630 11020 13720 11260
rect 13960 11020 14050 11260
rect 14290 11020 14380 11260
rect 14620 11020 14710 11260
rect 14950 11020 15040 11260
rect 15280 11020 15370 11260
rect 15610 11020 15700 11260
rect 15940 11020 16030 11260
rect 16270 11020 16360 11260
rect 16600 11020 16690 11260
rect 16930 11020 17020 11260
rect 17260 11020 17350 11260
rect 17590 11020 17680 11260
rect 17920 11020 18010 11260
rect 18250 11020 18340 11260
rect 18580 11020 18670 11260
rect 18910 11020 19000 11260
rect 19240 11020 19330 11260
rect 19570 11020 19880 11260
rect 7640 10930 19880 11020
rect 7640 10690 7780 10930
rect 8020 10690 8110 10930
rect 8350 10690 8440 10930
rect 8680 10690 8770 10930
rect 9010 10690 9100 10930
rect 9340 10690 9430 10930
rect 9670 10690 9760 10930
rect 10000 10690 10090 10930
rect 10330 10690 10420 10930
rect 10660 10690 10750 10930
rect 10990 10690 11080 10930
rect 11320 10690 11410 10930
rect 11650 10690 11740 10930
rect 11980 10690 12070 10930
rect 12310 10690 12400 10930
rect 12640 10690 12730 10930
rect 12970 10690 13060 10930
rect 13300 10690 13390 10930
rect 13630 10690 13720 10930
rect 13960 10690 14050 10930
rect 14290 10690 14380 10930
rect 14620 10690 14710 10930
rect 14950 10690 15040 10930
rect 15280 10690 15370 10930
rect 15610 10690 15700 10930
rect 15940 10690 16030 10930
rect 16270 10690 16360 10930
rect 16600 10690 16690 10930
rect 16930 10690 17020 10930
rect 17260 10690 17350 10930
rect 17590 10690 17680 10930
rect 17920 10690 18010 10930
rect 18250 10690 18340 10930
rect 18580 10690 18670 10930
rect 18910 10690 19000 10930
rect 19240 10690 19330 10930
rect 19570 10690 19880 10930
rect 7640 10600 19880 10690
rect 7640 10360 7780 10600
rect 8020 10360 8110 10600
rect 8350 10360 8440 10600
rect 8680 10360 8770 10600
rect 9010 10360 9100 10600
rect 9340 10360 9430 10600
rect 9670 10360 9760 10600
rect 10000 10360 10090 10600
rect 10330 10360 10420 10600
rect 10660 10360 10750 10600
rect 10990 10360 11080 10600
rect 11320 10360 11410 10600
rect 11650 10360 11740 10600
rect 11980 10360 12070 10600
rect 12310 10360 12400 10600
rect 12640 10360 12730 10600
rect 12970 10360 13060 10600
rect 13300 10360 13390 10600
rect 13630 10360 13720 10600
rect 13960 10360 14050 10600
rect 14290 10360 14380 10600
rect 14620 10360 14710 10600
rect 14950 10360 15040 10600
rect 15280 10360 15370 10600
rect 15610 10360 15700 10600
rect 15940 10360 16030 10600
rect 16270 10360 16360 10600
rect 16600 10360 16690 10600
rect 16930 10360 17020 10600
rect 17260 10360 17350 10600
rect 17590 10360 17680 10600
rect 17920 10360 18010 10600
rect 18250 10360 18340 10600
rect 18580 10360 18670 10600
rect 18910 10360 19000 10600
rect 19240 10360 19330 10600
rect 19570 10360 19880 10600
rect 7640 10270 19880 10360
rect 7640 10030 7780 10270
rect 8020 10030 8110 10270
rect 8350 10030 8440 10270
rect 8680 10030 8770 10270
rect 9010 10030 9100 10270
rect 9340 10030 9430 10270
rect 9670 10030 9760 10270
rect 10000 10030 10090 10270
rect 10330 10030 10420 10270
rect 10660 10030 10750 10270
rect 10990 10030 11080 10270
rect 11320 10030 11410 10270
rect 11650 10030 11740 10270
rect 11980 10030 12070 10270
rect 12310 10030 12400 10270
rect 12640 10030 12730 10270
rect 12970 10030 13060 10270
rect 13300 10030 13390 10270
rect 13630 10030 13720 10270
rect 13960 10030 14050 10270
rect 14290 10030 14380 10270
rect 14620 10030 14710 10270
rect 14950 10030 15040 10270
rect 15280 10030 15370 10270
rect 15610 10030 15700 10270
rect 15940 10030 16030 10270
rect 16270 10030 16360 10270
rect 16600 10030 16690 10270
rect 16930 10030 17020 10270
rect 17260 10030 17350 10270
rect 17590 10030 17680 10270
rect 17920 10030 18010 10270
rect 18250 10030 18340 10270
rect 18580 10030 18670 10270
rect 18910 10030 19000 10270
rect 19240 10030 19330 10270
rect 19570 10030 19880 10270
rect 7640 9940 19880 10030
rect 7640 9700 7780 9940
rect 8020 9700 8110 9940
rect 8350 9700 8440 9940
rect 8680 9700 8770 9940
rect 9010 9700 9100 9940
rect 9340 9700 9430 9940
rect 9670 9700 9760 9940
rect 10000 9700 10090 9940
rect 10330 9700 10420 9940
rect 10660 9700 10750 9940
rect 10990 9700 11080 9940
rect 11320 9700 11410 9940
rect 11650 9700 11740 9940
rect 11980 9700 12070 9940
rect 12310 9700 12400 9940
rect 12640 9700 12730 9940
rect 12970 9700 13060 9940
rect 13300 9700 13390 9940
rect 13630 9700 13720 9940
rect 13960 9700 14050 9940
rect 14290 9700 14380 9940
rect 14620 9700 14710 9940
rect 14950 9700 15040 9940
rect 15280 9700 15370 9940
rect 15610 9700 15700 9940
rect 15940 9700 16030 9940
rect 16270 9700 16360 9940
rect 16600 9700 16690 9940
rect 16930 9700 17020 9940
rect 17260 9700 17350 9940
rect 17590 9700 17680 9940
rect 17920 9700 18010 9940
rect 18250 9700 18340 9940
rect 18580 9700 18670 9940
rect 18910 9700 19000 9940
rect 19240 9700 19330 9940
rect 19570 9700 19880 9940
rect 7640 9610 19880 9700
rect 7640 9370 7780 9610
rect 8020 9370 8110 9610
rect 8350 9370 8440 9610
rect 8680 9370 8770 9610
rect 9010 9370 9100 9610
rect 9340 9370 9430 9610
rect 9670 9370 9760 9610
rect 10000 9370 10090 9610
rect 10330 9370 10420 9610
rect 10660 9370 10750 9610
rect 10990 9370 11080 9610
rect 11320 9370 11410 9610
rect 11650 9370 11740 9610
rect 11980 9370 12070 9610
rect 12310 9370 12400 9610
rect 12640 9370 12730 9610
rect 12970 9370 13060 9610
rect 13300 9370 13390 9610
rect 13630 9370 13720 9610
rect 13960 9370 14050 9610
rect 14290 9370 14380 9610
rect 14620 9370 14710 9610
rect 14950 9370 15040 9610
rect 15280 9370 15370 9610
rect 15610 9370 15700 9610
rect 15940 9370 16030 9610
rect 16270 9370 16360 9610
rect 16600 9370 16690 9610
rect 16930 9370 17020 9610
rect 17260 9370 17350 9610
rect 17590 9370 17680 9610
rect 17920 9370 18010 9610
rect 18250 9370 18340 9610
rect 18580 9370 18670 9610
rect 18910 9370 19000 9610
rect 19240 9370 19330 9610
rect 19570 9370 19880 9610
rect 7640 9280 19880 9370
rect 7640 9040 7780 9280
rect 8020 9040 8110 9280
rect 8350 9040 8440 9280
rect 8680 9040 8770 9280
rect 9010 9040 9100 9280
rect 9340 9040 9430 9280
rect 9670 9040 9760 9280
rect 10000 9040 10090 9280
rect 10330 9040 10420 9280
rect 10660 9040 10750 9280
rect 10990 9040 11080 9280
rect 11320 9040 11410 9280
rect 11650 9040 11740 9280
rect 11980 9040 12070 9280
rect 12310 9040 12400 9280
rect 12640 9040 12730 9280
rect 12970 9040 13060 9280
rect 13300 9040 13390 9280
rect 13630 9040 13720 9280
rect 13960 9040 14050 9280
rect 14290 9040 14380 9280
rect 14620 9040 14710 9280
rect 14950 9040 15040 9280
rect 15280 9040 15370 9280
rect 15610 9040 15700 9280
rect 15940 9040 16030 9280
rect 16270 9040 16360 9280
rect 16600 9040 16690 9280
rect 16930 9040 17020 9280
rect 17260 9040 17350 9280
rect 17590 9040 17680 9280
rect 17920 9040 18010 9280
rect 18250 9040 18340 9280
rect 18580 9040 18670 9280
rect 18910 9040 19000 9280
rect 19240 9040 19330 9280
rect 19570 9040 19880 9280
rect 7640 8720 19880 9040
rect 31130 7830 37830 7880
rect 31130 7590 31180 7830
rect 31420 7590 31510 7830
rect 31750 7590 31840 7830
rect 32080 7590 32170 7830
rect 32410 7590 32500 7830
rect 32740 7590 32830 7830
rect 33070 7590 33160 7830
rect 33400 7590 33490 7830
rect 33730 7590 33820 7830
rect 34060 7590 34150 7830
rect 34390 7590 34480 7830
rect 34720 7590 34810 7830
rect 35050 7590 35140 7830
rect 35380 7590 35470 7830
rect 35710 7590 35800 7830
rect 36040 7590 36130 7830
rect 36370 7590 36460 7830
rect 36700 7590 36790 7830
rect 37030 7590 37120 7830
rect 37360 7590 37450 7830
rect 37690 7590 37830 7830
rect 31130 7500 37830 7590
rect 31130 7260 31180 7500
rect 31420 7260 31510 7500
rect 31750 7260 31840 7500
rect 32080 7260 32170 7500
rect 32410 7260 32500 7500
rect 32740 7260 32830 7500
rect 33070 7260 33160 7500
rect 33400 7260 33490 7500
rect 33730 7260 33820 7500
rect 34060 7260 34150 7500
rect 34390 7260 34480 7500
rect 34720 7260 34810 7500
rect 35050 7260 35140 7500
rect 35380 7260 35470 7500
rect 35710 7260 35800 7500
rect 36040 7260 36130 7500
rect 36370 7260 36460 7500
rect 36700 7260 36790 7500
rect 37030 7260 37120 7500
rect 37360 7260 37450 7500
rect 37690 7260 37830 7500
rect 31130 7170 37830 7260
rect 31130 6930 31180 7170
rect 31420 6930 31510 7170
rect 31750 6930 31840 7170
rect 32080 6930 32170 7170
rect 32410 6930 32500 7170
rect 32740 6930 32830 7170
rect 33070 6930 33160 7170
rect 33400 6930 33490 7170
rect 33730 6930 33820 7170
rect 34060 6930 34150 7170
rect 34390 6930 34480 7170
rect 34720 6930 34810 7170
rect 35050 6930 35140 7170
rect 35380 6930 35470 7170
rect 35710 6930 35800 7170
rect 36040 6930 36130 7170
rect 36370 6930 36460 7170
rect 36700 6930 36790 7170
rect 37030 6930 37120 7170
rect 37360 6930 37450 7170
rect 37690 6930 37830 7170
rect 31130 6840 37830 6930
rect 31130 6600 31180 6840
rect 31420 6600 31510 6840
rect 31750 6600 31840 6840
rect 32080 6600 32170 6840
rect 32410 6600 32500 6840
rect 32740 6600 32830 6840
rect 33070 6600 33160 6840
rect 33400 6600 33490 6840
rect 33730 6600 33820 6840
rect 34060 6600 34150 6840
rect 34390 6600 34480 6840
rect 34720 6600 34810 6840
rect 35050 6600 35140 6840
rect 35380 6600 35470 6840
rect 35710 6600 35800 6840
rect 36040 6600 36130 6840
rect 36370 6600 36460 6840
rect 36700 6600 36790 6840
rect 37030 6600 37120 6840
rect 37360 6600 37450 6840
rect 37690 6600 37830 6840
rect 31130 6510 37830 6600
rect 31130 6270 31180 6510
rect 31420 6270 31510 6510
rect 31750 6270 31840 6510
rect 32080 6270 32170 6510
rect 32410 6270 32500 6510
rect 32740 6270 32830 6510
rect 33070 6270 33160 6510
rect 33400 6270 33490 6510
rect 33730 6270 33820 6510
rect 34060 6270 34150 6510
rect 34390 6270 34480 6510
rect 34720 6270 34810 6510
rect 35050 6270 35140 6510
rect 35380 6270 35470 6510
rect 35710 6270 35800 6510
rect 36040 6270 36130 6510
rect 36370 6270 36460 6510
rect 36700 6270 36790 6510
rect 37030 6270 37120 6510
rect 37360 6270 37450 6510
rect 37690 6270 37830 6510
rect 31130 6180 37830 6270
rect 31130 5940 31180 6180
rect 31420 5940 31510 6180
rect 31750 5940 31840 6180
rect 32080 5940 32170 6180
rect 32410 5940 32500 6180
rect 32740 5940 32830 6180
rect 33070 5940 33160 6180
rect 33400 5940 33490 6180
rect 33730 5940 33820 6180
rect 34060 5940 34150 6180
rect 34390 5940 34480 6180
rect 34720 5940 34810 6180
rect 35050 5940 35140 6180
rect 35380 5940 35470 6180
rect 35710 5940 35800 6180
rect 36040 5940 36130 6180
rect 36370 5940 36460 6180
rect 36700 5940 36790 6180
rect 37030 5940 37120 6180
rect 37360 5940 37450 6180
rect 37690 5940 37830 6180
rect 31130 5850 37830 5940
rect 31130 5610 31180 5850
rect 31420 5610 31510 5850
rect 31750 5610 31840 5850
rect 32080 5610 32170 5850
rect 32410 5610 32500 5850
rect 32740 5610 32830 5850
rect 33070 5610 33160 5850
rect 33400 5610 33490 5850
rect 33730 5610 33820 5850
rect 34060 5610 34150 5850
rect 34390 5610 34480 5850
rect 34720 5610 34810 5850
rect 35050 5610 35140 5850
rect 35380 5610 35470 5850
rect 35710 5610 35800 5850
rect 36040 5610 36130 5850
rect 36370 5610 36460 5850
rect 36700 5610 36790 5850
rect 37030 5610 37120 5850
rect 37360 5610 37450 5850
rect 37690 5610 37830 5850
rect 31130 5520 37830 5610
rect 31130 5280 31180 5520
rect 31420 5280 31510 5520
rect 31750 5280 31840 5520
rect 32080 5280 32170 5520
rect 32410 5280 32500 5520
rect 32740 5280 32830 5520
rect 33070 5280 33160 5520
rect 33400 5280 33490 5520
rect 33730 5280 33820 5520
rect 34060 5280 34150 5520
rect 34390 5280 34480 5520
rect 34720 5280 34810 5520
rect 35050 5280 35140 5520
rect 35380 5280 35470 5520
rect 35710 5280 35800 5520
rect 36040 5280 36130 5520
rect 36370 5280 36460 5520
rect 36700 5280 36790 5520
rect 37030 5280 37120 5520
rect 37360 5280 37450 5520
rect 37690 5280 37830 5520
rect 31130 5190 37830 5280
rect 31130 4950 31180 5190
rect 31420 4950 31510 5190
rect 31750 4950 31840 5190
rect 32080 4950 32170 5190
rect 32410 4950 32500 5190
rect 32740 4950 32830 5190
rect 33070 4950 33160 5190
rect 33400 4950 33490 5190
rect 33730 4950 33820 5190
rect 34060 4950 34150 5190
rect 34390 4950 34480 5190
rect 34720 4950 34810 5190
rect 35050 4950 35140 5190
rect 35380 4950 35470 5190
rect 35710 4950 35800 5190
rect 36040 4950 36130 5190
rect 36370 4950 36460 5190
rect 36700 4950 36790 5190
rect 37030 4950 37120 5190
rect 37360 4950 37450 5190
rect 37690 4950 37830 5190
rect 31130 4860 37830 4950
rect 31130 4620 31180 4860
rect 31420 4620 31510 4860
rect 31750 4620 31840 4860
rect 32080 4620 32170 4860
rect 32410 4620 32500 4860
rect 32740 4620 32830 4860
rect 33070 4620 33160 4860
rect 33400 4620 33490 4860
rect 33730 4620 33820 4860
rect 34060 4620 34150 4860
rect 34390 4620 34480 4860
rect 34720 4620 34810 4860
rect 35050 4620 35140 4860
rect 35380 4620 35470 4860
rect 35710 4620 35800 4860
rect 36040 4620 36130 4860
rect 36370 4620 36460 4860
rect 36700 4620 36790 4860
rect 37030 4620 37120 4860
rect 37360 4620 37450 4860
rect 37690 4620 37830 4860
rect 31130 4530 37830 4620
rect 31130 4290 31180 4530
rect 31420 4290 31510 4530
rect 31750 4290 31840 4530
rect 32080 4290 32170 4530
rect 32410 4290 32500 4530
rect 32740 4290 32830 4530
rect 33070 4290 33160 4530
rect 33400 4290 33490 4530
rect 33730 4290 33820 4530
rect 34060 4290 34150 4530
rect 34390 4290 34480 4530
rect 34720 4290 34810 4530
rect 35050 4290 35140 4530
rect 35380 4290 35470 4530
rect 35710 4290 35800 4530
rect 36040 4290 36130 4530
rect 36370 4290 36460 4530
rect 36700 4290 36790 4530
rect 37030 4290 37120 4530
rect 37360 4290 37450 4530
rect 37690 4290 37830 4530
rect 31130 4200 37830 4290
rect 31130 3960 31180 4200
rect 31420 3960 31510 4200
rect 31750 3960 31840 4200
rect 32080 3960 32170 4200
rect 32410 3960 32500 4200
rect 32740 3960 32830 4200
rect 33070 3960 33160 4200
rect 33400 3960 33490 4200
rect 33730 3960 33820 4200
rect 34060 3960 34150 4200
rect 34390 3960 34480 4200
rect 34720 3960 34810 4200
rect 35050 3960 35140 4200
rect 35380 3960 35470 4200
rect 35710 3960 35800 4200
rect 36040 3960 36130 4200
rect 36370 3960 36460 4200
rect 36700 3960 36790 4200
rect 37030 3960 37120 4200
rect 37360 3960 37450 4200
rect 37690 3960 37830 4200
rect 31130 3870 37830 3960
rect 31130 3630 31180 3870
rect 31420 3630 31510 3870
rect 31750 3630 31840 3870
rect 32080 3630 32170 3870
rect 32410 3630 32500 3870
rect 32740 3630 32830 3870
rect 33070 3630 33160 3870
rect 33400 3630 33490 3870
rect 33730 3630 33820 3870
rect 34060 3630 34150 3870
rect 34390 3630 34480 3870
rect 34720 3630 34810 3870
rect 35050 3630 35140 3870
rect 35380 3630 35470 3870
rect 35710 3630 35800 3870
rect 36040 3630 36130 3870
rect 36370 3630 36460 3870
rect 36700 3630 36790 3870
rect 37030 3630 37120 3870
rect 37360 3630 37450 3870
rect 37690 3630 37830 3870
rect 31130 3540 37830 3630
rect 31130 3300 31180 3540
rect 31420 3300 31510 3540
rect 31750 3300 31840 3540
rect 32080 3300 32170 3540
rect 32410 3300 32500 3540
rect 32740 3300 32830 3540
rect 33070 3300 33160 3540
rect 33400 3300 33490 3540
rect 33730 3300 33820 3540
rect 34060 3300 34150 3540
rect 34390 3300 34480 3540
rect 34720 3300 34810 3540
rect 35050 3300 35140 3540
rect 35380 3300 35470 3540
rect 35710 3300 35800 3540
rect 36040 3300 36130 3540
rect 36370 3300 36460 3540
rect 36700 3300 36790 3540
rect 37030 3300 37120 3540
rect 37360 3300 37450 3540
rect 37690 3300 37830 3540
rect 31130 3210 37830 3300
rect 31130 2970 31180 3210
rect 31420 2970 31510 3210
rect 31750 2970 31840 3210
rect 32080 2970 32170 3210
rect 32410 2970 32500 3210
rect 32740 2970 32830 3210
rect 33070 2970 33160 3210
rect 33400 2970 33490 3210
rect 33730 2970 33820 3210
rect 34060 2970 34150 3210
rect 34390 2970 34480 3210
rect 34720 2970 34810 3210
rect 35050 2970 35140 3210
rect 35380 2970 35470 3210
rect 35710 2970 35800 3210
rect 36040 2970 36130 3210
rect 36370 2970 36460 3210
rect 36700 2970 36790 3210
rect 37030 2970 37120 3210
rect 37360 2970 37450 3210
rect 37690 2970 37830 3210
rect 31130 2880 37830 2970
rect 31130 2640 31180 2880
rect 31420 2640 31510 2880
rect 31750 2640 31840 2880
rect 32080 2640 32170 2880
rect 32410 2640 32500 2880
rect 32740 2640 32830 2880
rect 33070 2640 33160 2880
rect 33400 2640 33490 2880
rect 33730 2640 33820 2880
rect 34060 2640 34150 2880
rect 34390 2640 34480 2880
rect 34720 2640 34810 2880
rect 35050 2640 35140 2880
rect 35380 2640 35470 2880
rect 35710 2640 35800 2880
rect 36040 2640 36130 2880
rect 36370 2640 36460 2880
rect 36700 2640 36790 2880
rect 37030 2640 37120 2880
rect 37360 2640 37450 2880
rect 37690 2640 37830 2880
rect 31130 2550 37830 2640
rect 31130 2310 31180 2550
rect 31420 2310 31510 2550
rect 31750 2310 31840 2550
rect 32080 2310 32170 2550
rect 32410 2310 32500 2550
rect 32740 2310 32830 2550
rect 33070 2310 33160 2550
rect 33400 2310 33490 2550
rect 33730 2310 33820 2550
rect 34060 2310 34150 2550
rect 34390 2310 34480 2550
rect 34720 2310 34810 2550
rect 35050 2310 35140 2550
rect 35380 2310 35470 2550
rect 35710 2310 35800 2550
rect 36040 2310 36130 2550
rect 36370 2310 36460 2550
rect 36700 2310 36790 2550
rect 37030 2310 37120 2550
rect 37360 2310 37450 2550
rect 37690 2310 37830 2550
rect 31130 2220 37830 2310
rect 31130 1980 31180 2220
rect 31420 1980 31510 2220
rect 31750 1980 31840 2220
rect 32080 1980 32170 2220
rect 32410 1980 32500 2220
rect 32740 1980 32830 2220
rect 33070 1980 33160 2220
rect 33400 1980 33490 2220
rect 33730 1980 33820 2220
rect 34060 1980 34150 2220
rect 34390 1980 34480 2220
rect 34720 1980 34810 2220
rect 35050 1980 35140 2220
rect 35380 1980 35470 2220
rect 35710 1980 35800 2220
rect 36040 1980 36130 2220
rect 36370 1980 36460 2220
rect 36700 1980 36790 2220
rect 37030 1980 37120 2220
rect 37360 1980 37450 2220
rect 37690 1980 37830 2220
rect 31130 1890 37830 1980
rect 31130 1650 31180 1890
rect 31420 1650 31510 1890
rect 31750 1650 31840 1890
rect 32080 1650 32170 1890
rect 32410 1650 32500 1890
rect 32740 1650 32830 1890
rect 33070 1650 33160 1890
rect 33400 1650 33490 1890
rect 33730 1650 33820 1890
rect 34060 1650 34150 1890
rect 34390 1650 34480 1890
rect 34720 1650 34810 1890
rect 35050 1650 35140 1890
rect 35380 1650 35470 1890
rect 35710 1650 35800 1890
rect 36040 1650 36130 1890
rect 36370 1650 36460 1890
rect 36700 1650 36790 1890
rect 37030 1650 37120 1890
rect 37360 1650 37450 1890
rect 37690 1650 37830 1890
rect 31130 1560 37830 1650
rect 31130 1320 31180 1560
rect 31420 1320 31510 1560
rect 31750 1320 31840 1560
rect 32080 1320 32170 1560
rect 32410 1320 32500 1560
rect 32740 1320 32830 1560
rect 33070 1320 33160 1560
rect 33400 1320 33490 1560
rect 33730 1320 33820 1560
rect 34060 1320 34150 1560
rect 34390 1320 34480 1560
rect 34720 1320 34810 1560
rect 35050 1320 35140 1560
rect 35380 1320 35470 1560
rect 35710 1320 35800 1560
rect 36040 1320 36130 1560
rect 36370 1320 36460 1560
rect 36700 1320 36790 1560
rect 37030 1320 37120 1560
rect 37360 1320 37450 1560
rect 37690 1320 37830 1560
rect 31130 1180 37830 1320
rect 31130 230 37830 280
rect 31130 -10 31180 230
rect 31420 -10 31510 230
rect 31750 -10 31840 230
rect 32080 -10 32170 230
rect 32410 -10 32500 230
rect 32740 -10 32830 230
rect 33070 -10 33160 230
rect 33400 -10 33490 230
rect 33730 -10 33820 230
rect 34060 -10 34150 230
rect 34390 -10 34480 230
rect 34720 -10 34810 230
rect 35050 -10 35140 230
rect 35380 -10 35470 230
rect 35710 -10 35800 230
rect 36040 -10 36130 230
rect 36370 -10 36460 230
rect 36700 -10 36790 230
rect 37030 -10 37120 230
rect 37360 -10 37450 230
rect 37690 -10 37830 230
rect 31130 -100 37830 -10
rect 31130 -340 31180 -100
rect 31420 -340 31510 -100
rect 31750 -340 31840 -100
rect 32080 -340 32170 -100
rect 32410 -340 32500 -100
rect 32740 -340 32830 -100
rect 33070 -340 33160 -100
rect 33400 -340 33490 -100
rect 33730 -340 33820 -100
rect 34060 -340 34150 -100
rect 34390 -340 34480 -100
rect 34720 -340 34810 -100
rect 35050 -340 35140 -100
rect 35380 -340 35470 -100
rect 35710 -340 35800 -100
rect 36040 -340 36130 -100
rect 36370 -340 36460 -100
rect 36700 -340 36790 -100
rect 37030 -340 37120 -100
rect 37360 -340 37450 -100
rect 37690 -340 37830 -100
rect 31130 -430 37830 -340
rect 31130 -670 31180 -430
rect 31420 -670 31510 -430
rect 31750 -670 31840 -430
rect 32080 -670 32170 -430
rect 32410 -670 32500 -430
rect 32740 -670 32830 -430
rect 33070 -670 33160 -430
rect 33400 -670 33490 -430
rect 33730 -670 33820 -430
rect 34060 -670 34150 -430
rect 34390 -670 34480 -430
rect 34720 -670 34810 -430
rect 35050 -670 35140 -430
rect 35380 -670 35470 -430
rect 35710 -670 35800 -430
rect 36040 -670 36130 -430
rect 36370 -670 36460 -430
rect 36700 -670 36790 -430
rect 37030 -670 37120 -430
rect 37360 -670 37450 -430
rect 37690 -670 37830 -430
rect 31130 -760 37830 -670
rect 31130 -1000 31180 -760
rect 31420 -1000 31510 -760
rect 31750 -1000 31840 -760
rect 32080 -1000 32170 -760
rect 32410 -1000 32500 -760
rect 32740 -1000 32830 -760
rect 33070 -1000 33160 -760
rect 33400 -1000 33490 -760
rect 33730 -1000 33820 -760
rect 34060 -1000 34150 -760
rect 34390 -1000 34480 -760
rect 34720 -1000 34810 -760
rect 35050 -1000 35140 -760
rect 35380 -1000 35470 -760
rect 35710 -1000 35800 -760
rect 36040 -1000 36130 -760
rect 36370 -1000 36460 -760
rect 36700 -1000 36790 -760
rect 37030 -1000 37120 -760
rect 37360 -1000 37450 -760
rect 37690 -1000 37830 -760
rect 31130 -1090 37830 -1000
rect 31130 -1330 31180 -1090
rect 31420 -1330 31510 -1090
rect 31750 -1330 31840 -1090
rect 32080 -1330 32170 -1090
rect 32410 -1330 32500 -1090
rect 32740 -1330 32830 -1090
rect 33070 -1330 33160 -1090
rect 33400 -1330 33490 -1090
rect 33730 -1330 33820 -1090
rect 34060 -1330 34150 -1090
rect 34390 -1330 34480 -1090
rect 34720 -1330 34810 -1090
rect 35050 -1330 35140 -1090
rect 35380 -1330 35470 -1090
rect 35710 -1330 35800 -1090
rect 36040 -1330 36130 -1090
rect 36370 -1330 36460 -1090
rect 36700 -1330 36790 -1090
rect 37030 -1330 37120 -1090
rect 37360 -1330 37450 -1090
rect 37690 -1330 37830 -1090
rect 31130 -1420 37830 -1330
rect 31130 -1660 31180 -1420
rect 31420 -1660 31510 -1420
rect 31750 -1660 31840 -1420
rect 32080 -1660 32170 -1420
rect 32410 -1660 32500 -1420
rect 32740 -1660 32830 -1420
rect 33070 -1660 33160 -1420
rect 33400 -1660 33490 -1420
rect 33730 -1660 33820 -1420
rect 34060 -1660 34150 -1420
rect 34390 -1660 34480 -1420
rect 34720 -1660 34810 -1420
rect 35050 -1660 35140 -1420
rect 35380 -1660 35470 -1420
rect 35710 -1660 35800 -1420
rect 36040 -1660 36130 -1420
rect 36370 -1660 36460 -1420
rect 36700 -1660 36790 -1420
rect 37030 -1660 37120 -1420
rect 37360 -1660 37450 -1420
rect 37690 -1660 37830 -1420
rect 31130 -1750 37830 -1660
rect 31130 -1990 31180 -1750
rect 31420 -1990 31510 -1750
rect 31750 -1990 31840 -1750
rect 32080 -1990 32170 -1750
rect 32410 -1990 32500 -1750
rect 32740 -1990 32830 -1750
rect 33070 -1990 33160 -1750
rect 33400 -1990 33490 -1750
rect 33730 -1990 33820 -1750
rect 34060 -1990 34150 -1750
rect 34390 -1990 34480 -1750
rect 34720 -1990 34810 -1750
rect 35050 -1990 35140 -1750
rect 35380 -1990 35470 -1750
rect 35710 -1990 35800 -1750
rect 36040 -1990 36130 -1750
rect 36370 -1990 36460 -1750
rect 36700 -1990 36790 -1750
rect 37030 -1990 37120 -1750
rect 37360 -1990 37450 -1750
rect 37690 -1990 37830 -1750
rect 31130 -2080 37830 -1990
rect 31130 -2320 31180 -2080
rect 31420 -2320 31510 -2080
rect 31750 -2320 31840 -2080
rect 32080 -2320 32170 -2080
rect 32410 -2320 32500 -2080
rect 32740 -2320 32830 -2080
rect 33070 -2320 33160 -2080
rect 33400 -2320 33490 -2080
rect 33730 -2320 33820 -2080
rect 34060 -2320 34150 -2080
rect 34390 -2320 34480 -2080
rect 34720 -2320 34810 -2080
rect 35050 -2320 35140 -2080
rect 35380 -2320 35470 -2080
rect 35710 -2320 35800 -2080
rect 36040 -2320 36130 -2080
rect 36370 -2320 36460 -2080
rect 36700 -2320 36790 -2080
rect 37030 -2320 37120 -2080
rect 37360 -2320 37450 -2080
rect 37690 -2320 37830 -2080
rect 31130 -2410 37830 -2320
rect 31130 -2650 31180 -2410
rect 31420 -2650 31510 -2410
rect 31750 -2650 31840 -2410
rect 32080 -2650 32170 -2410
rect 32410 -2650 32500 -2410
rect 32740 -2650 32830 -2410
rect 33070 -2650 33160 -2410
rect 33400 -2650 33490 -2410
rect 33730 -2650 33820 -2410
rect 34060 -2650 34150 -2410
rect 34390 -2650 34480 -2410
rect 34720 -2650 34810 -2410
rect 35050 -2650 35140 -2410
rect 35380 -2650 35470 -2410
rect 35710 -2650 35800 -2410
rect 36040 -2650 36130 -2410
rect 36370 -2650 36460 -2410
rect 36700 -2650 36790 -2410
rect 37030 -2650 37120 -2410
rect 37360 -2650 37450 -2410
rect 37690 -2650 37830 -2410
rect 31130 -2740 37830 -2650
rect 31130 -2980 31180 -2740
rect 31420 -2980 31510 -2740
rect 31750 -2980 31840 -2740
rect 32080 -2980 32170 -2740
rect 32410 -2980 32500 -2740
rect 32740 -2980 32830 -2740
rect 33070 -2980 33160 -2740
rect 33400 -2980 33490 -2740
rect 33730 -2980 33820 -2740
rect 34060 -2980 34150 -2740
rect 34390 -2980 34480 -2740
rect 34720 -2980 34810 -2740
rect 35050 -2980 35140 -2740
rect 35380 -2980 35470 -2740
rect 35710 -2980 35800 -2740
rect 36040 -2980 36130 -2740
rect 36370 -2980 36460 -2740
rect 36700 -2980 36790 -2740
rect 37030 -2980 37120 -2740
rect 37360 -2980 37450 -2740
rect 37690 -2980 37830 -2740
rect 31130 -3070 37830 -2980
rect 31130 -3310 31180 -3070
rect 31420 -3310 31510 -3070
rect 31750 -3310 31840 -3070
rect 32080 -3310 32170 -3070
rect 32410 -3310 32500 -3070
rect 32740 -3310 32830 -3070
rect 33070 -3310 33160 -3070
rect 33400 -3310 33490 -3070
rect 33730 -3310 33820 -3070
rect 34060 -3310 34150 -3070
rect 34390 -3310 34480 -3070
rect 34720 -3310 34810 -3070
rect 35050 -3310 35140 -3070
rect 35380 -3310 35470 -3070
rect 35710 -3310 35800 -3070
rect 36040 -3310 36130 -3070
rect 36370 -3310 36460 -3070
rect 36700 -3310 36790 -3070
rect 37030 -3310 37120 -3070
rect 37360 -3310 37450 -3070
rect 37690 -3310 37830 -3070
rect 31130 -3400 37830 -3310
rect 31130 -3640 31180 -3400
rect 31420 -3640 31510 -3400
rect 31750 -3640 31840 -3400
rect 32080 -3640 32170 -3400
rect 32410 -3640 32500 -3400
rect 32740 -3640 32830 -3400
rect 33070 -3640 33160 -3400
rect 33400 -3640 33490 -3400
rect 33730 -3640 33820 -3400
rect 34060 -3640 34150 -3400
rect 34390 -3640 34480 -3400
rect 34720 -3640 34810 -3400
rect 35050 -3640 35140 -3400
rect 35380 -3640 35470 -3400
rect 35710 -3640 35800 -3400
rect 36040 -3640 36130 -3400
rect 36370 -3640 36460 -3400
rect 36700 -3640 36790 -3400
rect 37030 -3640 37120 -3400
rect 37360 -3640 37450 -3400
rect 37690 -3640 37830 -3400
rect 31130 -3730 37830 -3640
rect 31130 -3970 31180 -3730
rect 31420 -3970 31510 -3730
rect 31750 -3970 31840 -3730
rect 32080 -3970 32170 -3730
rect 32410 -3970 32500 -3730
rect 32740 -3970 32830 -3730
rect 33070 -3970 33160 -3730
rect 33400 -3970 33490 -3730
rect 33730 -3970 33820 -3730
rect 34060 -3970 34150 -3730
rect 34390 -3970 34480 -3730
rect 34720 -3970 34810 -3730
rect 35050 -3970 35140 -3730
rect 35380 -3970 35470 -3730
rect 35710 -3970 35800 -3730
rect 36040 -3970 36130 -3730
rect 36370 -3970 36460 -3730
rect 36700 -3970 36790 -3730
rect 37030 -3970 37120 -3730
rect 37360 -3970 37450 -3730
rect 37690 -3970 37830 -3730
rect 31130 -4060 37830 -3970
rect 31130 -4300 31180 -4060
rect 31420 -4300 31510 -4060
rect 31750 -4300 31840 -4060
rect 32080 -4300 32170 -4060
rect 32410 -4300 32500 -4060
rect 32740 -4300 32830 -4060
rect 33070 -4300 33160 -4060
rect 33400 -4300 33490 -4060
rect 33730 -4300 33820 -4060
rect 34060 -4300 34150 -4060
rect 34390 -4300 34480 -4060
rect 34720 -4300 34810 -4060
rect 35050 -4300 35140 -4060
rect 35380 -4300 35470 -4060
rect 35710 -4300 35800 -4060
rect 36040 -4300 36130 -4060
rect 36370 -4300 36460 -4060
rect 36700 -4300 36790 -4060
rect 37030 -4300 37120 -4060
rect 37360 -4300 37450 -4060
rect 37690 -4300 37830 -4060
rect 31130 -4390 37830 -4300
rect 31130 -4630 31180 -4390
rect 31420 -4630 31510 -4390
rect 31750 -4630 31840 -4390
rect 32080 -4630 32170 -4390
rect 32410 -4630 32500 -4390
rect 32740 -4630 32830 -4390
rect 33070 -4630 33160 -4390
rect 33400 -4630 33490 -4390
rect 33730 -4630 33820 -4390
rect 34060 -4630 34150 -4390
rect 34390 -4630 34480 -4390
rect 34720 -4630 34810 -4390
rect 35050 -4630 35140 -4390
rect 35380 -4630 35470 -4390
rect 35710 -4630 35800 -4390
rect 36040 -4630 36130 -4390
rect 36370 -4630 36460 -4390
rect 36700 -4630 36790 -4390
rect 37030 -4630 37120 -4390
rect 37360 -4630 37450 -4390
rect 37690 -4630 37830 -4390
rect -1320 -4840 230 -4660
rect -1320 -5080 -1180 -4840
rect -940 -5080 -850 -4840
rect -610 -5080 -520 -4840
rect -280 -5080 -190 -4840
rect 50 -5080 230 -4840
rect -1320 -5170 230 -5080
rect -1320 -5410 -1180 -5170
rect -940 -5410 -850 -5170
rect -610 -5410 -520 -5170
rect -280 -5410 -190 -5170
rect 50 -5410 230 -5170
rect -1320 -5500 230 -5410
rect -1320 -5740 -1180 -5500
rect -940 -5740 -850 -5500
rect -610 -5740 -520 -5500
rect -280 -5740 -190 -5500
rect 50 -5740 230 -5500
rect -1320 -5830 230 -5740
rect -1320 -6070 -1180 -5830
rect -940 -6070 -850 -5830
rect -610 -6070 -520 -5830
rect -280 -6070 -190 -5830
rect 50 -6070 230 -5830
rect -1320 -6210 230 -6070
rect 14550 -4840 16100 -4660
rect 14550 -5080 14730 -4840
rect 14970 -5080 15060 -4840
rect 15300 -5080 15390 -4840
rect 15630 -5080 15720 -4840
rect 15960 -5080 16100 -4840
rect 14550 -5170 16100 -5080
rect 14550 -5410 14730 -5170
rect 14970 -5410 15060 -5170
rect 15300 -5410 15390 -5170
rect 15630 -5410 15720 -5170
rect 15960 -5410 16100 -5170
rect 14550 -5500 16100 -5410
rect 14550 -5740 14730 -5500
rect 14970 -5740 15060 -5500
rect 15300 -5740 15390 -5500
rect 15630 -5740 15720 -5500
rect 15960 -5740 16100 -5500
rect 14550 -5830 16100 -5740
rect 14550 -6070 14730 -5830
rect 14970 -6070 15060 -5830
rect 15300 -6070 15390 -5830
rect 15630 -6070 15720 -5830
rect 15960 -6070 16100 -5830
rect 14550 -6210 16100 -6070
rect 31130 -4720 37830 -4630
rect 31130 -4960 31180 -4720
rect 31420 -4960 31510 -4720
rect 31750 -4960 31840 -4720
rect 32080 -4960 32170 -4720
rect 32410 -4960 32500 -4720
rect 32740 -4960 32830 -4720
rect 33070 -4960 33160 -4720
rect 33400 -4960 33490 -4720
rect 33730 -4960 33820 -4720
rect 34060 -4960 34150 -4720
rect 34390 -4960 34480 -4720
rect 34720 -4960 34810 -4720
rect 35050 -4960 35140 -4720
rect 35380 -4960 35470 -4720
rect 35710 -4960 35800 -4720
rect 36040 -4960 36130 -4720
rect 36370 -4960 36460 -4720
rect 36700 -4960 36790 -4720
rect 37030 -4960 37120 -4720
rect 37360 -4960 37450 -4720
rect 37690 -4960 37830 -4720
rect 31130 -5050 37830 -4960
rect 31130 -5290 31180 -5050
rect 31420 -5290 31510 -5050
rect 31750 -5290 31840 -5050
rect 32080 -5290 32170 -5050
rect 32410 -5290 32500 -5050
rect 32740 -5290 32830 -5050
rect 33070 -5290 33160 -5050
rect 33400 -5290 33490 -5050
rect 33730 -5290 33820 -5050
rect 34060 -5290 34150 -5050
rect 34390 -5290 34480 -5050
rect 34720 -5290 34810 -5050
rect 35050 -5290 35140 -5050
rect 35380 -5290 35470 -5050
rect 35710 -5290 35800 -5050
rect 36040 -5290 36130 -5050
rect 36370 -5290 36460 -5050
rect 36700 -5290 36790 -5050
rect 37030 -5290 37120 -5050
rect 37360 -5290 37450 -5050
rect 37690 -5290 37830 -5050
rect 31130 -5380 37830 -5290
rect 31130 -5620 31180 -5380
rect 31420 -5620 31510 -5380
rect 31750 -5620 31840 -5380
rect 32080 -5620 32170 -5380
rect 32410 -5620 32500 -5380
rect 32740 -5620 32830 -5380
rect 33070 -5620 33160 -5380
rect 33400 -5620 33490 -5380
rect 33730 -5620 33820 -5380
rect 34060 -5620 34150 -5380
rect 34390 -5620 34480 -5380
rect 34720 -5620 34810 -5380
rect 35050 -5620 35140 -5380
rect 35380 -5620 35470 -5380
rect 35710 -5620 35800 -5380
rect 36040 -5620 36130 -5380
rect 36370 -5620 36460 -5380
rect 36700 -5620 36790 -5380
rect 37030 -5620 37120 -5380
rect 37360 -5620 37450 -5380
rect 37690 -5620 37830 -5380
rect 31130 -5710 37830 -5620
rect 31130 -5950 31180 -5710
rect 31420 -5950 31510 -5710
rect 31750 -5950 31840 -5710
rect 32080 -5950 32170 -5710
rect 32410 -5950 32500 -5710
rect 32740 -5950 32830 -5710
rect 33070 -5950 33160 -5710
rect 33400 -5950 33490 -5710
rect 33730 -5950 33820 -5710
rect 34060 -5950 34150 -5710
rect 34390 -5950 34480 -5710
rect 34720 -5950 34810 -5710
rect 35050 -5950 35140 -5710
rect 35380 -5950 35470 -5710
rect 35710 -5950 35800 -5710
rect 36040 -5950 36130 -5710
rect 36370 -5950 36460 -5710
rect 36700 -5950 36790 -5710
rect 37030 -5950 37120 -5710
rect 37360 -5950 37450 -5710
rect 37690 -5950 37830 -5710
rect 31130 -6040 37830 -5950
rect 31130 -6280 31180 -6040
rect 31420 -6280 31510 -6040
rect 31750 -6280 31840 -6040
rect 32080 -6280 32170 -6040
rect 32410 -6280 32500 -6040
rect 32740 -6280 32830 -6040
rect 33070 -6280 33160 -6040
rect 33400 -6280 33490 -6040
rect 33730 -6280 33820 -6040
rect 34060 -6280 34150 -6040
rect 34390 -6280 34480 -6040
rect 34720 -6280 34810 -6040
rect 35050 -6280 35140 -6040
rect 35380 -6280 35470 -6040
rect 35710 -6280 35800 -6040
rect 36040 -6280 36130 -6040
rect 36370 -6280 36460 -6040
rect 36700 -6280 36790 -6040
rect 37030 -6280 37120 -6040
rect 37360 -6280 37450 -6040
rect 37690 -6280 37830 -6040
rect 31130 -6420 37830 -6280
<< mimcap2contact >>
rect -4670 20590 -4430 20830
rect -4340 20590 -4100 20830
rect -4010 20590 -3770 20830
rect -3680 20590 -3440 20830
rect -3350 20590 -3110 20830
rect -3020 20590 -2780 20830
rect -2690 20590 -2450 20830
rect -2360 20590 -2120 20830
rect -2030 20590 -1790 20830
rect -1700 20590 -1460 20830
rect -1370 20590 -1130 20830
rect -1040 20590 -800 20830
rect -710 20590 -470 20830
rect -380 20590 -140 20830
rect -50 20590 190 20830
rect 280 20590 520 20830
rect 610 20590 850 20830
rect 940 20590 1180 20830
rect 1270 20590 1510 20830
rect 1600 20590 1840 20830
rect 1930 20590 2170 20830
rect 2260 20590 2500 20830
rect 2590 20590 2830 20830
rect 2920 20590 3160 20830
rect 3250 20590 3490 20830
rect 3580 20590 3820 20830
rect 3910 20590 4150 20830
rect 4240 20590 4480 20830
rect 4570 20590 4810 20830
rect 4900 20590 5140 20830
rect 5230 20590 5470 20830
rect 5560 20590 5800 20830
rect 5890 20590 6130 20830
rect 6220 20590 6460 20830
rect 6550 20590 6790 20830
rect 6880 20590 7120 20830
rect -4670 20260 -4430 20500
rect -4340 20260 -4100 20500
rect -4010 20260 -3770 20500
rect -3680 20260 -3440 20500
rect -3350 20260 -3110 20500
rect -3020 20260 -2780 20500
rect -2690 20260 -2450 20500
rect -2360 20260 -2120 20500
rect -2030 20260 -1790 20500
rect -1700 20260 -1460 20500
rect -1370 20260 -1130 20500
rect -1040 20260 -800 20500
rect -710 20260 -470 20500
rect -380 20260 -140 20500
rect -50 20260 190 20500
rect 280 20260 520 20500
rect 610 20260 850 20500
rect 940 20260 1180 20500
rect 1270 20260 1510 20500
rect 1600 20260 1840 20500
rect 1930 20260 2170 20500
rect 2260 20260 2500 20500
rect 2590 20260 2830 20500
rect 2920 20260 3160 20500
rect 3250 20260 3490 20500
rect 3580 20260 3820 20500
rect 3910 20260 4150 20500
rect 4240 20260 4480 20500
rect 4570 20260 4810 20500
rect 4900 20260 5140 20500
rect 5230 20260 5470 20500
rect 5560 20260 5800 20500
rect 5890 20260 6130 20500
rect 6220 20260 6460 20500
rect 6550 20260 6790 20500
rect 6880 20260 7120 20500
rect -4670 19930 -4430 20170
rect -4340 19930 -4100 20170
rect -4010 19930 -3770 20170
rect -3680 19930 -3440 20170
rect -3350 19930 -3110 20170
rect -3020 19930 -2780 20170
rect -2690 19930 -2450 20170
rect -2360 19930 -2120 20170
rect -2030 19930 -1790 20170
rect -1700 19930 -1460 20170
rect -1370 19930 -1130 20170
rect -1040 19930 -800 20170
rect -710 19930 -470 20170
rect -380 19930 -140 20170
rect -50 19930 190 20170
rect 280 19930 520 20170
rect 610 19930 850 20170
rect 940 19930 1180 20170
rect 1270 19930 1510 20170
rect 1600 19930 1840 20170
rect 1930 19930 2170 20170
rect 2260 19930 2500 20170
rect 2590 19930 2830 20170
rect 2920 19930 3160 20170
rect 3250 19930 3490 20170
rect 3580 19930 3820 20170
rect 3910 19930 4150 20170
rect 4240 19930 4480 20170
rect 4570 19930 4810 20170
rect 4900 19930 5140 20170
rect 5230 19930 5470 20170
rect 5560 19930 5800 20170
rect 5890 19930 6130 20170
rect 6220 19930 6460 20170
rect 6550 19930 6790 20170
rect 6880 19930 7120 20170
rect -4670 19600 -4430 19840
rect -4340 19600 -4100 19840
rect -4010 19600 -3770 19840
rect -3680 19600 -3440 19840
rect -3350 19600 -3110 19840
rect -3020 19600 -2780 19840
rect -2690 19600 -2450 19840
rect -2360 19600 -2120 19840
rect -2030 19600 -1790 19840
rect -1700 19600 -1460 19840
rect -1370 19600 -1130 19840
rect -1040 19600 -800 19840
rect -710 19600 -470 19840
rect -380 19600 -140 19840
rect -50 19600 190 19840
rect 280 19600 520 19840
rect 610 19600 850 19840
rect 940 19600 1180 19840
rect 1270 19600 1510 19840
rect 1600 19600 1840 19840
rect 1930 19600 2170 19840
rect 2260 19600 2500 19840
rect 2590 19600 2830 19840
rect 2920 19600 3160 19840
rect 3250 19600 3490 19840
rect 3580 19600 3820 19840
rect 3910 19600 4150 19840
rect 4240 19600 4480 19840
rect 4570 19600 4810 19840
rect 4900 19600 5140 19840
rect 5230 19600 5470 19840
rect 5560 19600 5800 19840
rect 5890 19600 6130 19840
rect 6220 19600 6460 19840
rect 6550 19600 6790 19840
rect 6880 19600 7120 19840
rect -4670 19270 -4430 19510
rect -4340 19270 -4100 19510
rect -4010 19270 -3770 19510
rect -3680 19270 -3440 19510
rect -3350 19270 -3110 19510
rect -3020 19270 -2780 19510
rect -2690 19270 -2450 19510
rect -2360 19270 -2120 19510
rect -2030 19270 -1790 19510
rect -1700 19270 -1460 19510
rect -1370 19270 -1130 19510
rect -1040 19270 -800 19510
rect -710 19270 -470 19510
rect -380 19270 -140 19510
rect -50 19270 190 19510
rect 280 19270 520 19510
rect 610 19270 850 19510
rect 940 19270 1180 19510
rect 1270 19270 1510 19510
rect 1600 19270 1840 19510
rect 1930 19270 2170 19510
rect 2260 19270 2500 19510
rect 2590 19270 2830 19510
rect 2920 19270 3160 19510
rect 3250 19270 3490 19510
rect 3580 19270 3820 19510
rect 3910 19270 4150 19510
rect 4240 19270 4480 19510
rect 4570 19270 4810 19510
rect 4900 19270 5140 19510
rect 5230 19270 5470 19510
rect 5560 19270 5800 19510
rect 5890 19270 6130 19510
rect 6220 19270 6460 19510
rect 6550 19270 6790 19510
rect 6880 19270 7120 19510
rect -4670 18940 -4430 19180
rect -4340 18940 -4100 19180
rect -4010 18940 -3770 19180
rect -3680 18940 -3440 19180
rect -3350 18940 -3110 19180
rect -3020 18940 -2780 19180
rect -2690 18940 -2450 19180
rect -2360 18940 -2120 19180
rect -2030 18940 -1790 19180
rect -1700 18940 -1460 19180
rect -1370 18940 -1130 19180
rect -1040 18940 -800 19180
rect -710 18940 -470 19180
rect -380 18940 -140 19180
rect -50 18940 190 19180
rect 280 18940 520 19180
rect 610 18940 850 19180
rect 940 18940 1180 19180
rect 1270 18940 1510 19180
rect 1600 18940 1840 19180
rect 1930 18940 2170 19180
rect 2260 18940 2500 19180
rect 2590 18940 2830 19180
rect 2920 18940 3160 19180
rect 3250 18940 3490 19180
rect 3580 18940 3820 19180
rect 3910 18940 4150 19180
rect 4240 18940 4480 19180
rect 4570 18940 4810 19180
rect 4900 18940 5140 19180
rect 5230 18940 5470 19180
rect 5560 18940 5800 19180
rect 5890 18940 6130 19180
rect 6220 18940 6460 19180
rect 6550 18940 6790 19180
rect 6880 18940 7120 19180
rect -4670 18610 -4430 18850
rect -4340 18610 -4100 18850
rect -4010 18610 -3770 18850
rect -3680 18610 -3440 18850
rect -3350 18610 -3110 18850
rect -3020 18610 -2780 18850
rect -2690 18610 -2450 18850
rect -2360 18610 -2120 18850
rect -2030 18610 -1790 18850
rect -1700 18610 -1460 18850
rect -1370 18610 -1130 18850
rect -1040 18610 -800 18850
rect -710 18610 -470 18850
rect -380 18610 -140 18850
rect -50 18610 190 18850
rect 280 18610 520 18850
rect 610 18610 850 18850
rect 940 18610 1180 18850
rect 1270 18610 1510 18850
rect 1600 18610 1840 18850
rect 1930 18610 2170 18850
rect 2260 18610 2500 18850
rect 2590 18610 2830 18850
rect 2920 18610 3160 18850
rect 3250 18610 3490 18850
rect 3580 18610 3820 18850
rect 3910 18610 4150 18850
rect 4240 18610 4480 18850
rect 4570 18610 4810 18850
rect 4900 18610 5140 18850
rect 5230 18610 5470 18850
rect 5560 18610 5800 18850
rect 5890 18610 6130 18850
rect 6220 18610 6460 18850
rect 6550 18610 6790 18850
rect 6880 18610 7120 18850
rect -4670 18280 -4430 18520
rect -4340 18280 -4100 18520
rect -4010 18280 -3770 18520
rect -3680 18280 -3440 18520
rect -3350 18280 -3110 18520
rect -3020 18280 -2780 18520
rect -2690 18280 -2450 18520
rect -2360 18280 -2120 18520
rect -2030 18280 -1790 18520
rect -1700 18280 -1460 18520
rect -1370 18280 -1130 18520
rect -1040 18280 -800 18520
rect -710 18280 -470 18520
rect -380 18280 -140 18520
rect -50 18280 190 18520
rect 280 18280 520 18520
rect 610 18280 850 18520
rect 940 18280 1180 18520
rect 1270 18280 1510 18520
rect 1600 18280 1840 18520
rect 1930 18280 2170 18520
rect 2260 18280 2500 18520
rect 2590 18280 2830 18520
rect 2920 18280 3160 18520
rect 3250 18280 3490 18520
rect 3580 18280 3820 18520
rect 3910 18280 4150 18520
rect 4240 18280 4480 18520
rect 4570 18280 4810 18520
rect 4900 18280 5140 18520
rect 5230 18280 5470 18520
rect 5560 18280 5800 18520
rect 5890 18280 6130 18520
rect 6220 18280 6460 18520
rect 6550 18280 6790 18520
rect 6880 18280 7120 18520
rect -4670 17950 -4430 18190
rect -4340 17950 -4100 18190
rect -4010 17950 -3770 18190
rect -3680 17950 -3440 18190
rect -3350 17950 -3110 18190
rect -3020 17950 -2780 18190
rect -2690 17950 -2450 18190
rect -2360 17950 -2120 18190
rect -2030 17950 -1790 18190
rect -1700 17950 -1460 18190
rect -1370 17950 -1130 18190
rect -1040 17950 -800 18190
rect -710 17950 -470 18190
rect -380 17950 -140 18190
rect -50 17950 190 18190
rect 280 17950 520 18190
rect 610 17950 850 18190
rect 940 17950 1180 18190
rect 1270 17950 1510 18190
rect 1600 17950 1840 18190
rect 1930 17950 2170 18190
rect 2260 17950 2500 18190
rect 2590 17950 2830 18190
rect 2920 17950 3160 18190
rect 3250 17950 3490 18190
rect 3580 17950 3820 18190
rect 3910 17950 4150 18190
rect 4240 17950 4480 18190
rect 4570 17950 4810 18190
rect 4900 17950 5140 18190
rect 5230 17950 5470 18190
rect 5560 17950 5800 18190
rect 5890 17950 6130 18190
rect 6220 17950 6460 18190
rect 6550 17950 6790 18190
rect 6880 17950 7120 18190
rect -4670 17620 -4430 17860
rect -4340 17620 -4100 17860
rect -4010 17620 -3770 17860
rect -3680 17620 -3440 17860
rect -3350 17620 -3110 17860
rect -3020 17620 -2780 17860
rect -2690 17620 -2450 17860
rect -2360 17620 -2120 17860
rect -2030 17620 -1790 17860
rect -1700 17620 -1460 17860
rect -1370 17620 -1130 17860
rect -1040 17620 -800 17860
rect -710 17620 -470 17860
rect -380 17620 -140 17860
rect -50 17620 190 17860
rect 280 17620 520 17860
rect 610 17620 850 17860
rect 940 17620 1180 17860
rect 1270 17620 1510 17860
rect 1600 17620 1840 17860
rect 1930 17620 2170 17860
rect 2260 17620 2500 17860
rect 2590 17620 2830 17860
rect 2920 17620 3160 17860
rect 3250 17620 3490 17860
rect 3580 17620 3820 17860
rect 3910 17620 4150 17860
rect 4240 17620 4480 17860
rect 4570 17620 4810 17860
rect 4900 17620 5140 17860
rect 5230 17620 5470 17860
rect 5560 17620 5800 17860
rect 5890 17620 6130 17860
rect 6220 17620 6460 17860
rect 6550 17620 6790 17860
rect 6880 17620 7120 17860
rect -4670 17290 -4430 17530
rect -4340 17290 -4100 17530
rect -4010 17290 -3770 17530
rect -3680 17290 -3440 17530
rect -3350 17290 -3110 17530
rect -3020 17290 -2780 17530
rect -2690 17290 -2450 17530
rect -2360 17290 -2120 17530
rect -2030 17290 -1790 17530
rect -1700 17290 -1460 17530
rect -1370 17290 -1130 17530
rect -1040 17290 -800 17530
rect -710 17290 -470 17530
rect -380 17290 -140 17530
rect -50 17290 190 17530
rect 280 17290 520 17530
rect 610 17290 850 17530
rect 940 17290 1180 17530
rect 1270 17290 1510 17530
rect 1600 17290 1840 17530
rect 1930 17290 2170 17530
rect 2260 17290 2500 17530
rect 2590 17290 2830 17530
rect 2920 17290 3160 17530
rect 3250 17290 3490 17530
rect 3580 17290 3820 17530
rect 3910 17290 4150 17530
rect 4240 17290 4480 17530
rect 4570 17290 4810 17530
rect 4900 17290 5140 17530
rect 5230 17290 5470 17530
rect 5560 17290 5800 17530
rect 5890 17290 6130 17530
rect 6220 17290 6460 17530
rect 6550 17290 6790 17530
rect 6880 17290 7120 17530
rect -4670 16960 -4430 17200
rect -4340 16960 -4100 17200
rect -4010 16960 -3770 17200
rect -3680 16960 -3440 17200
rect -3350 16960 -3110 17200
rect -3020 16960 -2780 17200
rect -2690 16960 -2450 17200
rect -2360 16960 -2120 17200
rect -2030 16960 -1790 17200
rect -1700 16960 -1460 17200
rect -1370 16960 -1130 17200
rect -1040 16960 -800 17200
rect -710 16960 -470 17200
rect -380 16960 -140 17200
rect -50 16960 190 17200
rect 280 16960 520 17200
rect 610 16960 850 17200
rect 940 16960 1180 17200
rect 1270 16960 1510 17200
rect 1600 16960 1840 17200
rect 1930 16960 2170 17200
rect 2260 16960 2500 17200
rect 2590 16960 2830 17200
rect 2920 16960 3160 17200
rect 3250 16960 3490 17200
rect 3580 16960 3820 17200
rect 3910 16960 4150 17200
rect 4240 16960 4480 17200
rect 4570 16960 4810 17200
rect 4900 16960 5140 17200
rect 5230 16960 5470 17200
rect 5560 16960 5800 17200
rect 5890 16960 6130 17200
rect 6220 16960 6460 17200
rect 6550 16960 6790 17200
rect 6880 16960 7120 17200
rect -4670 16630 -4430 16870
rect -4340 16630 -4100 16870
rect -4010 16630 -3770 16870
rect -3680 16630 -3440 16870
rect -3350 16630 -3110 16870
rect -3020 16630 -2780 16870
rect -2690 16630 -2450 16870
rect -2360 16630 -2120 16870
rect -2030 16630 -1790 16870
rect -1700 16630 -1460 16870
rect -1370 16630 -1130 16870
rect -1040 16630 -800 16870
rect -710 16630 -470 16870
rect -380 16630 -140 16870
rect -50 16630 190 16870
rect 280 16630 520 16870
rect 610 16630 850 16870
rect 940 16630 1180 16870
rect 1270 16630 1510 16870
rect 1600 16630 1840 16870
rect 1930 16630 2170 16870
rect 2260 16630 2500 16870
rect 2590 16630 2830 16870
rect 2920 16630 3160 16870
rect 3250 16630 3490 16870
rect 3580 16630 3820 16870
rect 3910 16630 4150 16870
rect 4240 16630 4480 16870
rect 4570 16630 4810 16870
rect 4900 16630 5140 16870
rect 5230 16630 5470 16870
rect 5560 16630 5800 16870
rect 5890 16630 6130 16870
rect 6220 16630 6460 16870
rect 6550 16630 6790 16870
rect 6880 16630 7120 16870
rect -4670 16300 -4430 16540
rect -4340 16300 -4100 16540
rect -4010 16300 -3770 16540
rect -3680 16300 -3440 16540
rect -3350 16300 -3110 16540
rect -3020 16300 -2780 16540
rect -2690 16300 -2450 16540
rect -2360 16300 -2120 16540
rect -2030 16300 -1790 16540
rect -1700 16300 -1460 16540
rect -1370 16300 -1130 16540
rect -1040 16300 -800 16540
rect -710 16300 -470 16540
rect -380 16300 -140 16540
rect -50 16300 190 16540
rect 280 16300 520 16540
rect 610 16300 850 16540
rect 940 16300 1180 16540
rect 1270 16300 1510 16540
rect 1600 16300 1840 16540
rect 1930 16300 2170 16540
rect 2260 16300 2500 16540
rect 2590 16300 2830 16540
rect 2920 16300 3160 16540
rect 3250 16300 3490 16540
rect 3580 16300 3820 16540
rect 3910 16300 4150 16540
rect 4240 16300 4480 16540
rect 4570 16300 4810 16540
rect 4900 16300 5140 16540
rect 5230 16300 5470 16540
rect 5560 16300 5800 16540
rect 5890 16300 6130 16540
rect 6220 16300 6460 16540
rect 6550 16300 6790 16540
rect 6880 16300 7120 16540
rect -4670 15970 -4430 16210
rect -4340 15970 -4100 16210
rect -4010 15970 -3770 16210
rect -3680 15970 -3440 16210
rect -3350 15970 -3110 16210
rect -3020 15970 -2780 16210
rect -2690 15970 -2450 16210
rect -2360 15970 -2120 16210
rect -2030 15970 -1790 16210
rect -1700 15970 -1460 16210
rect -1370 15970 -1130 16210
rect -1040 15970 -800 16210
rect -710 15970 -470 16210
rect -380 15970 -140 16210
rect -50 15970 190 16210
rect 280 15970 520 16210
rect 610 15970 850 16210
rect 940 15970 1180 16210
rect 1270 15970 1510 16210
rect 1600 15970 1840 16210
rect 1930 15970 2170 16210
rect 2260 15970 2500 16210
rect 2590 15970 2830 16210
rect 2920 15970 3160 16210
rect 3250 15970 3490 16210
rect 3580 15970 3820 16210
rect 3910 15970 4150 16210
rect 4240 15970 4480 16210
rect 4570 15970 4810 16210
rect 4900 15970 5140 16210
rect 5230 15970 5470 16210
rect 5560 15970 5800 16210
rect 5890 15970 6130 16210
rect 6220 15970 6460 16210
rect 6550 15970 6790 16210
rect 6880 15970 7120 16210
rect -4670 15640 -4430 15880
rect -4340 15640 -4100 15880
rect -4010 15640 -3770 15880
rect -3680 15640 -3440 15880
rect -3350 15640 -3110 15880
rect -3020 15640 -2780 15880
rect -2690 15640 -2450 15880
rect -2360 15640 -2120 15880
rect -2030 15640 -1790 15880
rect -1700 15640 -1460 15880
rect -1370 15640 -1130 15880
rect -1040 15640 -800 15880
rect -710 15640 -470 15880
rect -380 15640 -140 15880
rect -50 15640 190 15880
rect 280 15640 520 15880
rect 610 15640 850 15880
rect 940 15640 1180 15880
rect 1270 15640 1510 15880
rect 1600 15640 1840 15880
rect 1930 15640 2170 15880
rect 2260 15640 2500 15880
rect 2590 15640 2830 15880
rect 2920 15640 3160 15880
rect 3250 15640 3490 15880
rect 3580 15640 3820 15880
rect 3910 15640 4150 15880
rect 4240 15640 4480 15880
rect 4570 15640 4810 15880
rect 4900 15640 5140 15880
rect 5230 15640 5470 15880
rect 5560 15640 5800 15880
rect 5890 15640 6130 15880
rect 6220 15640 6460 15880
rect 6550 15640 6790 15880
rect 6880 15640 7120 15880
rect -4670 15310 -4430 15550
rect -4340 15310 -4100 15550
rect -4010 15310 -3770 15550
rect -3680 15310 -3440 15550
rect -3350 15310 -3110 15550
rect -3020 15310 -2780 15550
rect -2690 15310 -2450 15550
rect -2360 15310 -2120 15550
rect -2030 15310 -1790 15550
rect -1700 15310 -1460 15550
rect -1370 15310 -1130 15550
rect -1040 15310 -800 15550
rect -710 15310 -470 15550
rect -380 15310 -140 15550
rect -50 15310 190 15550
rect 280 15310 520 15550
rect 610 15310 850 15550
rect 940 15310 1180 15550
rect 1270 15310 1510 15550
rect 1600 15310 1840 15550
rect 1930 15310 2170 15550
rect 2260 15310 2500 15550
rect 2590 15310 2830 15550
rect 2920 15310 3160 15550
rect 3250 15310 3490 15550
rect 3580 15310 3820 15550
rect 3910 15310 4150 15550
rect 4240 15310 4480 15550
rect 4570 15310 4810 15550
rect 4900 15310 5140 15550
rect 5230 15310 5470 15550
rect 5560 15310 5800 15550
rect 5890 15310 6130 15550
rect 6220 15310 6460 15550
rect 6550 15310 6790 15550
rect 6880 15310 7120 15550
rect -4670 14980 -4430 15220
rect -4340 14980 -4100 15220
rect -4010 14980 -3770 15220
rect -3680 14980 -3440 15220
rect -3350 14980 -3110 15220
rect -3020 14980 -2780 15220
rect -2690 14980 -2450 15220
rect -2360 14980 -2120 15220
rect -2030 14980 -1790 15220
rect -1700 14980 -1460 15220
rect -1370 14980 -1130 15220
rect -1040 14980 -800 15220
rect -710 14980 -470 15220
rect -380 14980 -140 15220
rect -50 14980 190 15220
rect 280 14980 520 15220
rect 610 14980 850 15220
rect 940 14980 1180 15220
rect 1270 14980 1510 15220
rect 1600 14980 1840 15220
rect 1930 14980 2170 15220
rect 2260 14980 2500 15220
rect 2590 14980 2830 15220
rect 2920 14980 3160 15220
rect 3250 14980 3490 15220
rect 3580 14980 3820 15220
rect 3910 14980 4150 15220
rect 4240 14980 4480 15220
rect 4570 14980 4810 15220
rect 4900 14980 5140 15220
rect 5230 14980 5470 15220
rect 5560 14980 5800 15220
rect 5890 14980 6130 15220
rect 6220 14980 6460 15220
rect 6550 14980 6790 15220
rect 6880 14980 7120 15220
rect -4670 14650 -4430 14890
rect -4340 14650 -4100 14890
rect -4010 14650 -3770 14890
rect -3680 14650 -3440 14890
rect -3350 14650 -3110 14890
rect -3020 14650 -2780 14890
rect -2690 14650 -2450 14890
rect -2360 14650 -2120 14890
rect -2030 14650 -1790 14890
rect -1700 14650 -1460 14890
rect -1370 14650 -1130 14890
rect -1040 14650 -800 14890
rect -710 14650 -470 14890
rect -380 14650 -140 14890
rect -50 14650 190 14890
rect 280 14650 520 14890
rect 610 14650 850 14890
rect 940 14650 1180 14890
rect 1270 14650 1510 14890
rect 1600 14650 1840 14890
rect 1930 14650 2170 14890
rect 2260 14650 2500 14890
rect 2590 14650 2830 14890
rect 2920 14650 3160 14890
rect 3250 14650 3490 14890
rect 3580 14650 3820 14890
rect 3910 14650 4150 14890
rect 4240 14650 4480 14890
rect 4570 14650 4810 14890
rect 4900 14650 5140 14890
rect 5230 14650 5470 14890
rect 5560 14650 5800 14890
rect 5890 14650 6130 14890
rect 6220 14650 6460 14890
rect 6550 14650 6790 14890
rect 6880 14650 7120 14890
rect -4670 14320 -4430 14560
rect -4340 14320 -4100 14560
rect -4010 14320 -3770 14560
rect -3680 14320 -3440 14560
rect -3350 14320 -3110 14560
rect -3020 14320 -2780 14560
rect -2690 14320 -2450 14560
rect -2360 14320 -2120 14560
rect -2030 14320 -1790 14560
rect -1700 14320 -1460 14560
rect -1370 14320 -1130 14560
rect -1040 14320 -800 14560
rect -710 14320 -470 14560
rect -380 14320 -140 14560
rect -50 14320 190 14560
rect 280 14320 520 14560
rect 610 14320 850 14560
rect 940 14320 1180 14560
rect 1270 14320 1510 14560
rect 1600 14320 1840 14560
rect 1930 14320 2170 14560
rect 2260 14320 2500 14560
rect 2590 14320 2830 14560
rect 2920 14320 3160 14560
rect 3250 14320 3490 14560
rect 3580 14320 3820 14560
rect 3910 14320 4150 14560
rect 4240 14320 4480 14560
rect 4570 14320 4810 14560
rect 4900 14320 5140 14560
rect 5230 14320 5470 14560
rect 5560 14320 5800 14560
rect 5890 14320 6130 14560
rect 6220 14320 6460 14560
rect 6550 14320 6790 14560
rect 6880 14320 7120 14560
rect -4670 13990 -4430 14230
rect -4340 13990 -4100 14230
rect -4010 13990 -3770 14230
rect -3680 13990 -3440 14230
rect -3350 13990 -3110 14230
rect -3020 13990 -2780 14230
rect -2690 13990 -2450 14230
rect -2360 13990 -2120 14230
rect -2030 13990 -1790 14230
rect -1700 13990 -1460 14230
rect -1370 13990 -1130 14230
rect -1040 13990 -800 14230
rect -710 13990 -470 14230
rect -380 13990 -140 14230
rect -50 13990 190 14230
rect 280 13990 520 14230
rect 610 13990 850 14230
rect 940 13990 1180 14230
rect 1270 13990 1510 14230
rect 1600 13990 1840 14230
rect 1930 13990 2170 14230
rect 2260 13990 2500 14230
rect 2590 13990 2830 14230
rect 2920 13990 3160 14230
rect 3250 13990 3490 14230
rect 3580 13990 3820 14230
rect 3910 13990 4150 14230
rect 4240 13990 4480 14230
rect 4570 13990 4810 14230
rect 4900 13990 5140 14230
rect 5230 13990 5470 14230
rect 5560 13990 5800 14230
rect 5890 13990 6130 14230
rect 6220 13990 6460 14230
rect 6550 13990 6790 14230
rect 6880 13990 7120 14230
rect -4670 13660 -4430 13900
rect -4340 13660 -4100 13900
rect -4010 13660 -3770 13900
rect -3680 13660 -3440 13900
rect -3350 13660 -3110 13900
rect -3020 13660 -2780 13900
rect -2690 13660 -2450 13900
rect -2360 13660 -2120 13900
rect -2030 13660 -1790 13900
rect -1700 13660 -1460 13900
rect -1370 13660 -1130 13900
rect -1040 13660 -800 13900
rect -710 13660 -470 13900
rect -380 13660 -140 13900
rect -50 13660 190 13900
rect 280 13660 520 13900
rect 610 13660 850 13900
rect 940 13660 1180 13900
rect 1270 13660 1510 13900
rect 1600 13660 1840 13900
rect 1930 13660 2170 13900
rect 2260 13660 2500 13900
rect 2590 13660 2830 13900
rect 2920 13660 3160 13900
rect 3250 13660 3490 13900
rect 3580 13660 3820 13900
rect 3910 13660 4150 13900
rect 4240 13660 4480 13900
rect 4570 13660 4810 13900
rect 4900 13660 5140 13900
rect 5230 13660 5470 13900
rect 5560 13660 5800 13900
rect 5890 13660 6130 13900
rect 6220 13660 6460 13900
rect 6550 13660 6790 13900
rect 6880 13660 7120 13900
rect -4670 13330 -4430 13570
rect -4340 13330 -4100 13570
rect -4010 13330 -3770 13570
rect -3680 13330 -3440 13570
rect -3350 13330 -3110 13570
rect -3020 13330 -2780 13570
rect -2690 13330 -2450 13570
rect -2360 13330 -2120 13570
rect -2030 13330 -1790 13570
rect -1700 13330 -1460 13570
rect -1370 13330 -1130 13570
rect -1040 13330 -800 13570
rect -710 13330 -470 13570
rect -380 13330 -140 13570
rect -50 13330 190 13570
rect 280 13330 520 13570
rect 610 13330 850 13570
rect 940 13330 1180 13570
rect 1270 13330 1510 13570
rect 1600 13330 1840 13570
rect 1930 13330 2170 13570
rect 2260 13330 2500 13570
rect 2590 13330 2830 13570
rect 2920 13330 3160 13570
rect 3250 13330 3490 13570
rect 3580 13330 3820 13570
rect 3910 13330 4150 13570
rect 4240 13330 4480 13570
rect 4570 13330 4810 13570
rect 4900 13330 5140 13570
rect 5230 13330 5470 13570
rect 5560 13330 5800 13570
rect 5890 13330 6130 13570
rect 6220 13330 6460 13570
rect 6550 13330 6790 13570
rect 6880 13330 7120 13570
rect -4670 13000 -4430 13240
rect -4340 13000 -4100 13240
rect -4010 13000 -3770 13240
rect -3680 13000 -3440 13240
rect -3350 13000 -3110 13240
rect -3020 13000 -2780 13240
rect -2690 13000 -2450 13240
rect -2360 13000 -2120 13240
rect -2030 13000 -1790 13240
rect -1700 13000 -1460 13240
rect -1370 13000 -1130 13240
rect -1040 13000 -800 13240
rect -710 13000 -470 13240
rect -380 13000 -140 13240
rect -50 13000 190 13240
rect 280 13000 520 13240
rect 610 13000 850 13240
rect 940 13000 1180 13240
rect 1270 13000 1510 13240
rect 1600 13000 1840 13240
rect 1930 13000 2170 13240
rect 2260 13000 2500 13240
rect 2590 13000 2830 13240
rect 2920 13000 3160 13240
rect 3250 13000 3490 13240
rect 3580 13000 3820 13240
rect 3910 13000 4150 13240
rect 4240 13000 4480 13240
rect 4570 13000 4810 13240
rect 4900 13000 5140 13240
rect 5230 13000 5470 13240
rect 5560 13000 5800 13240
rect 5890 13000 6130 13240
rect 6220 13000 6460 13240
rect 6550 13000 6790 13240
rect 6880 13000 7120 13240
rect -4670 12670 -4430 12910
rect -4340 12670 -4100 12910
rect -4010 12670 -3770 12910
rect -3680 12670 -3440 12910
rect -3350 12670 -3110 12910
rect -3020 12670 -2780 12910
rect -2690 12670 -2450 12910
rect -2360 12670 -2120 12910
rect -2030 12670 -1790 12910
rect -1700 12670 -1460 12910
rect -1370 12670 -1130 12910
rect -1040 12670 -800 12910
rect -710 12670 -470 12910
rect -380 12670 -140 12910
rect -50 12670 190 12910
rect 280 12670 520 12910
rect 610 12670 850 12910
rect 940 12670 1180 12910
rect 1270 12670 1510 12910
rect 1600 12670 1840 12910
rect 1930 12670 2170 12910
rect 2260 12670 2500 12910
rect 2590 12670 2830 12910
rect 2920 12670 3160 12910
rect 3250 12670 3490 12910
rect 3580 12670 3820 12910
rect 3910 12670 4150 12910
rect 4240 12670 4480 12910
rect 4570 12670 4810 12910
rect 4900 12670 5140 12910
rect 5230 12670 5470 12910
rect 5560 12670 5800 12910
rect 5890 12670 6130 12910
rect 6220 12670 6460 12910
rect 6550 12670 6790 12910
rect 6880 12670 7120 12910
rect -4670 12340 -4430 12580
rect -4340 12340 -4100 12580
rect -4010 12340 -3770 12580
rect -3680 12340 -3440 12580
rect -3350 12340 -3110 12580
rect -3020 12340 -2780 12580
rect -2690 12340 -2450 12580
rect -2360 12340 -2120 12580
rect -2030 12340 -1790 12580
rect -1700 12340 -1460 12580
rect -1370 12340 -1130 12580
rect -1040 12340 -800 12580
rect -710 12340 -470 12580
rect -380 12340 -140 12580
rect -50 12340 190 12580
rect 280 12340 520 12580
rect 610 12340 850 12580
rect 940 12340 1180 12580
rect 1270 12340 1510 12580
rect 1600 12340 1840 12580
rect 1930 12340 2170 12580
rect 2260 12340 2500 12580
rect 2590 12340 2830 12580
rect 2920 12340 3160 12580
rect 3250 12340 3490 12580
rect 3580 12340 3820 12580
rect 3910 12340 4150 12580
rect 4240 12340 4480 12580
rect 4570 12340 4810 12580
rect 4900 12340 5140 12580
rect 5230 12340 5470 12580
rect 5560 12340 5800 12580
rect 5890 12340 6130 12580
rect 6220 12340 6460 12580
rect 6550 12340 6790 12580
rect 6880 12340 7120 12580
rect -4670 12010 -4430 12250
rect -4340 12010 -4100 12250
rect -4010 12010 -3770 12250
rect -3680 12010 -3440 12250
rect -3350 12010 -3110 12250
rect -3020 12010 -2780 12250
rect -2690 12010 -2450 12250
rect -2360 12010 -2120 12250
rect -2030 12010 -1790 12250
rect -1700 12010 -1460 12250
rect -1370 12010 -1130 12250
rect -1040 12010 -800 12250
rect -710 12010 -470 12250
rect -380 12010 -140 12250
rect -50 12010 190 12250
rect 280 12010 520 12250
rect 610 12010 850 12250
rect 940 12010 1180 12250
rect 1270 12010 1510 12250
rect 1600 12010 1840 12250
rect 1930 12010 2170 12250
rect 2260 12010 2500 12250
rect 2590 12010 2830 12250
rect 2920 12010 3160 12250
rect 3250 12010 3490 12250
rect 3580 12010 3820 12250
rect 3910 12010 4150 12250
rect 4240 12010 4480 12250
rect 4570 12010 4810 12250
rect 4900 12010 5140 12250
rect 5230 12010 5470 12250
rect 5560 12010 5800 12250
rect 5890 12010 6130 12250
rect 6220 12010 6460 12250
rect 6550 12010 6790 12250
rect 6880 12010 7120 12250
rect -4670 11680 -4430 11920
rect -4340 11680 -4100 11920
rect -4010 11680 -3770 11920
rect -3680 11680 -3440 11920
rect -3350 11680 -3110 11920
rect -3020 11680 -2780 11920
rect -2690 11680 -2450 11920
rect -2360 11680 -2120 11920
rect -2030 11680 -1790 11920
rect -1700 11680 -1460 11920
rect -1370 11680 -1130 11920
rect -1040 11680 -800 11920
rect -710 11680 -470 11920
rect -380 11680 -140 11920
rect -50 11680 190 11920
rect 280 11680 520 11920
rect 610 11680 850 11920
rect 940 11680 1180 11920
rect 1270 11680 1510 11920
rect 1600 11680 1840 11920
rect 1930 11680 2170 11920
rect 2260 11680 2500 11920
rect 2590 11680 2830 11920
rect 2920 11680 3160 11920
rect 3250 11680 3490 11920
rect 3580 11680 3820 11920
rect 3910 11680 4150 11920
rect 4240 11680 4480 11920
rect 4570 11680 4810 11920
rect 4900 11680 5140 11920
rect 5230 11680 5470 11920
rect 5560 11680 5800 11920
rect 5890 11680 6130 11920
rect 6220 11680 6460 11920
rect 6550 11680 6790 11920
rect 6880 11680 7120 11920
rect -4670 11350 -4430 11590
rect -4340 11350 -4100 11590
rect -4010 11350 -3770 11590
rect -3680 11350 -3440 11590
rect -3350 11350 -3110 11590
rect -3020 11350 -2780 11590
rect -2690 11350 -2450 11590
rect -2360 11350 -2120 11590
rect -2030 11350 -1790 11590
rect -1700 11350 -1460 11590
rect -1370 11350 -1130 11590
rect -1040 11350 -800 11590
rect -710 11350 -470 11590
rect -380 11350 -140 11590
rect -50 11350 190 11590
rect 280 11350 520 11590
rect 610 11350 850 11590
rect 940 11350 1180 11590
rect 1270 11350 1510 11590
rect 1600 11350 1840 11590
rect 1930 11350 2170 11590
rect 2260 11350 2500 11590
rect 2590 11350 2830 11590
rect 2920 11350 3160 11590
rect 3250 11350 3490 11590
rect 3580 11350 3820 11590
rect 3910 11350 4150 11590
rect 4240 11350 4480 11590
rect 4570 11350 4810 11590
rect 4900 11350 5140 11590
rect 5230 11350 5470 11590
rect 5560 11350 5800 11590
rect 5890 11350 6130 11590
rect 6220 11350 6460 11590
rect 6550 11350 6790 11590
rect 6880 11350 7120 11590
rect -4670 11020 -4430 11260
rect -4340 11020 -4100 11260
rect -4010 11020 -3770 11260
rect -3680 11020 -3440 11260
rect -3350 11020 -3110 11260
rect -3020 11020 -2780 11260
rect -2690 11020 -2450 11260
rect -2360 11020 -2120 11260
rect -2030 11020 -1790 11260
rect -1700 11020 -1460 11260
rect -1370 11020 -1130 11260
rect -1040 11020 -800 11260
rect -710 11020 -470 11260
rect -380 11020 -140 11260
rect -50 11020 190 11260
rect 280 11020 520 11260
rect 610 11020 850 11260
rect 940 11020 1180 11260
rect 1270 11020 1510 11260
rect 1600 11020 1840 11260
rect 1930 11020 2170 11260
rect 2260 11020 2500 11260
rect 2590 11020 2830 11260
rect 2920 11020 3160 11260
rect 3250 11020 3490 11260
rect 3580 11020 3820 11260
rect 3910 11020 4150 11260
rect 4240 11020 4480 11260
rect 4570 11020 4810 11260
rect 4900 11020 5140 11260
rect 5230 11020 5470 11260
rect 5560 11020 5800 11260
rect 5890 11020 6130 11260
rect 6220 11020 6460 11260
rect 6550 11020 6790 11260
rect 6880 11020 7120 11260
rect -4670 10690 -4430 10930
rect -4340 10690 -4100 10930
rect -4010 10690 -3770 10930
rect -3680 10690 -3440 10930
rect -3350 10690 -3110 10930
rect -3020 10690 -2780 10930
rect -2690 10690 -2450 10930
rect -2360 10690 -2120 10930
rect -2030 10690 -1790 10930
rect -1700 10690 -1460 10930
rect -1370 10690 -1130 10930
rect -1040 10690 -800 10930
rect -710 10690 -470 10930
rect -380 10690 -140 10930
rect -50 10690 190 10930
rect 280 10690 520 10930
rect 610 10690 850 10930
rect 940 10690 1180 10930
rect 1270 10690 1510 10930
rect 1600 10690 1840 10930
rect 1930 10690 2170 10930
rect 2260 10690 2500 10930
rect 2590 10690 2830 10930
rect 2920 10690 3160 10930
rect 3250 10690 3490 10930
rect 3580 10690 3820 10930
rect 3910 10690 4150 10930
rect 4240 10690 4480 10930
rect 4570 10690 4810 10930
rect 4900 10690 5140 10930
rect 5230 10690 5470 10930
rect 5560 10690 5800 10930
rect 5890 10690 6130 10930
rect 6220 10690 6460 10930
rect 6550 10690 6790 10930
rect 6880 10690 7120 10930
rect -4670 10360 -4430 10600
rect -4340 10360 -4100 10600
rect -4010 10360 -3770 10600
rect -3680 10360 -3440 10600
rect -3350 10360 -3110 10600
rect -3020 10360 -2780 10600
rect -2690 10360 -2450 10600
rect -2360 10360 -2120 10600
rect -2030 10360 -1790 10600
rect -1700 10360 -1460 10600
rect -1370 10360 -1130 10600
rect -1040 10360 -800 10600
rect -710 10360 -470 10600
rect -380 10360 -140 10600
rect -50 10360 190 10600
rect 280 10360 520 10600
rect 610 10360 850 10600
rect 940 10360 1180 10600
rect 1270 10360 1510 10600
rect 1600 10360 1840 10600
rect 1930 10360 2170 10600
rect 2260 10360 2500 10600
rect 2590 10360 2830 10600
rect 2920 10360 3160 10600
rect 3250 10360 3490 10600
rect 3580 10360 3820 10600
rect 3910 10360 4150 10600
rect 4240 10360 4480 10600
rect 4570 10360 4810 10600
rect 4900 10360 5140 10600
rect 5230 10360 5470 10600
rect 5560 10360 5800 10600
rect 5890 10360 6130 10600
rect 6220 10360 6460 10600
rect 6550 10360 6790 10600
rect 6880 10360 7120 10600
rect -4670 10030 -4430 10270
rect -4340 10030 -4100 10270
rect -4010 10030 -3770 10270
rect -3680 10030 -3440 10270
rect -3350 10030 -3110 10270
rect -3020 10030 -2780 10270
rect -2690 10030 -2450 10270
rect -2360 10030 -2120 10270
rect -2030 10030 -1790 10270
rect -1700 10030 -1460 10270
rect -1370 10030 -1130 10270
rect -1040 10030 -800 10270
rect -710 10030 -470 10270
rect -380 10030 -140 10270
rect -50 10030 190 10270
rect 280 10030 520 10270
rect 610 10030 850 10270
rect 940 10030 1180 10270
rect 1270 10030 1510 10270
rect 1600 10030 1840 10270
rect 1930 10030 2170 10270
rect 2260 10030 2500 10270
rect 2590 10030 2830 10270
rect 2920 10030 3160 10270
rect 3250 10030 3490 10270
rect 3580 10030 3820 10270
rect 3910 10030 4150 10270
rect 4240 10030 4480 10270
rect 4570 10030 4810 10270
rect 4900 10030 5140 10270
rect 5230 10030 5470 10270
rect 5560 10030 5800 10270
rect 5890 10030 6130 10270
rect 6220 10030 6460 10270
rect 6550 10030 6790 10270
rect 6880 10030 7120 10270
rect -4670 9700 -4430 9940
rect -4340 9700 -4100 9940
rect -4010 9700 -3770 9940
rect -3680 9700 -3440 9940
rect -3350 9700 -3110 9940
rect -3020 9700 -2780 9940
rect -2690 9700 -2450 9940
rect -2360 9700 -2120 9940
rect -2030 9700 -1790 9940
rect -1700 9700 -1460 9940
rect -1370 9700 -1130 9940
rect -1040 9700 -800 9940
rect -710 9700 -470 9940
rect -380 9700 -140 9940
rect -50 9700 190 9940
rect 280 9700 520 9940
rect 610 9700 850 9940
rect 940 9700 1180 9940
rect 1270 9700 1510 9940
rect 1600 9700 1840 9940
rect 1930 9700 2170 9940
rect 2260 9700 2500 9940
rect 2590 9700 2830 9940
rect 2920 9700 3160 9940
rect 3250 9700 3490 9940
rect 3580 9700 3820 9940
rect 3910 9700 4150 9940
rect 4240 9700 4480 9940
rect 4570 9700 4810 9940
rect 4900 9700 5140 9940
rect 5230 9700 5470 9940
rect 5560 9700 5800 9940
rect 5890 9700 6130 9940
rect 6220 9700 6460 9940
rect 6550 9700 6790 9940
rect 6880 9700 7120 9940
rect -4670 9370 -4430 9610
rect -4340 9370 -4100 9610
rect -4010 9370 -3770 9610
rect -3680 9370 -3440 9610
rect -3350 9370 -3110 9610
rect -3020 9370 -2780 9610
rect -2690 9370 -2450 9610
rect -2360 9370 -2120 9610
rect -2030 9370 -1790 9610
rect -1700 9370 -1460 9610
rect -1370 9370 -1130 9610
rect -1040 9370 -800 9610
rect -710 9370 -470 9610
rect -380 9370 -140 9610
rect -50 9370 190 9610
rect 280 9370 520 9610
rect 610 9370 850 9610
rect 940 9370 1180 9610
rect 1270 9370 1510 9610
rect 1600 9370 1840 9610
rect 1930 9370 2170 9610
rect 2260 9370 2500 9610
rect 2590 9370 2830 9610
rect 2920 9370 3160 9610
rect 3250 9370 3490 9610
rect 3580 9370 3820 9610
rect 3910 9370 4150 9610
rect 4240 9370 4480 9610
rect 4570 9370 4810 9610
rect 4900 9370 5140 9610
rect 5230 9370 5470 9610
rect 5560 9370 5800 9610
rect 5890 9370 6130 9610
rect 6220 9370 6460 9610
rect 6550 9370 6790 9610
rect 6880 9370 7120 9610
rect -4670 9040 -4430 9280
rect -4340 9040 -4100 9280
rect -4010 9040 -3770 9280
rect -3680 9040 -3440 9280
rect -3350 9040 -3110 9280
rect -3020 9040 -2780 9280
rect -2690 9040 -2450 9280
rect -2360 9040 -2120 9280
rect -2030 9040 -1790 9280
rect -1700 9040 -1460 9280
rect -1370 9040 -1130 9280
rect -1040 9040 -800 9280
rect -710 9040 -470 9280
rect -380 9040 -140 9280
rect -50 9040 190 9280
rect 280 9040 520 9280
rect 610 9040 850 9280
rect 940 9040 1180 9280
rect 1270 9040 1510 9280
rect 1600 9040 1840 9280
rect 1930 9040 2170 9280
rect 2260 9040 2500 9280
rect 2590 9040 2830 9280
rect 2920 9040 3160 9280
rect 3250 9040 3490 9280
rect 3580 9040 3820 9280
rect 3910 9040 4150 9280
rect 4240 9040 4480 9280
rect 4570 9040 4810 9280
rect 4900 9040 5140 9280
rect 5230 9040 5470 9280
rect 5560 9040 5800 9280
rect 5890 9040 6130 9280
rect 6220 9040 6460 9280
rect 6550 9040 6790 9280
rect 6880 9040 7120 9280
rect 7780 20590 8020 20830
rect 8110 20590 8350 20830
rect 8440 20590 8680 20830
rect 8770 20590 9010 20830
rect 9100 20590 9340 20830
rect 9430 20590 9670 20830
rect 9760 20590 10000 20830
rect 10090 20590 10330 20830
rect 10420 20590 10660 20830
rect 10750 20590 10990 20830
rect 11080 20590 11320 20830
rect 11410 20590 11650 20830
rect 11740 20590 11980 20830
rect 12070 20590 12310 20830
rect 12400 20590 12640 20830
rect 12730 20590 12970 20830
rect 13060 20590 13300 20830
rect 13390 20590 13630 20830
rect 13720 20590 13960 20830
rect 14050 20590 14290 20830
rect 14380 20590 14620 20830
rect 14710 20590 14950 20830
rect 15040 20590 15280 20830
rect 15370 20590 15610 20830
rect 15700 20590 15940 20830
rect 16030 20590 16270 20830
rect 16360 20590 16600 20830
rect 16690 20590 16930 20830
rect 17020 20590 17260 20830
rect 17350 20590 17590 20830
rect 17680 20590 17920 20830
rect 18010 20590 18250 20830
rect 18340 20590 18580 20830
rect 18670 20590 18910 20830
rect 19000 20590 19240 20830
rect 19330 20590 19570 20830
rect 7780 20260 8020 20500
rect 8110 20260 8350 20500
rect 8440 20260 8680 20500
rect 8770 20260 9010 20500
rect 9100 20260 9340 20500
rect 9430 20260 9670 20500
rect 9760 20260 10000 20500
rect 10090 20260 10330 20500
rect 10420 20260 10660 20500
rect 10750 20260 10990 20500
rect 11080 20260 11320 20500
rect 11410 20260 11650 20500
rect 11740 20260 11980 20500
rect 12070 20260 12310 20500
rect 12400 20260 12640 20500
rect 12730 20260 12970 20500
rect 13060 20260 13300 20500
rect 13390 20260 13630 20500
rect 13720 20260 13960 20500
rect 14050 20260 14290 20500
rect 14380 20260 14620 20500
rect 14710 20260 14950 20500
rect 15040 20260 15280 20500
rect 15370 20260 15610 20500
rect 15700 20260 15940 20500
rect 16030 20260 16270 20500
rect 16360 20260 16600 20500
rect 16690 20260 16930 20500
rect 17020 20260 17260 20500
rect 17350 20260 17590 20500
rect 17680 20260 17920 20500
rect 18010 20260 18250 20500
rect 18340 20260 18580 20500
rect 18670 20260 18910 20500
rect 19000 20260 19240 20500
rect 19330 20260 19570 20500
rect 7780 19930 8020 20170
rect 8110 19930 8350 20170
rect 8440 19930 8680 20170
rect 8770 19930 9010 20170
rect 9100 19930 9340 20170
rect 9430 19930 9670 20170
rect 9760 19930 10000 20170
rect 10090 19930 10330 20170
rect 10420 19930 10660 20170
rect 10750 19930 10990 20170
rect 11080 19930 11320 20170
rect 11410 19930 11650 20170
rect 11740 19930 11980 20170
rect 12070 19930 12310 20170
rect 12400 19930 12640 20170
rect 12730 19930 12970 20170
rect 13060 19930 13300 20170
rect 13390 19930 13630 20170
rect 13720 19930 13960 20170
rect 14050 19930 14290 20170
rect 14380 19930 14620 20170
rect 14710 19930 14950 20170
rect 15040 19930 15280 20170
rect 15370 19930 15610 20170
rect 15700 19930 15940 20170
rect 16030 19930 16270 20170
rect 16360 19930 16600 20170
rect 16690 19930 16930 20170
rect 17020 19930 17260 20170
rect 17350 19930 17590 20170
rect 17680 19930 17920 20170
rect 18010 19930 18250 20170
rect 18340 19930 18580 20170
rect 18670 19930 18910 20170
rect 19000 19930 19240 20170
rect 19330 19930 19570 20170
rect 7780 19600 8020 19840
rect 8110 19600 8350 19840
rect 8440 19600 8680 19840
rect 8770 19600 9010 19840
rect 9100 19600 9340 19840
rect 9430 19600 9670 19840
rect 9760 19600 10000 19840
rect 10090 19600 10330 19840
rect 10420 19600 10660 19840
rect 10750 19600 10990 19840
rect 11080 19600 11320 19840
rect 11410 19600 11650 19840
rect 11740 19600 11980 19840
rect 12070 19600 12310 19840
rect 12400 19600 12640 19840
rect 12730 19600 12970 19840
rect 13060 19600 13300 19840
rect 13390 19600 13630 19840
rect 13720 19600 13960 19840
rect 14050 19600 14290 19840
rect 14380 19600 14620 19840
rect 14710 19600 14950 19840
rect 15040 19600 15280 19840
rect 15370 19600 15610 19840
rect 15700 19600 15940 19840
rect 16030 19600 16270 19840
rect 16360 19600 16600 19840
rect 16690 19600 16930 19840
rect 17020 19600 17260 19840
rect 17350 19600 17590 19840
rect 17680 19600 17920 19840
rect 18010 19600 18250 19840
rect 18340 19600 18580 19840
rect 18670 19600 18910 19840
rect 19000 19600 19240 19840
rect 19330 19600 19570 19840
rect 7780 19270 8020 19510
rect 8110 19270 8350 19510
rect 8440 19270 8680 19510
rect 8770 19270 9010 19510
rect 9100 19270 9340 19510
rect 9430 19270 9670 19510
rect 9760 19270 10000 19510
rect 10090 19270 10330 19510
rect 10420 19270 10660 19510
rect 10750 19270 10990 19510
rect 11080 19270 11320 19510
rect 11410 19270 11650 19510
rect 11740 19270 11980 19510
rect 12070 19270 12310 19510
rect 12400 19270 12640 19510
rect 12730 19270 12970 19510
rect 13060 19270 13300 19510
rect 13390 19270 13630 19510
rect 13720 19270 13960 19510
rect 14050 19270 14290 19510
rect 14380 19270 14620 19510
rect 14710 19270 14950 19510
rect 15040 19270 15280 19510
rect 15370 19270 15610 19510
rect 15700 19270 15940 19510
rect 16030 19270 16270 19510
rect 16360 19270 16600 19510
rect 16690 19270 16930 19510
rect 17020 19270 17260 19510
rect 17350 19270 17590 19510
rect 17680 19270 17920 19510
rect 18010 19270 18250 19510
rect 18340 19270 18580 19510
rect 18670 19270 18910 19510
rect 19000 19270 19240 19510
rect 19330 19270 19570 19510
rect 7780 18940 8020 19180
rect 8110 18940 8350 19180
rect 8440 18940 8680 19180
rect 8770 18940 9010 19180
rect 9100 18940 9340 19180
rect 9430 18940 9670 19180
rect 9760 18940 10000 19180
rect 10090 18940 10330 19180
rect 10420 18940 10660 19180
rect 10750 18940 10990 19180
rect 11080 18940 11320 19180
rect 11410 18940 11650 19180
rect 11740 18940 11980 19180
rect 12070 18940 12310 19180
rect 12400 18940 12640 19180
rect 12730 18940 12970 19180
rect 13060 18940 13300 19180
rect 13390 18940 13630 19180
rect 13720 18940 13960 19180
rect 14050 18940 14290 19180
rect 14380 18940 14620 19180
rect 14710 18940 14950 19180
rect 15040 18940 15280 19180
rect 15370 18940 15610 19180
rect 15700 18940 15940 19180
rect 16030 18940 16270 19180
rect 16360 18940 16600 19180
rect 16690 18940 16930 19180
rect 17020 18940 17260 19180
rect 17350 18940 17590 19180
rect 17680 18940 17920 19180
rect 18010 18940 18250 19180
rect 18340 18940 18580 19180
rect 18670 18940 18910 19180
rect 19000 18940 19240 19180
rect 19330 18940 19570 19180
rect 7780 18610 8020 18850
rect 8110 18610 8350 18850
rect 8440 18610 8680 18850
rect 8770 18610 9010 18850
rect 9100 18610 9340 18850
rect 9430 18610 9670 18850
rect 9760 18610 10000 18850
rect 10090 18610 10330 18850
rect 10420 18610 10660 18850
rect 10750 18610 10990 18850
rect 11080 18610 11320 18850
rect 11410 18610 11650 18850
rect 11740 18610 11980 18850
rect 12070 18610 12310 18850
rect 12400 18610 12640 18850
rect 12730 18610 12970 18850
rect 13060 18610 13300 18850
rect 13390 18610 13630 18850
rect 13720 18610 13960 18850
rect 14050 18610 14290 18850
rect 14380 18610 14620 18850
rect 14710 18610 14950 18850
rect 15040 18610 15280 18850
rect 15370 18610 15610 18850
rect 15700 18610 15940 18850
rect 16030 18610 16270 18850
rect 16360 18610 16600 18850
rect 16690 18610 16930 18850
rect 17020 18610 17260 18850
rect 17350 18610 17590 18850
rect 17680 18610 17920 18850
rect 18010 18610 18250 18850
rect 18340 18610 18580 18850
rect 18670 18610 18910 18850
rect 19000 18610 19240 18850
rect 19330 18610 19570 18850
rect 7780 18280 8020 18520
rect 8110 18280 8350 18520
rect 8440 18280 8680 18520
rect 8770 18280 9010 18520
rect 9100 18280 9340 18520
rect 9430 18280 9670 18520
rect 9760 18280 10000 18520
rect 10090 18280 10330 18520
rect 10420 18280 10660 18520
rect 10750 18280 10990 18520
rect 11080 18280 11320 18520
rect 11410 18280 11650 18520
rect 11740 18280 11980 18520
rect 12070 18280 12310 18520
rect 12400 18280 12640 18520
rect 12730 18280 12970 18520
rect 13060 18280 13300 18520
rect 13390 18280 13630 18520
rect 13720 18280 13960 18520
rect 14050 18280 14290 18520
rect 14380 18280 14620 18520
rect 14710 18280 14950 18520
rect 15040 18280 15280 18520
rect 15370 18280 15610 18520
rect 15700 18280 15940 18520
rect 16030 18280 16270 18520
rect 16360 18280 16600 18520
rect 16690 18280 16930 18520
rect 17020 18280 17260 18520
rect 17350 18280 17590 18520
rect 17680 18280 17920 18520
rect 18010 18280 18250 18520
rect 18340 18280 18580 18520
rect 18670 18280 18910 18520
rect 19000 18280 19240 18520
rect 19330 18280 19570 18520
rect 7780 17950 8020 18190
rect 8110 17950 8350 18190
rect 8440 17950 8680 18190
rect 8770 17950 9010 18190
rect 9100 17950 9340 18190
rect 9430 17950 9670 18190
rect 9760 17950 10000 18190
rect 10090 17950 10330 18190
rect 10420 17950 10660 18190
rect 10750 17950 10990 18190
rect 11080 17950 11320 18190
rect 11410 17950 11650 18190
rect 11740 17950 11980 18190
rect 12070 17950 12310 18190
rect 12400 17950 12640 18190
rect 12730 17950 12970 18190
rect 13060 17950 13300 18190
rect 13390 17950 13630 18190
rect 13720 17950 13960 18190
rect 14050 17950 14290 18190
rect 14380 17950 14620 18190
rect 14710 17950 14950 18190
rect 15040 17950 15280 18190
rect 15370 17950 15610 18190
rect 15700 17950 15940 18190
rect 16030 17950 16270 18190
rect 16360 17950 16600 18190
rect 16690 17950 16930 18190
rect 17020 17950 17260 18190
rect 17350 17950 17590 18190
rect 17680 17950 17920 18190
rect 18010 17950 18250 18190
rect 18340 17950 18580 18190
rect 18670 17950 18910 18190
rect 19000 17950 19240 18190
rect 19330 17950 19570 18190
rect 7780 17620 8020 17860
rect 8110 17620 8350 17860
rect 8440 17620 8680 17860
rect 8770 17620 9010 17860
rect 9100 17620 9340 17860
rect 9430 17620 9670 17860
rect 9760 17620 10000 17860
rect 10090 17620 10330 17860
rect 10420 17620 10660 17860
rect 10750 17620 10990 17860
rect 11080 17620 11320 17860
rect 11410 17620 11650 17860
rect 11740 17620 11980 17860
rect 12070 17620 12310 17860
rect 12400 17620 12640 17860
rect 12730 17620 12970 17860
rect 13060 17620 13300 17860
rect 13390 17620 13630 17860
rect 13720 17620 13960 17860
rect 14050 17620 14290 17860
rect 14380 17620 14620 17860
rect 14710 17620 14950 17860
rect 15040 17620 15280 17860
rect 15370 17620 15610 17860
rect 15700 17620 15940 17860
rect 16030 17620 16270 17860
rect 16360 17620 16600 17860
rect 16690 17620 16930 17860
rect 17020 17620 17260 17860
rect 17350 17620 17590 17860
rect 17680 17620 17920 17860
rect 18010 17620 18250 17860
rect 18340 17620 18580 17860
rect 18670 17620 18910 17860
rect 19000 17620 19240 17860
rect 19330 17620 19570 17860
rect 7780 17290 8020 17530
rect 8110 17290 8350 17530
rect 8440 17290 8680 17530
rect 8770 17290 9010 17530
rect 9100 17290 9340 17530
rect 9430 17290 9670 17530
rect 9760 17290 10000 17530
rect 10090 17290 10330 17530
rect 10420 17290 10660 17530
rect 10750 17290 10990 17530
rect 11080 17290 11320 17530
rect 11410 17290 11650 17530
rect 11740 17290 11980 17530
rect 12070 17290 12310 17530
rect 12400 17290 12640 17530
rect 12730 17290 12970 17530
rect 13060 17290 13300 17530
rect 13390 17290 13630 17530
rect 13720 17290 13960 17530
rect 14050 17290 14290 17530
rect 14380 17290 14620 17530
rect 14710 17290 14950 17530
rect 15040 17290 15280 17530
rect 15370 17290 15610 17530
rect 15700 17290 15940 17530
rect 16030 17290 16270 17530
rect 16360 17290 16600 17530
rect 16690 17290 16930 17530
rect 17020 17290 17260 17530
rect 17350 17290 17590 17530
rect 17680 17290 17920 17530
rect 18010 17290 18250 17530
rect 18340 17290 18580 17530
rect 18670 17290 18910 17530
rect 19000 17290 19240 17530
rect 19330 17290 19570 17530
rect 7780 16960 8020 17200
rect 8110 16960 8350 17200
rect 8440 16960 8680 17200
rect 8770 16960 9010 17200
rect 9100 16960 9340 17200
rect 9430 16960 9670 17200
rect 9760 16960 10000 17200
rect 10090 16960 10330 17200
rect 10420 16960 10660 17200
rect 10750 16960 10990 17200
rect 11080 16960 11320 17200
rect 11410 16960 11650 17200
rect 11740 16960 11980 17200
rect 12070 16960 12310 17200
rect 12400 16960 12640 17200
rect 12730 16960 12970 17200
rect 13060 16960 13300 17200
rect 13390 16960 13630 17200
rect 13720 16960 13960 17200
rect 14050 16960 14290 17200
rect 14380 16960 14620 17200
rect 14710 16960 14950 17200
rect 15040 16960 15280 17200
rect 15370 16960 15610 17200
rect 15700 16960 15940 17200
rect 16030 16960 16270 17200
rect 16360 16960 16600 17200
rect 16690 16960 16930 17200
rect 17020 16960 17260 17200
rect 17350 16960 17590 17200
rect 17680 16960 17920 17200
rect 18010 16960 18250 17200
rect 18340 16960 18580 17200
rect 18670 16960 18910 17200
rect 19000 16960 19240 17200
rect 19330 16960 19570 17200
rect 7780 16630 8020 16870
rect 8110 16630 8350 16870
rect 8440 16630 8680 16870
rect 8770 16630 9010 16870
rect 9100 16630 9340 16870
rect 9430 16630 9670 16870
rect 9760 16630 10000 16870
rect 10090 16630 10330 16870
rect 10420 16630 10660 16870
rect 10750 16630 10990 16870
rect 11080 16630 11320 16870
rect 11410 16630 11650 16870
rect 11740 16630 11980 16870
rect 12070 16630 12310 16870
rect 12400 16630 12640 16870
rect 12730 16630 12970 16870
rect 13060 16630 13300 16870
rect 13390 16630 13630 16870
rect 13720 16630 13960 16870
rect 14050 16630 14290 16870
rect 14380 16630 14620 16870
rect 14710 16630 14950 16870
rect 15040 16630 15280 16870
rect 15370 16630 15610 16870
rect 15700 16630 15940 16870
rect 16030 16630 16270 16870
rect 16360 16630 16600 16870
rect 16690 16630 16930 16870
rect 17020 16630 17260 16870
rect 17350 16630 17590 16870
rect 17680 16630 17920 16870
rect 18010 16630 18250 16870
rect 18340 16630 18580 16870
rect 18670 16630 18910 16870
rect 19000 16630 19240 16870
rect 19330 16630 19570 16870
rect 7780 16300 8020 16540
rect 8110 16300 8350 16540
rect 8440 16300 8680 16540
rect 8770 16300 9010 16540
rect 9100 16300 9340 16540
rect 9430 16300 9670 16540
rect 9760 16300 10000 16540
rect 10090 16300 10330 16540
rect 10420 16300 10660 16540
rect 10750 16300 10990 16540
rect 11080 16300 11320 16540
rect 11410 16300 11650 16540
rect 11740 16300 11980 16540
rect 12070 16300 12310 16540
rect 12400 16300 12640 16540
rect 12730 16300 12970 16540
rect 13060 16300 13300 16540
rect 13390 16300 13630 16540
rect 13720 16300 13960 16540
rect 14050 16300 14290 16540
rect 14380 16300 14620 16540
rect 14710 16300 14950 16540
rect 15040 16300 15280 16540
rect 15370 16300 15610 16540
rect 15700 16300 15940 16540
rect 16030 16300 16270 16540
rect 16360 16300 16600 16540
rect 16690 16300 16930 16540
rect 17020 16300 17260 16540
rect 17350 16300 17590 16540
rect 17680 16300 17920 16540
rect 18010 16300 18250 16540
rect 18340 16300 18580 16540
rect 18670 16300 18910 16540
rect 19000 16300 19240 16540
rect 19330 16300 19570 16540
rect 7780 15970 8020 16210
rect 8110 15970 8350 16210
rect 8440 15970 8680 16210
rect 8770 15970 9010 16210
rect 9100 15970 9340 16210
rect 9430 15970 9670 16210
rect 9760 15970 10000 16210
rect 10090 15970 10330 16210
rect 10420 15970 10660 16210
rect 10750 15970 10990 16210
rect 11080 15970 11320 16210
rect 11410 15970 11650 16210
rect 11740 15970 11980 16210
rect 12070 15970 12310 16210
rect 12400 15970 12640 16210
rect 12730 15970 12970 16210
rect 13060 15970 13300 16210
rect 13390 15970 13630 16210
rect 13720 15970 13960 16210
rect 14050 15970 14290 16210
rect 14380 15970 14620 16210
rect 14710 15970 14950 16210
rect 15040 15970 15280 16210
rect 15370 15970 15610 16210
rect 15700 15970 15940 16210
rect 16030 15970 16270 16210
rect 16360 15970 16600 16210
rect 16690 15970 16930 16210
rect 17020 15970 17260 16210
rect 17350 15970 17590 16210
rect 17680 15970 17920 16210
rect 18010 15970 18250 16210
rect 18340 15970 18580 16210
rect 18670 15970 18910 16210
rect 19000 15970 19240 16210
rect 19330 15970 19570 16210
rect 7780 15640 8020 15880
rect 8110 15640 8350 15880
rect 8440 15640 8680 15880
rect 8770 15640 9010 15880
rect 9100 15640 9340 15880
rect 9430 15640 9670 15880
rect 9760 15640 10000 15880
rect 10090 15640 10330 15880
rect 10420 15640 10660 15880
rect 10750 15640 10990 15880
rect 11080 15640 11320 15880
rect 11410 15640 11650 15880
rect 11740 15640 11980 15880
rect 12070 15640 12310 15880
rect 12400 15640 12640 15880
rect 12730 15640 12970 15880
rect 13060 15640 13300 15880
rect 13390 15640 13630 15880
rect 13720 15640 13960 15880
rect 14050 15640 14290 15880
rect 14380 15640 14620 15880
rect 14710 15640 14950 15880
rect 15040 15640 15280 15880
rect 15370 15640 15610 15880
rect 15700 15640 15940 15880
rect 16030 15640 16270 15880
rect 16360 15640 16600 15880
rect 16690 15640 16930 15880
rect 17020 15640 17260 15880
rect 17350 15640 17590 15880
rect 17680 15640 17920 15880
rect 18010 15640 18250 15880
rect 18340 15640 18580 15880
rect 18670 15640 18910 15880
rect 19000 15640 19240 15880
rect 19330 15640 19570 15880
rect 7780 15310 8020 15550
rect 8110 15310 8350 15550
rect 8440 15310 8680 15550
rect 8770 15310 9010 15550
rect 9100 15310 9340 15550
rect 9430 15310 9670 15550
rect 9760 15310 10000 15550
rect 10090 15310 10330 15550
rect 10420 15310 10660 15550
rect 10750 15310 10990 15550
rect 11080 15310 11320 15550
rect 11410 15310 11650 15550
rect 11740 15310 11980 15550
rect 12070 15310 12310 15550
rect 12400 15310 12640 15550
rect 12730 15310 12970 15550
rect 13060 15310 13300 15550
rect 13390 15310 13630 15550
rect 13720 15310 13960 15550
rect 14050 15310 14290 15550
rect 14380 15310 14620 15550
rect 14710 15310 14950 15550
rect 15040 15310 15280 15550
rect 15370 15310 15610 15550
rect 15700 15310 15940 15550
rect 16030 15310 16270 15550
rect 16360 15310 16600 15550
rect 16690 15310 16930 15550
rect 17020 15310 17260 15550
rect 17350 15310 17590 15550
rect 17680 15310 17920 15550
rect 18010 15310 18250 15550
rect 18340 15310 18580 15550
rect 18670 15310 18910 15550
rect 19000 15310 19240 15550
rect 19330 15310 19570 15550
rect 7780 14980 8020 15220
rect 8110 14980 8350 15220
rect 8440 14980 8680 15220
rect 8770 14980 9010 15220
rect 9100 14980 9340 15220
rect 9430 14980 9670 15220
rect 9760 14980 10000 15220
rect 10090 14980 10330 15220
rect 10420 14980 10660 15220
rect 10750 14980 10990 15220
rect 11080 14980 11320 15220
rect 11410 14980 11650 15220
rect 11740 14980 11980 15220
rect 12070 14980 12310 15220
rect 12400 14980 12640 15220
rect 12730 14980 12970 15220
rect 13060 14980 13300 15220
rect 13390 14980 13630 15220
rect 13720 14980 13960 15220
rect 14050 14980 14290 15220
rect 14380 14980 14620 15220
rect 14710 14980 14950 15220
rect 15040 14980 15280 15220
rect 15370 14980 15610 15220
rect 15700 14980 15940 15220
rect 16030 14980 16270 15220
rect 16360 14980 16600 15220
rect 16690 14980 16930 15220
rect 17020 14980 17260 15220
rect 17350 14980 17590 15220
rect 17680 14980 17920 15220
rect 18010 14980 18250 15220
rect 18340 14980 18580 15220
rect 18670 14980 18910 15220
rect 19000 14980 19240 15220
rect 19330 14980 19570 15220
rect 7780 14650 8020 14890
rect 8110 14650 8350 14890
rect 8440 14650 8680 14890
rect 8770 14650 9010 14890
rect 9100 14650 9340 14890
rect 9430 14650 9670 14890
rect 9760 14650 10000 14890
rect 10090 14650 10330 14890
rect 10420 14650 10660 14890
rect 10750 14650 10990 14890
rect 11080 14650 11320 14890
rect 11410 14650 11650 14890
rect 11740 14650 11980 14890
rect 12070 14650 12310 14890
rect 12400 14650 12640 14890
rect 12730 14650 12970 14890
rect 13060 14650 13300 14890
rect 13390 14650 13630 14890
rect 13720 14650 13960 14890
rect 14050 14650 14290 14890
rect 14380 14650 14620 14890
rect 14710 14650 14950 14890
rect 15040 14650 15280 14890
rect 15370 14650 15610 14890
rect 15700 14650 15940 14890
rect 16030 14650 16270 14890
rect 16360 14650 16600 14890
rect 16690 14650 16930 14890
rect 17020 14650 17260 14890
rect 17350 14650 17590 14890
rect 17680 14650 17920 14890
rect 18010 14650 18250 14890
rect 18340 14650 18580 14890
rect 18670 14650 18910 14890
rect 19000 14650 19240 14890
rect 19330 14650 19570 14890
rect 7780 14320 8020 14560
rect 8110 14320 8350 14560
rect 8440 14320 8680 14560
rect 8770 14320 9010 14560
rect 9100 14320 9340 14560
rect 9430 14320 9670 14560
rect 9760 14320 10000 14560
rect 10090 14320 10330 14560
rect 10420 14320 10660 14560
rect 10750 14320 10990 14560
rect 11080 14320 11320 14560
rect 11410 14320 11650 14560
rect 11740 14320 11980 14560
rect 12070 14320 12310 14560
rect 12400 14320 12640 14560
rect 12730 14320 12970 14560
rect 13060 14320 13300 14560
rect 13390 14320 13630 14560
rect 13720 14320 13960 14560
rect 14050 14320 14290 14560
rect 14380 14320 14620 14560
rect 14710 14320 14950 14560
rect 15040 14320 15280 14560
rect 15370 14320 15610 14560
rect 15700 14320 15940 14560
rect 16030 14320 16270 14560
rect 16360 14320 16600 14560
rect 16690 14320 16930 14560
rect 17020 14320 17260 14560
rect 17350 14320 17590 14560
rect 17680 14320 17920 14560
rect 18010 14320 18250 14560
rect 18340 14320 18580 14560
rect 18670 14320 18910 14560
rect 19000 14320 19240 14560
rect 19330 14320 19570 14560
rect 7780 13990 8020 14230
rect 8110 13990 8350 14230
rect 8440 13990 8680 14230
rect 8770 13990 9010 14230
rect 9100 13990 9340 14230
rect 9430 13990 9670 14230
rect 9760 13990 10000 14230
rect 10090 13990 10330 14230
rect 10420 13990 10660 14230
rect 10750 13990 10990 14230
rect 11080 13990 11320 14230
rect 11410 13990 11650 14230
rect 11740 13990 11980 14230
rect 12070 13990 12310 14230
rect 12400 13990 12640 14230
rect 12730 13990 12970 14230
rect 13060 13990 13300 14230
rect 13390 13990 13630 14230
rect 13720 13990 13960 14230
rect 14050 13990 14290 14230
rect 14380 13990 14620 14230
rect 14710 13990 14950 14230
rect 15040 13990 15280 14230
rect 15370 13990 15610 14230
rect 15700 13990 15940 14230
rect 16030 13990 16270 14230
rect 16360 13990 16600 14230
rect 16690 13990 16930 14230
rect 17020 13990 17260 14230
rect 17350 13990 17590 14230
rect 17680 13990 17920 14230
rect 18010 13990 18250 14230
rect 18340 13990 18580 14230
rect 18670 13990 18910 14230
rect 19000 13990 19240 14230
rect 19330 13990 19570 14230
rect 7780 13660 8020 13900
rect 8110 13660 8350 13900
rect 8440 13660 8680 13900
rect 8770 13660 9010 13900
rect 9100 13660 9340 13900
rect 9430 13660 9670 13900
rect 9760 13660 10000 13900
rect 10090 13660 10330 13900
rect 10420 13660 10660 13900
rect 10750 13660 10990 13900
rect 11080 13660 11320 13900
rect 11410 13660 11650 13900
rect 11740 13660 11980 13900
rect 12070 13660 12310 13900
rect 12400 13660 12640 13900
rect 12730 13660 12970 13900
rect 13060 13660 13300 13900
rect 13390 13660 13630 13900
rect 13720 13660 13960 13900
rect 14050 13660 14290 13900
rect 14380 13660 14620 13900
rect 14710 13660 14950 13900
rect 15040 13660 15280 13900
rect 15370 13660 15610 13900
rect 15700 13660 15940 13900
rect 16030 13660 16270 13900
rect 16360 13660 16600 13900
rect 16690 13660 16930 13900
rect 17020 13660 17260 13900
rect 17350 13660 17590 13900
rect 17680 13660 17920 13900
rect 18010 13660 18250 13900
rect 18340 13660 18580 13900
rect 18670 13660 18910 13900
rect 19000 13660 19240 13900
rect 19330 13660 19570 13900
rect 7780 13330 8020 13570
rect 8110 13330 8350 13570
rect 8440 13330 8680 13570
rect 8770 13330 9010 13570
rect 9100 13330 9340 13570
rect 9430 13330 9670 13570
rect 9760 13330 10000 13570
rect 10090 13330 10330 13570
rect 10420 13330 10660 13570
rect 10750 13330 10990 13570
rect 11080 13330 11320 13570
rect 11410 13330 11650 13570
rect 11740 13330 11980 13570
rect 12070 13330 12310 13570
rect 12400 13330 12640 13570
rect 12730 13330 12970 13570
rect 13060 13330 13300 13570
rect 13390 13330 13630 13570
rect 13720 13330 13960 13570
rect 14050 13330 14290 13570
rect 14380 13330 14620 13570
rect 14710 13330 14950 13570
rect 15040 13330 15280 13570
rect 15370 13330 15610 13570
rect 15700 13330 15940 13570
rect 16030 13330 16270 13570
rect 16360 13330 16600 13570
rect 16690 13330 16930 13570
rect 17020 13330 17260 13570
rect 17350 13330 17590 13570
rect 17680 13330 17920 13570
rect 18010 13330 18250 13570
rect 18340 13330 18580 13570
rect 18670 13330 18910 13570
rect 19000 13330 19240 13570
rect 19330 13330 19570 13570
rect 7780 13000 8020 13240
rect 8110 13000 8350 13240
rect 8440 13000 8680 13240
rect 8770 13000 9010 13240
rect 9100 13000 9340 13240
rect 9430 13000 9670 13240
rect 9760 13000 10000 13240
rect 10090 13000 10330 13240
rect 10420 13000 10660 13240
rect 10750 13000 10990 13240
rect 11080 13000 11320 13240
rect 11410 13000 11650 13240
rect 11740 13000 11980 13240
rect 12070 13000 12310 13240
rect 12400 13000 12640 13240
rect 12730 13000 12970 13240
rect 13060 13000 13300 13240
rect 13390 13000 13630 13240
rect 13720 13000 13960 13240
rect 14050 13000 14290 13240
rect 14380 13000 14620 13240
rect 14710 13000 14950 13240
rect 15040 13000 15280 13240
rect 15370 13000 15610 13240
rect 15700 13000 15940 13240
rect 16030 13000 16270 13240
rect 16360 13000 16600 13240
rect 16690 13000 16930 13240
rect 17020 13000 17260 13240
rect 17350 13000 17590 13240
rect 17680 13000 17920 13240
rect 18010 13000 18250 13240
rect 18340 13000 18580 13240
rect 18670 13000 18910 13240
rect 19000 13000 19240 13240
rect 19330 13000 19570 13240
rect 7780 12670 8020 12910
rect 8110 12670 8350 12910
rect 8440 12670 8680 12910
rect 8770 12670 9010 12910
rect 9100 12670 9340 12910
rect 9430 12670 9670 12910
rect 9760 12670 10000 12910
rect 10090 12670 10330 12910
rect 10420 12670 10660 12910
rect 10750 12670 10990 12910
rect 11080 12670 11320 12910
rect 11410 12670 11650 12910
rect 11740 12670 11980 12910
rect 12070 12670 12310 12910
rect 12400 12670 12640 12910
rect 12730 12670 12970 12910
rect 13060 12670 13300 12910
rect 13390 12670 13630 12910
rect 13720 12670 13960 12910
rect 14050 12670 14290 12910
rect 14380 12670 14620 12910
rect 14710 12670 14950 12910
rect 15040 12670 15280 12910
rect 15370 12670 15610 12910
rect 15700 12670 15940 12910
rect 16030 12670 16270 12910
rect 16360 12670 16600 12910
rect 16690 12670 16930 12910
rect 17020 12670 17260 12910
rect 17350 12670 17590 12910
rect 17680 12670 17920 12910
rect 18010 12670 18250 12910
rect 18340 12670 18580 12910
rect 18670 12670 18910 12910
rect 19000 12670 19240 12910
rect 19330 12670 19570 12910
rect 7780 12340 8020 12580
rect 8110 12340 8350 12580
rect 8440 12340 8680 12580
rect 8770 12340 9010 12580
rect 9100 12340 9340 12580
rect 9430 12340 9670 12580
rect 9760 12340 10000 12580
rect 10090 12340 10330 12580
rect 10420 12340 10660 12580
rect 10750 12340 10990 12580
rect 11080 12340 11320 12580
rect 11410 12340 11650 12580
rect 11740 12340 11980 12580
rect 12070 12340 12310 12580
rect 12400 12340 12640 12580
rect 12730 12340 12970 12580
rect 13060 12340 13300 12580
rect 13390 12340 13630 12580
rect 13720 12340 13960 12580
rect 14050 12340 14290 12580
rect 14380 12340 14620 12580
rect 14710 12340 14950 12580
rect 15040 12340 15280 12580
rect 15370 12340 15610 12580
rect 15700 12340 15940 12580
rect 16030 12340 16270 12580
rect 16360 12340 16600 12580
rect 16690 12340 16930 12580
rect 17020 12340 17260 12580
rect 17350 12340 17590 12580
rect 17680 12340 17920 12580
rect 18010 12340 18250 12580
rect 18340 12340 18580 12580
rect 18670 12340 18910 12580
rect 19000 12340 19240 12580
rect 19330 12340 19570 12580
rect 7780 12010 8020 12250
rect 8110 12010 8350 12250
rect 8440 12010 8680 12250
rect 8770 12010 9010 12250
rect 9100 12010 9340 12250
rect 9430 12010 9670 12250
rect 9760 12010 10000 12250
rect 10090 12010 10330 12250
rect 10420 12010 10660 12250
rect 10750 12010 10990 12250
rect 11080 12010 11320 12250
rect 11410 12010 11650 12250
rect 11740 12010 11980 12250
rect 12070 12010 12310 12250
rect 12400 12010 12640 12250
rect 12730 12010 12970 12250
rect 13060 12010 13300 12250
rect 13390 12010 13630 12250
rect 13720 12010 13960 12250
rect 14050 12010 14290 12250
rect 14380 12010 14620 12250
rect 14710 12010 14950 12250
rect 15040 12010 15280 12250
rect 15370 12010 15610 12250
rect 15700 12010 15940 12250
rect 16030 12010 16270 12250
rect 16360 12010 16600 12250
rect 16690 12010 16930 12250
rect 17020 12010 17260 12250
rect 17350 12010 17590 12250
rect 17680 12010 17920 12250
rect 18010 12010 18250 12250
rect 18340 12010 18580 12250
rect 18670 12010 18910 12250
rect 19000 12010 19240 12250
rect 19330 12010 19570 12250
rect 7780 11680 8020 11920
rect 8110 11680 8350 11920
rect 8440 11680 8680 11920
rect 8770 11680 9010 11920
rect 9100 11680 9340 11920
rect 9430 11680 9670 11920
rect 9760 11680 10000 11920
rect 10090 11680 10330 11920
rect 10420 11680 10660 11920
rect 10750 11680 10990 11920
rect 11080 11680 11320 11920
rect 11410 11680 11650 11920
rect 11740 11680 11980 11920
rect 12070 11680 12310 11920
rect 12400 11680 12640 11920
rect 12730 11680 12970 11920
rect 13060 11680 13300 11920
rect 13390 11680 13630 11920
rect 13720 11680 13960 11920
rect 14050 11680 14290 11920
rect 14380 11680 14620 11920
rect 14710 11680 14950 11920
rect 15040 11680 15280 11920
rect 15370 11680 15610 11920
rect 15700 11680 15940 11920
rect 16030 11680 16270 11920
rect 16360 11680 16600 11920
rect 16690 11680 16930 11920
rect 17020 11680 17260 11920
rect 17350 11680 17590 11920
rect 17680 11680 17920 11920
rect 18010 11680 18250 11920
rect 18340 11680 18580 11920
rect 18670 11680 18910 11920
rect 19000 11680 19240 11920
rect 19330 11680 19570 11920
rect 7780 11350 8020 11590
rect 8110 11350 8350 11590
rect 8440 11350 8680 11590
rect 8770 11350 9010 11590
rect 9100 11350 9340 11590
rect 9430 11350 9670 11590
rect 9760 11350 10000 11590
rect 10090 11350 10330 11590
rect 10420 11350 10660 11590
rect 10750 11350 10990 11590
rect 11080 11350 11320 11590
rect 11410 11350 11650 11590
rect 11740 11350 11980 11590
rect 12070 11350 12310 11590
rect 12400 11350 12640 11590
rect 12730 11350 12970 11590
rect 13060 11350 13300 11590
rect 13390 11350 13630 11590
rect 13720 11350 13960 11590
rect 14050 11350 14290 11590
rect 14380 11350 14620 11590
rect 14710 11350 14950 11590
rect 15040 11350 15280 11590
rect 15370 11350 15610 11590
rect 15700 11350 15940 11590
rect 16030 11350 16270 11590
rect 16360 11350 16600 11590
rect 16690 11350 16930 11590
rect 17020 11350 17260 11590
rect 17350 11350 17590 11590
rect 17680 11350 17920 11590
rect 18010 11350 18250 11590
rect 18340 11350 18580 11590
rect 18670 11350 18910 11590
rect 19000 11350 19240 11590
rect 19330 11350 19570 11590
rect 7780 11020 8020 11260
rect 8110 11020 8350 11260
rect 8440 11020 8680 11260
rect 8770 11020 9010 11260
rect 9100 11020 9340 11260
rect 9430 11020 9670 11260
rect 9760 11020 10000 11260
rect 10090 11020 10330 11260
rect 10420 11020 10660 11260
rect 10750 11020 10990 11260
rect 11080 11020 11320 11260
rect 11410 11020 11650 11260
rect 11740 11020 11980 11260
rect 12070 11020 12310 11260
rect 12400 11020 12640 11260
rect 12730 11020 12970 11260
rect 13060 11020 13300 11260
rect 13390 11020 13630 11260
rect 13720 11020 13960 11260
rect 14050 11020 14290 11260
rect 14380 11020 14620 11260
rect 14710 11020 14950 11260
rect 15040 11020 15280 11260
rect 15370 11020 15610 11260
rect 15700 11020 15940 11260
rect 16030 11020 16270 11260
rect 16360 11020 16600 11260
rect 16690 11020 16930 11260
rect 17020 11020 17260 11260
rect 17350 11020 17590 11260
rect 17680 11020 17920 11260
rect 18010 11020 18250 11260
rect 18340 11020 18580 11260
rect 18670 11020 18910 11260
rect 19000 11020 19240 11260
rect 19330 11020 19570 11260
rect 7780 10690 8020 10930
rect 8110 10690 8350 10930
rect 8440 10690 8680 10930
rect 8770 10690 9010 10930
rect 9100 10690 9340 10930
rect 9430 10690 9670 10930
rect 9760 10690 10000 10930
rect 10090 10690 10330 10930
rect 10420 10690 10660 10930
rect 10750 10690 10990 10930
rect 11080 10690 11320 10930
rect 11410 10690 11650 10930
rect 11740 10690 11980 10930
rect 12070 10690 12310 10930
rect 12400 10690 12640 10930
rect 12730 10690 12970 10930
rect 13060 10690 13300 10930
rect 13390 10690 13630 10930
rect 13720 10690 13960 10930
rect 14050 10690 14290 10930
rect 14380 10690 14620 10930
rect 14710 10690 14950 10930
rect 15040 10690 15280 10930
rect 15370 10690 15610 10930
rect 15700 10690 15940 10930
rect 16030 10690 16270 10930
rect 16360 10690 16600 10930
rect 16690 10690 16930 10930
rect 17020 10690 17260 10930
rect 17350 10690 17590 10930
rect 17680 10690 17920 10930
rect 18010 10690 18250 10930
rect 18340 10690 18580 10930
rect 18670 10690 18910 10930
rect 19000 10690 19240 10930
rect 19330 10690 19570 10930
rect 7780 10360 8020 10600
rect 8110 10360 8350 10600
rect 8440 10360 8680 10600
rect 8770 10360 9010 10600
rect 9100 10360 9340 10600
rect 9430 10360 9670 10600
rect 9760 10360 10000 10600
rect 10090 10360 10330 10600
rect 10420 10360 10660 10600
rect 10750 10360 10990 10600
rect 11080 10360 11320 10600
rect 11410 10360 11650 10600
rect 11740 10360 11980 10600
rect 12070 10360 12310 10600
rect 12400 10360 12640 10600
rect 12730 10360 12970 10600
rect 13060 10360 13300 10600
rect 13390 10360 13630 10600
rect 13720 10360 13960 10600
rect 14050 10360 14290 10600
rect 14380 10360 14620 10600
rect 14710 10360 14950 10600
rect 15040 10360 15280 10600
rect 15370 10360 15610 10600
rect 15700 10360 15940 10600
rect 16030 10360 16270 10600
rect 16360 10360 16600 10600
rect 16690 10360 16930 10600
rect 17020 10360 17260 10600
rect 17350 10360 17590 10600
rect 17680 10360 17920 10600
rect 18010 10360 18250 10600
rect 18340 10360 18580 10600
rect 18670 10360 18910 10600
rect 19000 10360 19240 10600
rect 19330 10360 19570 10600
rect 7780 10030 8020 10270
rect 8110 10030 8350 10270
rect 8440 10030 8680 10270
rect 8770 10030 9010 10270
rect 9100 10030 9340 10270
rect 9430 10030 9670 10270
rect 9760 10030 10000 10270
rect 10090 10030 10330 10270
rect 10420 10030 10660 10270
rect 10750 10030 10990 10270
rect 11080 10030 11320 10270
rect 11410 10030 11650 10270
rect 11740 10030 11980 10270
rect 12070 10030 12310 10270
rect 12400 10030 12640 10270
rect 12730 10030 12970 10270
rect 13060 10030 13300 10270
rect 13390 10030 13630 10270
rect 13720 10030 13960 10270
rect 14050 10030 14290 10270
rect 14380 10030 14620 10270
rect 14710 10030 14950 10270
rect 15040 10030 15280 10270
rect 15370 10030 15610 10270
rect 15700 10030 15940 10270
rect 16030 10030 16270 10270
rect 16360 10030 16600 10270
rect 16690 10030 16930 10270
rect 17020 10030 17260 10270
rect 17350 10030 17590 10270
rect 17680 10030 17920 10270
rect 18010 10030 18250 10270
rect 18340 10030 18580 10270
rect 18670 10030 18910 10270
rect 19000 10030 19240 10270
rect 19330 10030 19570 10270
rect 7780 9700 8020 9940
rect 8110 9700 8350 9940
rect 8440 9700 8680 9940
rect 8770 9700 9010 9940
rect 9100 9700 9340 9940
rect 9430 9700 9670 9940
rect 9760 9700 10000 9940
rect 10090 9700 10330 9940
rect 10420 9700 10660 9940
rect 10750 9700 10990 9940
rect 11080 9700 11320 9940
rect 11410 9700 11650 9940
rect 11740 9700 11980 9940
rect 12070 9700 12310 9940
rect 12400 9700 12640 9940
rect 12730 9700 12970 9940
rect 13060 9700 13300 9940
rect 13390 9700 13630 9940
rect 13720 9700 13960 9940
rect 14050 9700 14290 9940
rect 14380 9700 14620 9940
rect 14710 9700 14950 9940
rect 15040 9700 15280 9940
rect 15370 9700 15610 9940
rect 15700 9700 15940 9940
rect 16030 9700 16270 9940
rect 16360 9700 16600 9940
rect 16690 9700 16930 9940
rect 17020 9700 17260 9940
rect 17350 9700 17590 9940
rect 17680 9700 17920 9940
rect 18010 9700 18250 9940
rect 18340 9700 18580 9940
rect 18670 9700 18910 9940
rect 19000 9700 19240 9940
rect 19330 9700 19570 9940
rect 7780 9370 8020 9610
rect 8110 9370 8350 9610
rect 8440 9370 8680 9610
rect 8770 9370 9010 9610
rect 9100 9370 9340 9610
rect 9430 9370 9670 9610
rect 9760 9370 10000 9610
rect 10090 9370 10330 9610
rect 10420 9370 10660 9610
rect 10750 9370 10990 9610
rect 11080 9370 11320 9610
rect 11410 9370 11650 9610
rect 11740 9370 11980 9610
rect 12070 9370 12310 9610
rect 12400 9370 12640 9610
rect 12730 9370 12970 9610
rect 13060 9370 13300 9610
rect 13390 9370 13630 9610
rect 13720 9370 13960 9610
rect 14050 9370 14290 9610
rect 14380 9370 14620 9610
rect 14710 9370 14950 9610
rect 15040 9370 15280 9610
rect 15370 9370 15610 9610
rect 15700 9370 15940 9610
rect 16030 9370 16270 9610
rect 16360 9370 16600 9610
rect 16690 9370 16930 9610
rect 17020 9370 17260 9610
rect 17350 9370 17590 9610
rect 17680 9370 17920 9610
rect 18010 9370 18250 9610
rect 18340 9370 18580 9610
rect 18670 9370 18910 9610
rect 19000 9370 19240 9610
rect 19330 9370 19570 9610
rect 7780 9040 8020 9280
rect 8110 9040 8350 9280
rect 8440 9040 8680 9280
rect 8770 9040 9010 9280
rect 9100 9040 9340 9280
rect 9430 9040 9670 9280
rect 9760 9040 10000 9280
rect 10090 9040 10330 9280
rect 10420 9040 10660 9280
rect 10750 9040 10990 9280
rect 11080 9040 11320 9280
rect 11410 9040 11650 9280
rect 11740 9040 11980 9280
rect 12070 9040 12310 9280
rect 12400 9040 12640 9280
rect 12730 9040 12970 9280
rect 13060 9040 13300 9280
rect 13390 9040 13630 9280
rect 13720 9040 13960 9280
rect 14050 9040 14290 9280
rect 14380 9040 14620 9280
rect 14710 9040 14950 9280
rect 15040 9040 15280 9280
rect 15370 9040 15610 9280
rect 15700 9040 15940 9280
rect 16030 9040 16270 9280
rect 16360 9040 16600 9280
rect 16690 9040 16930 9280
rect 17020 9040 17260 9280
rect 17350 9040 17590 9280
rect 17680 9040 17920 9280
rect 18010 9040 18250 9280
rect 18340 9040 18580 9280
rect 18670 9040 18910 9280
rect 19000 9040 19240 9280
rect 19330 9040 19570 9280
rect 31180 7590 31420 7830
rect 31510 7590 31750 7830
rect 31840 7590 32080 7830
rect 32170 7590 32410 7830
rect 32500 7590 32740 7830
rect 32830 7590 33070 7830
rect 33160 7590 33400 7830
rect 33490 7590 33730 7830
rect 33820 7590 34060 7830
rect 34150 7590 34390 7830
rect 34480 7590 34720 7830
rect 34810 7590 35050 7830
rect 35140 7590 35380 7830
rect 35470 7590 35710 7830
rect 35800 7590 36040 7830
rect 36130 7590 36370 7830
rect 36460 7590 36700 7830
rect 36790 7590 37030 7830
rect 37120 7590 37360 7830
rect 37450 7590 37690 7830
rect 31180 7260 31420 7500
rect 31510 7260 31750 7500
rect 31840 7260 32080 7500
rect 32170 7260 32410 7500
rect 32500 7260 32740 7500
rect 32830 7260 33070 7500
rect 33160 7260 33400 7500
rect 33490 7260 33730 7500
rect 33820 7260 34060 7500
rect 34150 7260 34390 7500
rect 34480 7260 34720 7500
rect 34810 7260 35050 7500
rect 35140 7260 35380 7500
rect 35470 7260 35710 7500
rect 35800 7260 36040 7500
rect 36130 7260 36370 7500
rect 36460 7260 36700 7500
rect 36790 7260 37030 7500
rect 37120 7260 37360 7500
rect 37450 7260 37690 7500
rect 31180 6930 31420 7170
rect 31510 6930 31750 7170
rect 31840 6930 32080 7170
rect 32170 6930 32410 7170
rect 32500 6930 32740 7170
rect 32830 6930 33070 7170
rect 33160 6930 33400 7170
rect 33490 6930 33730 7170
rect 33820 6930 34060 7170
rect 34150 6930 34390 7170
rect 34480 6930 34720 7170
rect 34810 6930 35050 7170
rect 35140 6930 35380 7170
rect 35470 6930 35710 7170
rect 35800 6930 36040 7170
rect 36130 6930 36370 7170
rect 36460 6930 36700 7170
rect 36790 6930 37030 7170
rect 37120 6930 37360 7170
rect 37450 6930 37690 7170
rect 31180 6600 31420 6840
rect 31510 6600 31750 6840
rect 31840 6600 32080 6840
rect 32170 6600 32410 6840
rect 32500 6600 32740 6840
rect 32830 6600 33070 6840
rect 33160 6600 33400 6840
rect 33490 6600 33730 6840
rect 33820 6600 34060 6840
rect 34150 6600 34390 6840
rect 34480 6600 34720 6840
rect 34810 6600 35050 6840
rect 35140 6600 35380 6840
rect 35470 6600 35710 6840
rect 35800 6600 36040 6840
rect 36130 6600 36370 6840
rect 36460 6600 36700 6840
rect 36790 6600 37030 6840
rect 37120 6600 37360 6840
rect 37450 6600 37690 6840
rect 31180 6270 31420 6510
rect 31510 6270 31750 6510
rect 31840 6270 32080 6510
rect 32170 6270 32410 6510
rect 32500 6270 32740 6510
rect 32830 6270 33070 6510
rect 33160 6270 33400 6510
rect 33490 6270 33730 6510
rect 33820 6270 34060 6510
rect 34150 6270 34390 6510
rect 34480 6270 34720 6510
rect 34810 6270 35050 6510
rect 35140 6270 35380 6510
rect 35470 6270 35710 6510
rect 35800 6270 36040 6510
rect 36130 6270 36370 6510
rect 36460 6270 36700 6510
rect 36790 6270 37030 6510
rect 37120 6270 37360 6510
rect 37450 6270 37690 6510
rect 31180 5940 31420 6180
rect 31510 5940 31750 6180
rect 31840 5940 32080 6180
rect 32170 5940 32410 6180
rect 32500 5940 32740 6180
rect 32830 5940 33070 6180
rect 33160 5940 33400 6180
rect 33490 5940 33730 6180
rect 33820 5940 34060 6180
rect 34150 5940 34390 6180
rect 34480 5940 34720 6180
rect 34810 5940 35050 6180
rect 35140 5940 35380 6180
rect 35470 5940 35710 6180
rect 35800 5940 36040 6180
rect 36130 5940 36370 6180
rect 36460 5940 36700 6180
rect 36790 5940 37030 6180
rect 37120 5940 37360 6180
rect 37450 5940 37690 6180
rect 31180 5610 31420 5850
rect 31510 5610 31750 5850
rect 31840 5610 32080 5850
rect 32170 5610 32410 5850
rect 32500 5610 32740 5850
rect 32830 5610 33070 5850
rect 33160 5610 33400 5850
rect 33490 5610 33730 5850
rect 33820 5610 34060 5850
rect 34150 5610 34390 5850
rect 34480 5610 34720 5850
rect 34810 5610 35050 5850
rect 35140 5610 35380 5850
rect 35470 5610 35710 5850
rect 35800 5610 36040 5850
rect 36130 5610 36370 5850
rect 36460 5610 36700 5850
rect 36790 5610 37030 5850
rect 37120 5610 37360 5850
rect 37450 5610 37690 5850
rect 31180 5280 31420 5520
rect 31510 5280 31750 5520
rect 31840 5280 32080 5520
rect 32170 5280 32410 5520
rect 32500 5280 32740 5520
rect 32830 5280 33070 5520
rect 33160 5280 33400 5520
rect 33490 5280 33730 5520
rect 33820 5280 34060 5520
rect 34150 5280 34390 5520
rect 34480 5280 34720 5520
rect 34810 5280 35050 5520
rect 35140 5280 35380 5520
rect 35470 5280 35710 5520
rect 35800 5280 36040 5520
rect 36130 5280 36370 5520
rect 36460 5280 36700 5520
rect 36790 5280 37030 5520
rect 37120 5280 37360 5520
rect 37450 5280 37690 5520
rect 31180 4950 31420 5190
rect 31510 4950 31750 5190
rect 31840 4950 32080 5190
rect 32170 4950 32410 5190
rect 32500 4950 32740 5190
rect 32830 4950 33070 5190
rect 33160 4950 33400 5190
rect 33490 4950 33730 5190
rect 33820 4950 34060 5190
rect 34150 4950 34390 5190
rect 34480 4950 34720 5190
rect 34810 4950 35050 5190
rect 35140 4950 35380 5190
rect 35470 4950 35710 5190
rect 35800 4950 36040 5190
rect 36130 4950 36370 5190
rect 36460 4950 36700 5190
rect 36790 4950 37030 5190
rect 37120 4950 37360 5190
rect 37450 4950 37690 5190
rect 31180 4620 31420 4860
rect 31510 4620 31750 4860
rect 31840 4620 32080 4860
rect 32170 4620 32410 4860
rect 32500 4620 32740 4860
rect 32830 4620 33070 4860
rect 33160 4620 33400 4860
rect 33490 4620 33730 4860
rect 33820 4620 34060 4860
rect 34150 4620 34390 4860
rect 34480 4620 34720 4860
rect 34810 4620 35050 4860
rect 35140 4620 35380 4860
rect 35470 4620 35710 4860
rect 35800 4620 36040 4860
rect 36130 4620 36370 4860
rect 36460 4620 36700 4860
rect 36790 4620 37030 4860
rect 37120 4620 37360 4860
rect 37450 4620 37690 4860
rect 31180 4290 31420 4530
rect 31510 4290 31750 4530
rect 31840 4290 32080 4530
rect 32170 4290 32410 4530
rect 32500 4290 32740 4530
rect 32830 4290 33070 4530
rect 33160 4290 33400 4530
rect 33490 4290 33730 4530
rect 33820 4290 34060 4530
rect 34150 4290 34390 4530
rect 34480 4290 34720 4530
rect 34810 4290 35050 4530
rect 35140 4290 35380 4530
rect 35470 4290 35710 4530
rect 35800 4290 36040 4530
rect 36130 4290 36370 4530
rect 36460 4290 36700 4530
rect 36790 4290 37030 4530
rect 37120 4290 37360 4530
rect 37450 4290 37690 4530
rect 31180 3960 31420 4200
rect 31510 3960 31750 4200
rect 31840 3960 32080 4200
rect 32170 3960 32410 4200
rect 32500 3960 32740 4200
rect 32830 3960 33070 4200
rect 33160 3960 33400 4200
rect 33490 3960 33730 4200
rect 33820 3960 34060 4200
rect 34150 3960 34390 4200
rect 34480 3960 34720 4200
rect 34810 3960 35050 4200
rect 35140 3960 35380 4200
rect 35470 3960 35710 4200
rect 35800 3960 36040 4200
rect 36130 3960 36370 4200
rect 36460 3960 36700 4200
rect 36790 3960 37030 4200
rect 37120 3960 37360 4200
rect 37450 3960 37690 4200
rect 31180 3630 31420 3870
rect 31510 3630 31750 3870
rect 31840 3630 32080 3870
rect 32170 3630 32410 3870
rect 32500 3630 32740 3870
rect 32830 3630 33070 3870
rect 33160 3630 33400 3870
rect 33490 3630 33730 3870
rect 33820 3630 34060 3870
rect 34150 3630 34390 3870
rect 34480 3630 34720 3870
rect 34810 3630 35050 3870
rect 35140 3630 35380 3870
rect 35470 3630 35710 3870
rect 35800 3630 36040 3870
rect 36130 3630 36370 3870
rect 36460 3630 36700 3870
rect 36790 3630 37030 3870
rect 37120 3630 37360 3870
rect 37450 3630 37690 3870
rect 31180 3300 31420 3540
rect 31510 3300 31750 3540
rect 31840 3300 32080 3540
rect 32170 3300 32410 3540
rect 32500 3300 32740 3540
rect 32830 3300 33070 3540
rect 33160 3300 33400 3540
rect 33490 3300 33730 3540
rect 33820 3300 34060 3540
rect 34150 3300 34390 3540
rect 34480 3300 34720 3540
rect 34810 3300 35050 3540
rect 35140 3300 35380 3540
rect 35470 3300 35710 3540
rect 35800 3300 36040 3540
rect 36130 3300 36370 3540
rect 36460 3300 36700 3540
rect 36790 3300 37030 3540
rect 37120 3300 37360 3540
rect 37450 3300 37690 3540
rect 31180 2970 31420 3210
rect 31510 2970 31750 3210
rect 31840 2970 32080 3210
rect 32170 2970 32410 3210
rect 32500 2970 32740 3210
rect 32830 2970 33070 3210
rect 33160 2970 33400 3210
rect 33490 2970 33730 3210
rect 33820 2970 34060 3210
rect 34150 2970 34390 3210
rect 34480 2970 34720 3210
rect 34810 2970 35050 3210
rect 35140 2970 35380 3210
rect 35470 2970 35710 3210
rect 35800 2970 36040 3210
rect 36130 2970 36370 3210
rect 36460 2970 36700 3210
rect 36790 2970 37030 3210
rect 37120 2970 37360 3210
rect 37450 2970 37690 3210
rect 31180 2640 31420 2880
rect 31510 2640 31750 2880
rect 31840 2640 32080 2880
rect 32170 2640 32410 2880
rect 32500 2640 32740 2880
rect 32830 2640 33070 2880
rect 33160 2640 33400 2880
rect 33490 2640 33730 2880
rect 33820 2640 34060 2880
rect 34150 2640 34390 2880
rect 34480 2640 34720 2880
rect 34810 2640 35050 2880
rect 35140 2640 35380 2880
rect 35470 2640 35710 2880
rect 35800 2640 36040 2880
rect 36130 2640 36370 2880
rect 36460 2640 36700 2880
rect 36790 2640 37030 2880
rect 37120 2640 37360 2880
rect 37450 2640 37690 2880
rect 31180 2310 31420 2550
rect 31510 2310 31750 2550
rect 31840 2310 32080 2550
rect 32170 2310 32410 2550
rect 32500 2310 32740 2550
rect 32830 2310 33070 2550
rect 33160 2310 33400 2550
rect 33490 2310 33730 2550
rect 33820 2310 34060 2550
rect 34150 2310 34390 2550
rect 34480 2310 34720 2550
rect 34810 2310 35050 2550
rect 35140 2310 35380 2550
rect 35470 2310 35710 2550
rect 35800 2310 36040 2550
rect 36130 2310 36370 2550
rect 36460 2310 36700 2550
rect 36790 2310 37030 2550
rect 37120 2310 37360 2550
rect 37450 2310 37690 2550
rect 31180 1980 31420 2220
rect 31510 1980 31750 2220
rect 31840 1980 32080 2220
rect 32170 1980 32410 2220
rect 32500 1980 32740 2220
rect 32830 1980 33070 2220
rect 33160 1980 33400 2220
rect 33490 1980 33730 2220
rect 33820 1980 34060 2220
rect 34150 1980 34390 2220
rect 34480 1980 34720 2220
rect 34810 1980 35050 2220
rect 35140 1980 35380 2220
rect 35470 1980 35710 2220
rect 35800 1980 36040 2220
rect 36130 1980 36370 2220
rect 36460 1980 36700 2220
rect 36790 1980 37030 2220
rect 37120 1980 37360 2220
rect 37450 1980 37690 2220
rect 31180 1650 31420 1890
rect 31510 1650 31750 1890
rect 31840 1650 32080 1890
rect 32170 1650 32410 1890
rect 32500 1650 32740 1890
rect 32830 1650 33070 1890
rect 33160 1650 33400 1890
rect 33490 1650 33730 1890
rect 33820 1650 34060 1890
rect 34150 1650 34390 1890
rect 34480 1650 34720 1890
rect 34810 1650 35050 1890
rect 35140 1650 35380 1890
rect 35470 1650 35710 1890
rect 35800 1650 36040 1890
rect 36130 1650 36370 1890
rect 36460 1650 36700 1890
rect 36790 1650 37030 1890
rect 37120 1650 37360 1890
rect 37450 1650 37690 1890
rect 31180 1320 31420 1560
rect 31510 1320 31750 1560
rect 31840 1320 32080 1560
rect 32170 1320 32410 1560
rect 32500 1320 32740 1560
rect 32830 1320 33070 1560
rect 33160 1320 33400 1560
rect 33490 1320 33730 1560
rect 33820 1320 34060 1560
rect 34150 1320 34390 1560
rect 34480 1320 34720 1560
rect 34810 1320 35050 1560
rect 35140 1320 35380 1560
rect 35470 1320 35710 1560
rect 35800 1320 36040 1560
rect 36130 1320 36370 1560
rect 36460 1320 36700 1560
rect 36790 1320 37030 1560
rect 37120 1320 37360 1560
rect 37450 1320 37690 1560
rect 31180 -10 31420 230
rect 31510 -10 31750 230
rect 31840 -10 32080 230
rect 32170 -10 32410 230
rect 32500 -10 32740 230
rect 32830 -10 33070 230
rect 33160 -10 33400 230
rect 33490 -10 33730 230
rect 33820 -10 34060 230
rect 34150 -10 34390 230
rect 34480 -10 34720 230
rect 34810 -10 35050 230
rect 35140 -10 35380 230
rect 35470 -10 35710 230
rect 35800 -10 36040 230
rect 36130 -10 36370 230
rect 36460 -10 36700 230
rect 36790 -10 37030 230
rect 37120 -10 37360 230
rect 37450 -10 37690 230
rect 31180 -340 31420 -100
rect 31510 -340 31750 -100
rect 31840 -340 32080 -100
rect 32170 -340 32410 -100
rect 32500 -340 32740 -100
rect 32830 -340 33070 -100
rect 33160 -340 33400 -100
rect 33490 -340 33730 -100
rect 33820 -340 34060 -100
rect 34150 -340 34390 -100
rect 34480 -340 34720 -100
rect 34810 -340 35050 -100
rect 35140 -340 35380 -100
rect 35470 -340 35710 -100
rect 35800 -340 36040 -100
rect 36130 -340 36370 -100
rect 36460 -340 36700 -100
rect 36790 -340 37030 -100
rect 37120 -340 37360 -100
rect 37450 -340 37690 -100
rect 31180 -670 31420 -430
rect 31510 -670 31750 -430
rect 31840 -670 32080 -430
rect 32170 -670 32410 -430
rect 32500 -670 32740 -430
rect 32830 -670 33070 -430
rect 33160 -670 33400 -430
rect 33490 -670 33730 -430
rect 33820 -670 34060 -430
rect 34150 -670 34390 -430
rect 34480 -670 34720 -430
rect 34810 -670 35050 -430
rect 35140 -670 35380 -430
rect 35470 -670 35710 -430
rect 35800 -670 36040 -430
rect 36130 -670 36370 -430
rect 36460 -670 36700 -430
rect 36790 -670 37030 -430
rect 37120 -670 37360 -430
rect 37450 -670 37690 -430
rect 31180 -1000 31420 -760
rect 31510 -1000 31750 -760
rect 31840 -1000 32080 -760
rect 32170 -1000 32410 -760
rect 32500 -1000 32740 -760
rect 32830 -1000 33070 -760
rect 33160 -1000 33400 -760
rect 33490 -1000 33730 -760
rect 33820 -1000 34060 -760
rect 34150 -1000 34390 -760
rect 34480 -1000 34720 -760
rect 34810 -1000 35050 -760
rect 35140 -1000 35380 -760
rect 35470 -1000 35710 -760
rect 35800 -1000 36040 -760
rect 36130 -1000 36370 -760
rect 36460 -1000 36700 -760
rect 36790 -1000 37030 -760
rect 37120 -1000 37360 -760
rect 37450 -1000 37690 -760
rect 31180 -1330 31420 -1090
rect 31510 -1330 31750 -1090
rect 31840 -1330 32080 -1090
rect 32170 -1330 32410 -1090
rect 32500 -1330 32740 -1090
rect 32830 -1330 33070 -1090
rect 33160 -1330 33400 -1090
rect 33490 -1330 33730 -1090
rect 33820 -1330 34060 -1090
rect 34150 -1330 34390 -1090
rect 34480 -1330 34720 -1090
rect 34810 -1330 35050 -1090
rect 35140 -1330 35380 -1090
rect 35470 -1330 35710 -1090
rect 35800 -1330 36040 -1090
rect 36130 -1330 36370 -1090
rect 36460 -1330 36700 -1090
rect 36790 -1330 37030 -1090
rect 37120 -1330 37360 -1090
rect 37450 -1330 37690 -1090
rect 31180 -1660 31420 -1420
rect 31510 -1660 31750 -1420
rect 31840 -1660 32080 -1420
rect 32170 -1660 32410 -1420
rect 32500 -1660 32740 -1420
rect 32830 -1660 33070 -1420
rect 33160 -1660 33400 -1420
rect 33490 -1660 33730 -1420
rect 33820 -1660 34060 -1420
rect 34150 -1660 34390 -1420
rect 34480 -1660 34720 -1420
rect 34810 -1660 35050 -1420
rect 35140 -1660 35380 -1420
rect 35470 -1660 35710 -1420
rect 35800 -1660 36040 -1420
rect 36130 -1660 36370 -1420
rect 36460 -1660 36700 -1420
rect 36790 -1660 37030 -1420
rect 37120 -1660 37360 -1420
rect 37450 -1660 37690 -1420
rect 31180 -1990 31420 -1750
rect 31510 -1990 31750 -1750
rect 31840 -1990 32080 -1750
rect 32170 -1990 32410 -1750
rect 32500 -1990 32740 -1750
rect 32830 -1990 33070 -1750
rect 33160 -1990 33400 -1750
rect 33490 -1990 33730 -1750
rect 33820 -1990 34060 -1750
rect 34150 -1990 34390 -1750
rect 34480 -1990 34720 -1750
rect 34810 -1990 35050 -1750
rect 35140 -1990 35380 -1750
rect 35470 -1990 35710 -1750
rect 35800 -1990 36040 -1750
rect 36130 -1990 36370 -1750
rect 36460 -1990 36700 -1750
rect 36790 -1990 37030 -1750
rect 37120 -1990 37360 -1750
rect 37450 -1990 37690 -1750
rect 31180 -2320 31420 -2080
rect 31510 -2320 31750 -2080
rect 31840 -2320 32080 -2080
rect 32170 -2320 32410 -2080
rect 32500 -2320 32740 -2080
rect 32830 -2320 33070 -2080
rect 33160 -2320 33400 -2080
rect 33490 -2320 33730 -2080
rect 33820 -2320 34060 -2080
rect 34150 -2320 34390 -2080
rect 34480 -2320 34720 -2080
rect 34810 -2320 35050 -2080
rect 35140 -2320 35380 -2080
rect 35470 -2320 35710 -2080
rect 35800 -2320 36040 -2080
rect 36130 -2320 36370 -2080
rect 36460 -2320 36700 -2080
rect 36790 -2320 37030 -2080
rect 37120 -2320 37360 -2080
rect 37450 -2320 37690 -2080
rect 31180 -2650 31420 -2410
rect 31510 -2650 31750 -2410
rect 31840 -2650 32080 -2410
rect 32170 -2650 32410 -2410
rect 32500 -2650 32740 -2410
rect 32830 -2650 33070 -2410
rect 33160 -2650 33400 -2410
rect 33490 -2650 33730 -2410
rect 33820 -2650 34060 -2410
rect 34150 -2650 34390 -2410
rect 34480 -2650 34720 -2410
rect 34810 -2650 35050 -2410
rect 35140 -2650 35380 -2410
rect 35470 -2650 35710 -2410
rect 35800 -2650 36040 -2410
rect 36130 -2650 36370 -2410
rect 36460 -2650 36700 -2410
rect 36790 -2650 37030 -2410
rect 37120 -2650 37360 -2410
rect 37450 -2650 37690 -2410
rect 31180 -2980 31420 -2740
rect 31510 -2980 31750 -2740
rect 31840 -2980 32080 -2740
rect 32170 -2980 32410 -2740
rect 32500 -2980 32740 -2740
rect 32830 -2980 33070 -2740
rect 33160 -2980 33400 -2740
rect 33490 -2980 33730 -2740
rect 33820 -2980 34060 -2740
rect 34150 -2980 34390 -2740
rect 34480 -2980 34720 -2740
rect 34810 -2980 35050 -2740
rect 35140 -2980 35380 -2740
rect 35470 -2980 35710 -2740
rect 35800 -2980 36040 -2740
rect 36130 -2980 36370 -2740
rect 36460 -2980 36700 -2740
rect 36790 -2980 37030 -2740
rect 37120 -2980 37360 -2740
rect 37450 -2980 37690 -2740
rect 31180 -3310 31420 -3070
rect 31510 -3310 31750 -3070
rect 31840 -3310 32080 -3070
rect 32170 -3310 32410 -3070
rect 32500 -3310 32740 -3070
rect 32830 -3310 33070 -3070
rect 33160 -3310 33400 -3070
rect 33490 -3310 33730 -3070
rect 33820 -3310 34060 -3070
rect 34150 -3310 34390 -3070
rect 34480 -3310 34720 -3070
rect 34810 -3310 35050 -3070
rect 35140 -3310 35380 -3070
rect 35470 -3310 35710 -3070
rect 35800 -3310 36040 -3070
rect 36130 -3310 36370 -3070
rect 36460 -3310 36700 -3070
rect 36790 -3310 37030 -3070
rect 37120 -3310 37360 -3070
rect 37450 -3310 37690 -3070
rect 31180 -3640 31420 -3400
rect 31510 -3640 31750 -3400
rect 31840 -3640 32080 -3400
rect 32170 -3640 32410 -3400
rect 32500 -3640 32740 -3400
rect 32830 -3640 33070 -3400
rect 33160 -3640 33400 -3400
rect 33490 -3640 33730 -3400
rect 33820 -3640 34060 -3400
rect 34150 -3640 34390 -3400
rect 34480 -3640 34720 -3400
rect 34810 -3640 35050 -3400
rect 35140 -3640 35380 -3400
rect 35470 -3640 35710 -3400
rect 35800 -3640 36040 -3400
rect 36130 -3640 36370 -3400
rect 36460 -3640 36700 -3400
rect 36790 -3640 37030 -3400
rect 37120 -3640 37360 -3400
rect 37450 -3640 37690 -3400
rect 31180 -3970 31420 -3730
rect 31510 -3970 31750 -3730
rect 31840 -3970 32080 -3730
rect 32170 -3970 32410 -3730
rect 32500 -3970 32740 -3730
rect 32830 -3970 33070 -3730
rect 33160 -3970 33400 -3730
rect 33490 -3970 33730 -3730
rect 33820 -3970 34060 -3730
rect 34150 -3970 34390 -3730
rect 34480 -3970 34720 -3730
rect 34810 -3970 35050 -3730
rect 35140 -3970 35380 -3730
rect 35470 -3970 35710 -3730
rect 35800 -3970 36040 -3730
rect 36130 -3970 36370 -3730
rect 36460 -3970 36700 -3730
rect 36790 -3970 37030 -3730
rect 37120 -3970 37360 -3730
rect 37450 -3970 37690 -3730
rect 31180 -4300 31420 -4060
rect 31510 -4300 31750 -4060
rect 31840 -4300 32080 -4060
rect 32170 -4300 32410 -4060
rect 32500 -4300 32740 -4060
rect 32830 -4300 33070 -4060
rect 33160 -4300 33400 -4060
rect 33490 -4300 33730 -4060
rect 33820 -4300 34060 -4060
rect 34150 -4300 34390 -4060
rect 34480 -4300 34720 -4060
rect 34810 -4300 35050 -4060
rect 35140 -4300 35380 -4060
rect 35470 -4300 35710 -4060
rect 35800 -4300 36040 -4060
rect 36130 -4300 36370 -4060
rect 36460 -4300 36700 -4060
rect 36790 -4300 37030 -4060
rect 37120 -4300 37360 -4060
rect 37450 -4300 37690 -4060
rect 31180 -4630 31420 -4390
rect 31510 -4630 31750 -4390
rect 31840 -4630 32080 -4390
rect 32170 -4630 32410 -4390
rect 32500 -4630 32740 -4390
rect 32830 -4630 33070 -4390
rect 33160 -4630 33400 -4390
rect 33490 -4630 33730 -4390
rect 33820 -4630 34060 -4390
rect 34150 -4630 34390 -4390
rect 34480 -4630 34720 -4390
rect 34810 -4630 35050 -4390
rect 35140 -4630 35380 -4390
rect 35470 -4630 35710 -4390
rect 35800 -4630 36040 -4390
rect 36130 -4630 36370 -4390
rect 36460 -4630 36700 -4390
rect 36790 -4630 37030 -4390
rect 37120 -4630 37360 -4390
rect 37450 -4630 37690 -4390
rect -1180 -5080 -940 -4840
rect -850 -5080 -610 -4840
rect -520 -5080 -280 -4840
rect -190 -5080 50 -4840
rect -1180 -5410 -940 -5170
rect -850 -5410 -610 -5170
rect -520 -5410 -280 -5170
rect -190 -5410 50 -5170
rect -1180 -5740 -940 -5500
rect -850 -5740 -610 -5500
rect -520 -5740 -280 -5500
rect -190 -5740 50 -5500
rect -1180 -6070 -940 -5830
rect -850 -6070 -610 -5830
rect -520 -6070 -280 -5830
rect -190 -6070 50 -5830
rect 14730 -5080 14970 -4840
rect 15060 -5080 15300 -4840
rect 15390 -5080 15630 -4840
rect 15720 -5080 15960 -4840
rect 14730 -5410 14970 -5170
rect 15060 -5410 15300 -5170
rect 15390 -5410 15630 -5170
rect 15720 -5410 15960 -5170
rect 14730 -5740 14970 -5500
rect 15060 -5740 15300 -5500
rect 15390 -5740 15630 -5500
rect 15720 -5740 15960 -5500
rect 14730 -6070 14970 -5830
rect 15060 -6070 15300 -5830
rect 15390 -6070 15630 -5830
rect 15720 -6070 15960 -5830
rect 31180 -4960 31420 -4720
rect 31510 -4960 31750 -4720
rect 31840 -4960 32080 -4720
rect 32170 -4960 32410 -4720
rect 32500 -4960 32740 -4720
rect 32830 -4960 33070 -4720
rect 33160 -4960 33400 -4720
rect 33490 -4960 33730 -4720
rect 33820 -4960 34060 -4720
rect 34150 -4960 34390 -4720
rect 34480 -4960 34720 -4720
rect 34810 -4960 35050 -4720
rect 35140 -4960 35380 -4720
rect 35470 -4960 35710 -4720
rect 35800 -4960 36040 -4720
rect 36130 -4960 36370 -4720
rect 36460 -4960 36700 -4720
rect 36790 -4960 37030 -4720
rect 37120 -4960 37360 -4720
rect 37450 -4960 37690 -4720
rect 31180 -5290 31420 -5050
rect 31510 -5290 31750 -5050
rect 31840 -5290 32080 -5050
rect 32170 -5290 32410 -5050
rect 32500 -5290 32740 -5050
rect 32830 -5290 33070 -5050
rect 33160 -5290 33400 -5050
rect 33490 -5290 33730 -5050
rect 33820 -5290 34060 -5050
rect 34150 -5290 34390 -5050
rect 34480 -5290 34720 -5050
rect 34810 -5290 35050 -5050
rect 35140 -5290 35380 -5050
rect 35470 -5290 35710 -5050
rect 35800 -5290 36040 -5050
rect 36130 -5290 36370 -5050
rect 36460 -5290 36700 -5050
rect 36790 -5290 37030 -5050
rect 37120 -5290 37360 -5050
rect 37450 -5290 37690 -5050
rect 31180 -5620 31420 -5380
rect 31510 -5620 31750 -5380
rect 31840 -5620 32080 -5380
rect 32170 -5620 32410 -5380
rect 32500 -5620 32740 -5380
rect 32830 -5620 33070 -5380
rect 33160 -5620 33400 -5380
rect 33490 -5620 33730 -5380
rect 33820 -5620 34060 -5380
rect 34150 -5620 34390 -5380
rect 34480 -5620 34720 -5380
rect 34810 -5620 35050 -5380
rect 35140 -5620 35380 -5380
rect 35470 -5620 35710 -5380
rect 35800 -5620 36040 -5380
rect 36130 -5620 36370 -5380
rect 36460 -5620 36700 -5380
rect 36790 -5620 37030 -5380
rect 37120 -5620 37360 -5380
rect 37450 -5620 37690 -5380
rect 31180 -5950 31420 -5710
rect 31510 -5950 31750 -5710
rect 31840 -5950 32080 -5710
rect 32170 -5950 32410 -5710
rect 32500 -5950 32740 -5710
rect 32830 -5950 33070 -5710
rect 33160 -5950 33400 -5710
rect 33490 -5950 33730 -5710
rect 33820 -5950 34060 -5710
rect 34150 -5950 34390 -5710
rect 34480 -5950 34720 -5710
rect 34810 -5950 35050 -5710
rect 35140 -5950 35380 -5710
rect 35470 -5950 35710 -5710
rect 35800 -5950 36040 -5710
rect 36130 -5950 36370 -5710
rect 36460 -5950 36700 -5710
rect 36790 -5950 37030 -5710
rect 37120 -5950 37360 -5710
rect 37450 -5950 37690 -5710
rect 31180 -6280 31420 -6040
rect 31510 -6280 31750 -6040
rect 31840 -6280 32080 -6040
rect 32170 -6280 32410 -6040
rect 32500 -6280 32740 -6040
rect 32830 -6280 33070 -6040
rect 33160 -6280 33400 -6040
rect 33490 -6280 33730 -6040
rect 33820 -6280 34060 -6040
rect 34150 -6280 34390 -6040
rect 34480 -6280 34720 -6040
rect 34810 -6280 35050 -6040
rect 35140 -6280 35380 -6040
rect 35470 -6280 35710 -6040
rect 35800 -6280 36040 -6040
rect 36130 -6280 36370 -6040
rect 36460 -6280 36700 -6040
rect 36790 -6280 37030 -6040
rect 37120 -6280 37360 -6040
rect 37450 -6280 37690 -6040
<< metal5 >>
rect -5020 21610 7290 21640
rect -5020 21370 -4650 21610
rect -4410 21370 -4320 21610
rect -4080 21370 -3990 21610
rect -3750 21370 -3660 21610
rect -3420 21370 -3330 21610
rect -3090 21370 -3000 21610
rect -2760 21370 -2670 21610
rect -2430 21370 -2340 21610
rect -2100 21370 -2010 21610
rect -1770 21370 -1640 21610
rect -1400 21370 -1310 21610
rect -1070 21370 -980 21610
rect -740 21370 -650 21610
rect -410 21370 -320 21610
rect -80 21370 10 21610
rect 250 21370 340 21610
rect 580 21370 670 21610
rect 910 21370 1000 21610
rect 1240 21370 1370 21610
rect 1610 21370 1700 21610
rect 1940 21370 2030 21610
rect 2270 21370 2360 21610
rect 2600 21370 2690 21610
rect 2930 21370 3020 21610
rect 3260 21370 3350 21610
rect 3590 21370 3680 21610
rect 3920 21370 4010 21610
rect 4250 21370 4380 21610
rect 4620 21370 4710 21610
rect 4950 21370 5040 21610
rect 5280 21370 5370 21610
rect 5610 21370 5700 21610
rect 5940 21370 6030 21610
rect 6270 21370 6360 21610
rect 6600 21370 6690 21610
rect 6930 21370 7020 21610
rect 7260 21370 7290 21610
rect -5020 20830 7290 21370
rect -5020 20590 -4670 20830
rect -4430 20590 -4340 20830
rect -4100 20590 -4010 20830
rect -3770 20590 -3680 20830
rect -3440 20590 -3350 20830
rect -3110 20590 -3020 20830
rect -2780 20590 -2690 20830
rect -2450 20590 -2360 20830
rect -2120 20590 -2030 20830
rect -1790 20590 -1700 20830
rect -1460 20590 -1370 20830
rect -1130 20590 -1040 20830
rect -800 20590 -710 20830
rect -470 20590 -380 20830
rect -140 20590 -50 20830
rect 190 20590 280 20830
rect 520 20590 610 20830
rect 850 20590 940 20830
rect 1180 20590 1270 20830
rect 1510 20590 1600 20830
rect 1840 20590 1930 20830
rect 2170 20590 2260 20830
rect 2500 20590 2590 20830
rect 2830 20590 2920 20830
rect 3160 20590 3250 20830
rect 3490 20590 3580 20830
rect 3820 20590 3910 20830
rect 4150 20590 4240 20830
rect 4480 20590 4570 20830
rect 4810 20590 4900 20830
rect 5140 20590 5230 20830
rect 5470 20590 5560 20830
rect 5800 20590 5890 20830
rect 6130 20590 6220 20830
rect 6460 20590 6550 20830
rect 6790 20590 6880 20830
rect 7120 20590 7290 20830
rect -5020 20500 7290 20590
rect -5020 20260 -4670 20500
rect -4430 20260 -4340 20500
rect -4100 20260 -4010 20500
rect -3770 20260 -3680 20500
rect -3440 20260 -3350 20500
rect -3110 20260 -3020 20500
rect -2780 20260 -2690 20500
rect -2450 20260 -2360 20500
rect -2120 20260 -2030 20500
rect -1790 20260 -1700 20500
rect -1460 20260 -1370 20500
rect -1130 20260 -1040 20500
rect -800 20260 -710 20500
rect -470 20260 -380 20500
rect -140 20260 -50 20500
rect 190 20260 280 20500
rect 520 20260 610 20500
rect 850 20260 940 20500
rect 1180 20260 1270 20500
rect 1510 20260 1600 20500
rect 1840 20260 1930 20500
rect 2170 20260 2260 20500
rect 2500 20260 2590 20500
rect 2830 20260 2920 20500
rect 3160 20260 3250 20500
rect 3490 20260 3580 20500
rect 3820 20260 3910 20500
rect 4150 20260 4240 20500
rect 4480 20260 4570 20500
rect 4810 20260 4900 20500
rect 5140 20260 5230 20500
rect 5470 20260 5560 20500
rect 5800 20260 5890 20500
rect 6130 20260 6220 20500
rect 6460 20260 6550 20500
rect 6790 20260 6880 20500
rect 7120 20260 7290 20500
rect -5020 20170 7290 20260
rect -5020 19930 -4670 20170
rect -4430 19930 -4340 20170
rect -4100 19930 -4010 20170
rect -3770 19930 -3680 20170
rect -3440 19930 -3350 20170
rect -3110 19930 -3020 20170
rect -2780 19930 -2690 20170
rect -2450 19930 -2360 20170
rect -2120 19930 -2030 20170
rect -1790 19930 -1700 20170
rect -1460 19930 -1370 20170
rect -1130 19930 -1040 20170
rect -800 19930 -710 20170
rect -470 19930 -380 20170
rect -140 19930 -50 20170
rect 190 19930 280 20170
rect 520 19930 610 20170
rect 850 19930 940 20170
rect 1180 19930 1270 20170
rect 1510 19930 1600 20170
rect 1840 19930 1930 20170
rect 2170 19930 2260 20170
rect 2500 19930 2590 20170
rect 2830 19930 2920 20170
rect 3160 19930 3250 20170
rect 3490 19930 3580 20170
rect 3820 19930 3910 20170
rect 4150 19930 4240 20170
rect 4480 19930 4570 20170
rect 4810 19930 4900 20170
rect 5140 19930 5230 20170
rect 5470 19930 5560 20170
rect 5800 19930 5890 20170
rect 6130 19930 6220 20170
rect 6460 19930 6550 20170
rect 6790 19930 6880 20170
rect 7120 19930 7290 20170
rect -5020 19840 7290 19930
rect -5020 19600 -4670 19840
rect -4430 19600 -4340 19840
rect -4100 19600 -4010 19840
rect -3770 19600 -3680 19840
rect -3440 19600 -3350 19840
rect -3110 19600 -3020 19840
rect -2780 19600 -2690 19840
rect -2450 19600 -2360 19840
rect -2120 19600 -2030 19840
rect -1790 19600 -1700 19840
rect -1460 19600 -1370 19840
rect -1130 19600 -1040 19840
rect -800 19600 -710 19840
rect -470 19600 -380 19840
rect -140 19600 -50 19840
rect 190 19600 280 19840
rect 520 19600 610 19840
rect 850 19600 940 19840
rect 1180 19600 1270 19840
rect 1510 19600 1600 19840
rect 1840 19600 1930 19840
rect 2170 19600 2260 19840
rect 2500 19600 2590 19840
rect 2830 19600 2920 19840
rect 3160 19600 3250 19840
rect 3490 19600 3580 19840
rect 3820 19600 3910 19840
rect 4150 19600 4240 19840
rect 4480 19600 4570 19840
rect 4810 19600 4900 19840
rect 5140 19600 5230 19840
rect 5470 19600 5560 19840
rect 5800 19600 5890 19840
rect 6130 19600 6220 19840
rect 6460 19600 6550 19840
rect 6790 19600 6880 19840
rect 7120 19600 7290 19840
rect -5020 19510 7290 19600
rect -5020 19270 -4670 19510
rect -4430 19270 -4340 19510
rect -4100 19270 -4010 19510
rect -3770 19270 -3680 19510
rect -3440 19270 -3350 19510
rect -3110 19270 -3020 19510
rect -2780 19270 -2690 19510
rect -2450 19270 -2360 19510
rect -2120 19270 -2030 19510
rect -1790 19270 -1700 19510
rect -1460 19270 -1370 19510
rect -1130 19270 -1040 19510
rect -800 19270 -710 19510
rect -470 19270 -380 19510
rect -140 19270 -50 19510
rect 190 19270 280 19510
rect 520 19270 610 19510
rect 850 19270 940 19510
rect 1180 19270 1270 19510
rect 1510 19270 1600 19510
rect 1840 19270 1930 19510
rect 2170 19270 2260 19510
rect 2500 19270 2590 19510
rect 2830 19270 2920 19510
rect 3160 19270 3250 19510
rect 3490 19270 3580 19510
rect 3820 19270 3910 19510
rect 4150 19270 4240 19510
rect 4480 19270 4570 19510
rect 4810 19270 4900 19510
rect 5140 19270 5230 19510
rect 5470 19270 5560 19510
rect 5800 19270 5890 19510
rect 6130 19270 6220 19510
rect 6460 19270 6550 19510
rect 6790 19270 6880 19510
rect 7120 19270 7290 19510
rect -5020 19180 7290 19270
rect -5020 18940 -4670 19180
rect -4430 18940 -4340 19180
rect -4100 18940 -4010 19180
rect -3770 18940 -3680 19180
rect -3440 18940 -3350 19180
rect -3110 18940 -3020 19180
rect -2780 18940 -2690 19180
rect -2450 18940 -2360 19180
rect -2120 18940 -2030 19180
rect -1790 18940 -1700 19180
rect -1460 18940 -1370 19180
rect -1130 18940 -1040 19180
rect -800 18940 -710 19180
rect -470 18940 -380 19180
rect -140 18940 -50 19180
rect 190 18940 280 19180
rect 520 18940 610 19180
rect 850 18940 940 19180
rect 1180 18940 1270 19180
rect 1510 18940 1600 19180
rect 1840 18940 1930 19180
rect 2170 18940 2260 19180
rect 2500 18940 2590 19180
rect 2830 18940 2920 19180
rect 3160 18940 3250 19180
rect 3490 18940 3580 19180
rect 3820 18940 3910 19180
rect 4150 18940 4240 19180
rect 4480 18940 4570 19180
rect 4810 18940 4900 19180
rect 5140 18940 5230 19180
rect 5470 18940 5560 19180
rect 5800 18940 5890 19180
rect 6130 18940 6220 19180
rect 6460 18940 6550 19180
rect 6790 18940 6880 19180
rect 7120 18940 7290 19180
rect -5020 18850 7290 18940
rect -5020 18610 -4670 18850
rect -4430 18610 -4340 18850
rect -4100 18610 -4010 18850
rect -3770 18610 -3680 18850
rect -3440 18610 -3350 18850
rect -3110 18610 -3020 18850
rect -2780 18610 -2690 18850
rect -2450 18610 -2360 18850
rect -2120 18610 -2030 18850
rect -1790 18610 -1700 18850
rect -1460 18610 -1370 18850
rect -1130 18610 -1040 18850
rect -800 18610 -710 18850
rect -470 18610 -380 18850
rect -140 18610 -50 18850
rect 190 18610 280 18850
rect 520 18610 610 18850
rect 850 18610 940 18850
rect 1180 18610 1270 18850
rect 1510 18610 1600 18850
rect 1840 18610 1930 18850
rect 2170 18610 2260 18850
rect 2500 18610 2590 18850
rect 2830 18610 2920 18850
rect 3160 18610 3250 18850
rect 3490 18610 3580 18850
rect 3820 18610 3910 18850
rect 4150 18610 4240 18850
rect 4480 18610 4570 18850
rect 4810 18610 4900 18850
rect 5140 18610 5230 18850
rect 5470 18610 5560 18850
rect 5800 18610 5890 18850
rect 6130 18610 6220 18850
rect 6460 18610 6550 18850
rect 6790 18610 6880 18850
rect 7120 18610 7290 18850
rect -5020 18520 7290 18610
rect -5020 18280 -4670 18520
rect -4430 18280 -4340 18520
rect -4100 18280 -4010 18520
rect -3770 18280 -3680 18520
rect -3440 18280 -3350 18520
rect -3110 18280 -3020 18520
rect -2780 18280 -2690 18520
rect -2450 18280 -2360 18520
rect -2120 18280 -2030 18520
rect -1790 18280 -1700 18520
rect -1460 18280 -1370 18520
rect -1130 18280 -1040 18520
rect -800 18280 -710 18520
rect -470 18280 -380 18520
rect -140 18280 -50 18520
rect 190 18280 280 18520
rect 520 18280 610 18520
rect 850 18280 940 18520
rect 1180 18280 1270 18520
rect 1510 18280 1600 18520
rect 1840 18280 1930 18520
rect 2170 18280 2260 18520
rect 2500 18280 2590 18520
rect 2830 18280 2920 18520
rect 3160 18280 3250 18520
rect 3490 18280 3580 18520
rect 3820 18280 3910 18520
rect 4150 18280 4240 18520
rect 4480 18280 4570 18520
rect 4810 18280 4900 18520
rect 5140 18280 5230 18520
rect 5470 18280 5560 18520
rect 5800 18280 5890 18520
rect 6130 18280 6220 18520
rect 6460 18280 6550 18520
rect 6790 18280 6880 18520
rect 7120 18280 7290 18520
rect -5020 18190 7290 18280
rect -5020 17950 -4670 18190
rect -4430 17950 -4340 18190
rect -4100 17950 -4010 18190
rect -3770 17950 -3680 18190
rect -3440 17950 -3350 18190
rect -3110 17950 -3020 18190
rect -2780 17950 -2690 18190
rect -2450 17950 -2360 18190
rect -2120 17950 -2030 18190
rect -1790 17950 -1700 18190
rect -1460 17950 -1370 18190
rect -1130 17950 -1040 18190
rect -800 17950 -710 18190
rect -470 17950 -380 18190
rect -140 17950 -50 18190
rect 190 17950 280 18190
rect 520 17950 610 18190
rect 850 17950 940 18190
rect 1180 17950 1270 18190
rect 1510 17950 1600 18190
rect 1840 17950 1930 18190
rect 2170 17950 2260 18190
rect 2500 17950 2590 18190
rect 2830 17950 2920 18190
rect 3160 17950 3250 18190
rect 3490 17950 3580 18190
rect 3820 17950 3910 18190
rect 4150 17950 4240 18190
rect 4480 17950 4570 18190
rect 4810 17950 4900 18190
rect 5140 17950 5230 18190
rect 5470 17950 5560 18190
rect 5800 17950 5890 18190
rect 6130 17950 6220 18190
rect 6460 17950 6550 18190
rect 6790 17950 6880 18190
rect 7120 17950 7290 18190
rect -5020 17860 7290 17950
rect -5020 17620 -4670 17860
rect -4430 17620 -4340 17860
rect -4100 17620 -4010 17860
rect -3770 17620 -3680 17860
rect -3440 17620 -3350 17860
rect -3110 17620 -3020 17860
rect -2780 17620 -2690 17860
rect -2450 17620 -2360 17860
rect -2120 17620 -2030 17860
rect -1790 17620 -1700 17860
rect -1460 17620 -1370 17860
rect -1130 17620 -1040 17860
rect -800 17620 -710 17860
rect -470 17620 -380 17860
rect -140 17620 -50 17860
rect 190 17620 280 17860
rect 520 17620 610 17860
rect 850 17620 940 17860
rect 1180 17620 1270 17860
rect 1510 17620 1600 17860
rect 1840 17620 1930 17860
rect 2170 17620 2260 17860
rect 2500 17620 2590 17860
rect 2830 17620 2920 17860
rect 3160 17620 3250 17860
rect 3490 17620 3580 17860
rect 3820 17620 3910 17860
rect 4150 17620 4240 17860
rect 4480 17620 4570 17860
rect 4810 17620 4900 17860
rect 5140 17620 5230 17860
rect 5470 17620 5560 17860
rect 5800 17620 5890 17860
rect 6130 17620 6220 17860
rect 6460 17620 6550 17860
rect 6790 17620 6880 17860
rect 7120 17620 7290 17860
rect -5020 17530 7290 17620
rect -5020 17290 -4670 17530
rect -4430 17290 -4340 17530
rect -4100 17290 -4010 17530
rect -3770 17290 -3680 17530
rect -3440 17290 -3350 17530
rect -3110 17290 -3020 17530
rect -2780 17290 -2690 17530
rect -2450 17290 -2360 17530
rect -2120 17290 -2030 17530
rect -1790 17290 -1700 17530
rect -1460 17290 -1370 17530
rect -1130 17290 -1040 17530
rect -800 17290 -710 17530
rect -470 17290 -380 17530
rect -140 17290 -50 17530
rect 190 17290 280 17530
rect 520 17290 610 17530
rect 850 17290 940 17530
rect 1180 17290 1270 17530
rect 1510 17290 1600 17530
rect 1840 17290 1930 17530
rect 2170 17290 2260 17530
rect 2500 17290 2590 17530
rect 2830 17290 2920 17530
rect 3160 17290 3250 17530
rect 3490 17290 3580 17530
rect 3820 17290 3910 17530
rect 4150 17290 4240 17530
rect 4480 17290 4570 17530
rect 4810 17290 4900 17530
rect 5140 17290 5230 17530
rect 5470 17290 5560 17530
rect 5800 17290 5890 17530
rect 6130 17290 6220 17530
rect 6460 17290 6550 17530
rect 6790 17290 6880 17530
rect 7120 17290 7290 17530
rect -5020 17200 7290 17290
rect -5020 16960 -4670 17200
rect -4430 16960 -4340 17200
rect -4100 16960 -4010 17200
rect -3770 16960 -3680 17200
rect -3440 16960 -3350 17200
rect -3110 16960 -3020 17200
rect -2780 16960 -2690 17200
rect -2450 16960 -2360 17200
rect -2120 16960 -2030 17200
rect -1790 16960 -1700 17200
rect -1460 16960 -1370 17200
rect -1130 16960 -1040 17200
rect -800 16960 -710 17200
rect -470 16960 -380 17200
rect -140 16960 -50 17200
rect 190 16960 280 17200
rect 520 16960 610 17200
rect 850 16960 940 17200
rect 1180 16960 1270 17200
rect 1510 16960 1600 17200
rect 1840 16960 1930 17200
rect 2170 16960 2260 17200
rect 2500 16960 2590 17200
rect 2830 16960 2920 17200
rect 3160 16960 3250 17200
rect 3490 16960 3580 17200
rect 3820 16960 3910 17200
rect 4150 16960 4240 17200
rect 4480 16960 4570 17200
rect 4810 16960 4900 17200
rect 5140 16960 5230 17200
rect 5470 16960 5560 17200
rect 5800 16960 5890 17200
rect 6130 16960 6220 17200
rect 6460 16960 6550 17200
rect 6790 16960 6880 17200
rect 7120 16960 7290 17200
rect -5020 16870 7290 16960
rect -5020 16630 -4670 16870
rect -4430 16630 -4340 16870
rect -4100 16630 -4010 16870
rect -3770 16630 -3680 16870
rect -3440 16630 -3350 16870
rect -3110 16630 -3020 16870
rect -2780 16630 -2690 16870
rect -2450 16630 -2360 16870
rect -2120 16630 -2030 16870
rect -1790 16630 -1700 16870
rect -1460 16630 -1370 16870
rect -1130 16630 -1040 16870
rect -800 16630 -710 16870
rect -470 16630 -380 16870
rect -140 16630 -50 16870
rect 190 16630 280 16870
rect 520 16630 610 16870
rect 850 16630 940 16870
rect 1180 16630 1270 16870
rect 1510 16630 1600 16870
rect 1840 16630 1930 16870
rect 2170 16630 2260 16870
rect 2500 16630 2590 16870
rect 2830 16630 2920 16870
rect 3160 16630 3250 16870
rect 3490 16630 3580 16870
rect 3820 16630 3910 16870
rect 4150 16630 4240 16870
rect 4480 16630 4570 16870
rect 4810 16630 4900 16870
rect 5140 16630 5230 16870
rect 5470 16630 5560 16870
rect 5800 16630 5890 16870
rect 6130 16630 6220 16870
rect 6460 16630 6550 16870
rect 6790 16630 6880 16870
rect 7120 16630 7290 16870
rect -5020 16540 7290 16630
rect -5020 16300 -4670 16540
rect -4430 16300 -4340 16540
rect -4100 16300 -4010 16540
rect -3770 16300 -3680 16540
rect -3440 16300 -3350 16540
rect -3110 16300 -3020 16540
rect -2780 16300 -2690 16540
rect -2450 16300 -2360 16540
rect -2120 16300 -2030 16540
rect -1790 16300 -1700 16540
rect -1460 16300 -1370 16540
rect -1130 16300 -1040 16540
rect -800 16300 -710 16540
rect -470 16300 -380 16540
rect -140 16300 -50 16540
rect 190 16300 280 16540
rect 520 16300 610 16540
rect 850 16300 940 16540
rect 1180 16300 1270 16540
rect 1510 16300 1600 16540
rect 1840 16300 1930 16540
rect 2170 16300 2260 16540
rect 2500 16300 2590 16540
rect 2830 16300 2920 16540
rect 3160 16300 3250 16540
rect 3490 16300 3580 16540
rect 3820 16300 3910 16540
rect 4150 16300 4240 16540
rect 4480 16300 4570 16540
rect 4810 16300 4900 16540
rect 5140 16300 5230 16540
rect 5470 16300 5560 16540
rect 5800 16300 5890 16540
rect 6130 16300 6220 16540
rect 6460 16300 6550 16540
rect 6790 16300 6880 16540
rect 7120 16300 7290 16540
rect -5020 16210 7290 16300
rect -5020 15970 -4670 16210
rect -4430 15970 -4340 16210
rect -4100 15970 -4010 16210
rect -3770 15970 -3680 16210
rect -3440 15970 -3350 16210
rect -3110 15970 -3020 16210
rect -2780 15970 -2690 16210
rect -2450 15970 -2360 16210
rect -2120 15970 -2030 16210
rect -1790 15970 -1700 16210
rect -1460 15970 -1370 16210
rect -1130 15970 -1040 16210
rect -800 15970 -710 16210
rect -470 15970 -380 16210
rect -140 15970 -50 16210
rect 190 15970 280 16210
rect 520 15970 610 16210
rect 850 15970 940 16210
rect 1180 15970 1270 16210
rect 1510 15970 1600 16210
rect 1840 15970 1930 16210
rect 2170 15970 2260 16210
rect 2500 15970 2590 16210
rect 2830 15970 2920 16210
rect 3160 15970 3250 16210
rect 3490 15970 3580 16210
rect 3820 15970 3910 16210
rect 4150 15970 4240 16210
rect 4480 15970 4570 16210
rect 4810 15970 4900 16210
rect 5140 15970 5230 16210
rect 5470 15970 5560 16210
rect 5800 15970 5890 16210
rect 6130 15970 6220 16210
rect 6460 15970 6550 16210
rect 6790 15970 6880 16210
rect 7120 15970 7290 16210
rect -5020 15880 7290 15970
rect -5020 15640 -4670 15880
rect -4430 15640 -4340 15880
rect -4100 15640 -4010 15880
rect -3770 15640 -3680 15880
rect -3440 15640 -3350 15880
rect -3110 15640 -3020 15880
rect -2780 15640 -2690 15880
rect -2450 15640 -2360 15880
rect -2120 15640 -2030 15880
rect -1790 15640 -1700 15880
rect -1460 15640 -1370 15880
rect -1130 15640 -1040 15880
rect -800 15640 -710 15880
rect -470 15640 -380 15880
rect -140 15640 -50 15880
rect 190 15640 280 15880
rect 520 15640 610 15880
rect 850 15640 940 15880
rect 1180 15640 1270 15880
rect 1510 15640 1600 15880
rect 1840 15640 1930 15880
rect 2170 15640 2260 15880
rect 2500 15640 2590 15880
rect 2830 15640 2920 15880
rect 3160 15640 3250 15880
rect 3490 15640 3580 15880
rect 3820 15640 3910 15880
rect 4150 15640 4240 15880
rect 4480 15640 4570 15880
rect 4810 15640 4900 15880
rect 5140 15640 5230 15880
rect 5470 15640 5560 15880
rect 5800 15640 5890 15880
rect 6130 15640 6220 15880
rect 6460 15640 6550 15880
rect 6790 15640 6880 15880
rect 7120 15640 7290 15880
rect -5020 15550 7290 15640
rect -5020 15310 -4670 15550
rect -4430 15310 -4340 15550
rect -4100 15310 -4010 15550
rect -3770 15310 -3680 15550
rect -3440 15310 -3350 15550
rect -3110 15310 -3020 15550
rect -2780 15310 -2690 15550
rect -2450 15310 -2360 15550
rect -2120 15310 -2030 15550
rect -1790 15310 -1700 15550
rect -1460 15310 -1370 15550
rect -1130 15310 -1040 15550
rect -800 15310 -710 15550
rect -470 15310 -380 15550
rect -140 15310 -50 15550
rect 190 15310 280 15550
rect 520 15310 610 15550
rect 850 15310 940 15550
rect 1180 15310 1270 15550
rect 1510 15310 1600 15550
rect 1840 15310 1930 15550
rect 2170 15310 2260 15550
rect 2500 15310 2590 15550
rect 2830 15310 2920 15550
rect 3160 15310 3250 15550
rect 3490 15310 3580 15550
rect 3820 15310 3910 15550
rect 4150 15310 4240 15550
rect 4480 15310 4570 15550
rect 4810 15310 4900 15550
rect 5140 15310 5230 15550
rect 5470 15310 5560 15550
rect 5800 15310 5890 15550
rect 6130 15310 6220 15550
rect 6460 15310 6550 15550
rect 6790 15310 6880 15550
rect 7120 15310 7290 15550
rect -5020 15220 7290 15310
rect -5020 14980 -4670 15220
rect -4430 14980 -4340 15220
rect -4100 14980 -4010 15220
rect -3770 14980 -3680 15220
rect -3440 14980 -3350 15220
rect -3110 14980 -3020 15220
rect -2780 14980 -2690 15220
rect -2450 14980 -2360 15220
rect -2120 14980 -2030 15220
rect -1790 14980 -1700 15220
rect -1460 14980 -1370 15220
rect -1130 14980 -1040 15220
rect -800 14980 -710 15220
rect -470 14980 -380 15220
rect -140 14980 -50 15220
rect 190 14980 280 15220
rect 520 14980 610 15220
rect 850 14980 940 15220
rect 1180 14980 1270 15220
rect 1510 14980 1600 15220
rect 1840 14980 1930 15220
rect 2170 14980 2260 15220
rect 2500 14980 2590 15220
rect 2830 14980 2920 15220
rect 3160 14980 3250 15220
rect 3490 14980 3580 15220
rect 3820 14980 3910 15220
rect 4150 14980 4240 15220
rect 4480 14980 4570 15220
rect 4810 14980 4900 15220
rect 5140 14980 5230 15220
rect 5470 14980 5560 15220
rect 5800 14980 5890 15220
rect 6130 14980 6220 15220
rect 6460 14980 6550 15220
rect 6790 14980 6880 15220
rect 7120 14980 7290 15220
rect -5020 14890 7290 14980
rect -5020 14650 -4670 14890
rect -4430 14650 -4340 14890
rect -4100 14650 -4010 14890
rect -3770 14650 -3680 14890
rect -3440 14650 -3350 14890
rect -3110 14650 -3020 14890
rect -2780 14650 -2690 14890
rect -2450 14650 -2360 14890
rect -2120 14650 -2030 14890
rect -1790 14650 -1700 14890
rect -1460 14650 -1370 14890
rect -1130 14650 -1040 14890
rect -800 14650 -710 14890
rect -470 14650 -380 14890
rect -140 14650 -50 14890
rect 190 14650 280 14890
rect 520 14650 610 14890
rect 850 14650 940 14890
rect 1180 14650 1270 14890
rect 1510 14650 1600 14890
rect 1840 14650 1930 14890
rect 2170 14650 2260 14890
rect 2500 14650 2590 14890
rect 2830 14650 2920 14890
rect 3160 14650 3250 14890
rect 3490 14650 3580 14890
rect 3820 14650 3910 14890
rect 4150 14650 4240 14890
rect 4480 14650 4570 14890
rect 4810 14650 4900 14890
rect 5140 14650 5230 14890
rect 5470 14650 5560 14890
rect 5800 14650 5890 14890
rect 6130 14650 6220 14890
rect 6460 14650 6550 14890
rect 6790 14650 6880 14890
rect 7120 14650 7290 14890
rect -5020 14560 7290 14650
rect -5020 14320 -4670 14560
rect -4430 14320 -4340 14560
rect -4100 14320 -4010 14560
rect -3770 14320 -3680 14560
rect -3440 14320 -3350 14560
rect -3110 14320 -3020 14560
rect -2780 14320 -2690 14560
rect -2450 14320 -2360 14560
rect -2120 14320 -2030 14560
rect -1790 14320 -1700 14560
rect -1460 14320 -1370 14560
rect -1130 14320 -1040 14560
rect -800 14320 -710 14560
rect -470 14320 -380 14560
rect -140 14320 -50 14560
rect 190 14320 280 14560
rect 520 14320 610 14560
rect 850 14320 940 14560
rect 1180 14320 1270 14560
rect 1510 14320 1600 14560
rect 1840 14320 1930 14560
rect 2170 14320 2260 14560
rect 2500 14320 2590 14560
rect 2830 14320 2920 14560
rect 3160 14320 3250 14560
rect 3490 14320 3580 14560
rect 3820 14320 3910 14560
rect 4150 14320 4240 14560
rect 4480 14320 4570 14560
rect 4810 14320 4900 14560
rect 5140 14320 5230 14560
rect 5470 14320 5560 14560
rect 5800 14320 5890 14560
rect 6130 14320 6220 14560
rect 6460 14320 6550 14560
rect 6790 14320 6880 14560
rect 7120 14320 7290 14560
rect -5020 14230 7290 14320
rect -5020 13990 -4670 14230
rect -4430 13990 -4340 14230
rect -4100 13990 -4010 14230
rect -3770 13990 -3680 14230
rect -3440 13990 -3350 14230
rect -3110 13990 -3020 14230
rect -2780 13990 -2690 14230
rect -2450 13990 -2360 14230
rect -2120 13990 -2030 14230
rect -1790 13990 -1700 14230
rect -1460 13990 -1370 14230
rect -1130 13990 -1040 14230
rect -800 13990 -710 14230
rect -470 13990 -380 14230
rect -140 13990 -50 14230
rect 190 13990 280 14230
rect 520 13990 610 14230
rect 850 13990 940 14230
rect 1180 13990 1270 14230
rect 1510 13990 1600 14230
rect 1840 13990 1930 14230
rect 2170 13990 2260 14230
rect 2500 13990 2590 14230
rect 2830 13990 2920 14230
rect 3160 13990 3250 14230
rect 3490 13990 3580 14230
rect 3820 13990 3910 14230
rect 4150 13990 4240 14230
rect 4480 13990 4570 14230
rect 4810 13990 4900 14230
rect 5140 13990 5230 14230
rect 5470 13990 5560 14230
rect 5800 13990 5890 14230
rect 6130 13990 6220 14230
rect 6460 13990 6550 14230
rect 6790 13990 6880 14230
rect 7120 13990 7290 14230
rect -5020 13900 7290 13990
rect -5020 13660 -4670 13900
rect -4430 13660 -4340 13900
rect -4100 13660 -4010 13900
rect -3770 13660 -3680 13900
rect -3440 13660 -3350 13900
rect -3110 13660 -3020 13900
rect -2780 13660 -2690 13900
rect -2450 13660 -2360 13900
rect -2120 13660 -2030 13900
rect -1790 13660 -1700 13900
rect -1460 13660 -1370 13900
rect -1130 13660 -1040 13900
rect -800 13660 -710 13900
rect -470 13660 -380 13900
rect -140 13660 -50 13900
rect 190 13660 280 13900
rect 520 13660 610 13900
rect 850 13660 940 13900
rect 1180 13660 1270 13900
rect 1510 13660 1600 13900
rect 1840 13660 1930 13900
rect 2170 13660 2260 13900
rect 2500 13660 2590 13900
rect 2830 13660 2920 13900
rect 3160 13660 3250 13900
rect 3490 13660 3580 13900
rect 3820 13660 3910 13900
rect 4150 13660 4240 13900
rect 4480 13660 4570 13900
rect 4810 13660 4900 13900
rect 5140 13660 5230 13900
rect 5470 13660 5560 13900
rect 5800 13660 5890 13900
rect 6130 13660 6220 13900
rect 6460 13660 6550 13900
rect 6790 13660 6880 13900
rect 7120 13660 7290 13900
rect -5020 13570 7290 13660
rect -5020 13330 -4670 13570
rect -4430 13330 -4340 13570
rect -4100 13330 -4010 13570
rect -3770 13330 -3680 13570
rect -3440 13330 -3350 13570
rect -3110 13330 -3020 13570
rect -2780 13330 -2690 13570
rect -2450 13330 -2360 13570
rect -2120 13330 -2030 13570
rect -1790 13330 -1700 13570
rect -1460 13330 -1370 13570
rect -1130 13330 -1040 13570
rect -800 13330 -710 13570
rect -470 13330 -380 13570
rect -140 13330 -50 13570
rect 190 13330 280 13570
rect 520 13330 610 13570
rect 850 13330 940 13570
rect 1180 13330 1270 13570
rect 1510 13330 1600 13570
rect 1840 13330 1930 13570
rect 2170 13330 2260 13570
rect 2500 13330 2590 13570
rect 2830 13330 2920 13570
rect 3160 13330 3250 13570
rect 3490 13330 3580 13570
rect 3820 13330 3910 13570
rect 4150 13330 4240 13570
rect 4480 13330 4570 13570
rect 4810 13330 4900 13570
rect 5140 13330 5230 13570
rect 5470 13330 5560 13570
rect 5800 13330 5890 13570
rect 6130 13330 6220 13570
rect 6460 13330 6550 13570
rect 6790 13330 6880 13570
rect 7120 13330 7290 13570
rect -5020 13240 7290 13330
rect -5020 13000 -4670 13240
rect -4430 13000 -4340 13240
rect -4100 13000 -4010 13240
rect -3770 13000 -3680 13240
rect -3440 13000 -3350 13240
rect -3110 13000 -3020 13240
rect -2780 13000 -2690 13240
rect -2450 13000 -2360 13240
rect -2120 13000 -2030 13240
rect -1790 13000 -1700 13240
rect -1460 13000 -1370 13240
rect -1130 13000 -1040 13240
rect -800 13000 -710 13240
rect -470 13000 -380 13240
rect -140 13000 -50 13240
rect 190 13000 280 13240
rect 520 13000 610 13240
rect 850 13000 940 13240
rect 1180 13000 1270 13240
rect 1510 13000 1600 13240
rect 1840 13000 1930 13240
rect 2170 13000 2260 13240
rect 2500 13000 2590 13240
rect 2830 13000 2920 13240
rect 3160 13000 3250 13240
rect 3490 13000 3580 13240
rect 3820 13000 3910 13240
rect 4150 13000 4240 13240
rect 4480 13000 4570 13240
rect 4810 13000 4900 13240
rect 5140 13000 5230 13240
rect 5470 13000 5560 13240
rect 5800 13000 5890 13240
rect 6130 13000 6220 13240
rect 6460 13000 6550 13240
rect 6790 13000 6880 13240
rect 7120 13000 7290 13240
rect -5020 12910 7290 13000
rect -5020 12670 -4670 12910
rect -4430 12670 -4340 12910
rect -4100 12670 -4010 12910
rect -3770 12670 -3680 12910
rect -3440 12670 -3350 12910
rect -3110 12670 -3020 12910
rect -2780 12670 -2690 12910
rect -2450 12670 -2360 12910
rect -2120 12670 -2030 12910
rect -1790 12670 -1700 12910
rect -1460 12670 -1370 12910
rect -1130 12670 -1040 12910
rect -800 12670 -710 12910
rect -470 12670 -380 12910
rect -140 12670 -50 12910
rect 190 12670 280 12910
rect 520 12670 610 12910
rect 850 12670 940 12910
rect 1180 12670 1270 12910
rect 1510 12670 1600 12910
rect 1840 12670 1930 12910
rect 2170 12670 2260 12910
rect 2500 12670 2590 12910
rect 2830 12670 2920 12910
rect 3160 12670 3250 12910
rect 3490 12670 3580 12910
rect 3820 12670 3910 12910
rect 4150 12670 4240 12910
rect 4480 12670 4570 12910
rect 4810 12670 4900 12910
rect 5140 12670 5230 12910
rect 5470 12670 5560 12910
rect 5800 12670 5890 12910
rect 6130 12670 6220 12910
rect 6460 12670 6550 12910
rect 6790 12670 6880 12910
rect 7120 12670 7290 12910
rect -5020 12580 7290 12670
rect -5020 12340 -4670 12580
rect -4430 12340 -4340 12580
rect -4100 12340 -4010 12580
rect -3770 12340 -3680 12580
rect -3440 12340 -3350 12580
rect -3110 12340 -3020 12580
rect -2780 12340 -2690 12580
rect -2450 12340 -2360 12580
rect -2120 12340 -2030 12580
rect -1790 12340 -1700 12580
rect -1460 12340 -1370 12580
rect -1130 12340 -1040 12580
rect -800 12340 -710 12580
rect -470 12340 -380 12580
rect -140 12340 -50 12580
rect 190 12340 280 12580
rect 520 12340 610 12580
rect 850 12340 940 12580
rect 1180 12340 1270 12580
rect 1510 12340 1600 12580
rect 1840 12340 1930 12580
rect 2170 12340 2260 12580
rect 2500 12340 2590 12580
rect 2830 12340 2920 12580
rect 3160 12340 3250 12580
rect 3490 12340 3580 12580
rect 3820 12340 3910 12580
rect 4150 12340 4240 12580
rect 4480 12340 4570 12580
rect 4810 12340 4900 12580
rect 5140 12340 5230 12580
rect 5470 12340 5560 12580
rect 5800 12340 5890 12580
rect 6130 12340 6220 12580
rect 6460 12340 6550 12580
rect 6790 12340 6880 12580
rect 7120 12340 7290 12580
rect -5020 12250 7290 12340
rect -5020 12010 -4670 12250
rect -4430 12010 -4340 12250
rect -4100 12010 -4010 12250
rect -3770 12010 -3680 12250
rect -3440 12010 -3350 12250
rect -3110 12010 -3020 12250
rect -2780 12010 -2690 12250
rect -2450 12010 -2360 12250
rect -2120 12010 -2030 12250
rect -1790 12010 -1700 12250
rect -1460 12010 -1370 12250
rect -1130 12010 -1040 12250
rect -800 12010 -710 12250
rect -470 12010 -380 12250
rect -140 12010 -50 12250
rect 190 12010 280 12250
rect 520 12010 610 12250
rect 850 12010 940 12250
rect 1180 12010 1270 12250
rect 1510 12010 1600 12250
rect 1840 12010 1930 12250
rect 2170 12010 2260 12250
rect 2500 12010 2590 12250
rect 2830 12010 2920 12250
rect 3160 12010 3250 12250
rect 3490 12010 3580 12250
rect 3820 12010 3910 12250
rect 4150 12010 4240 12250
rect 4480 12010 4570 12250
rect 4810 12010 4900 12250
rect 5140 12010 5230 12250
rect 5470 12010 5560 12250
rect 5800 12010 5890 12250
rect 6130 12010 6220 12250
rect 6460 12010 6550 12250
rect 6790 12010 6880 12250
rect 7120 12010 7290 12250
rect -5020 11920 7290 12010
rect -5020 11680 -4670 11920
rect -4430 11680 -4340 11920
rect -4100 11680 -4010 11920
rect -3770 11680 -3680 11920
rect -3440 11680 -3350 11920
rect -3110 11680 -3020 11920
rect -2780 11680 -2690 11920
rect -2450 11680 -2360 11920
rect -2120 11680 -2030 11920
rect -1790 11680 -1700 11920
rect -1460 11680 -1370 11920
rect -1130 11680 -1040 11920
rect -800 11680 -710 11920
rect -470 11680 -380 11920
rect -140 11680 -50 11920
rect 190 11680 280 11920
rect 520 11680 610 11920
rect 850 11680 940 11920
rect 1180 11680 1270 11920
rect 1510 11680 1600 11920
rect 1840 11680 1930 11920
rect 2170 11680 2260 11920
rect 2500 11680 2590 11920
rect 2830 11680 2920 11920
rect 3160 11680 3250 11920
rect 3490 11680 3580 11920
rect 3820 11680 3910 11920
rect 4150 11680 4240 11920
rect 4480 11680 4570 11920
rect 4810 11680 4900 11920
rect 5140 11680 5230 11920
rect 5470 11680 5560 11920
rect 5800 11680 5890 11920
rect 6130 11680 6220 11920
rect 6460 11680 6550 11920
rect 6790 11680 6880 11920
rect 7120 11680 7290 11920
rect -5020 11590 7290 11680
rect -5020 11350 -4670 11590
rect -4430 11350 -4340 11590
rect -4100 11350 -4010 11590
rect -3770 11350 -3680 11590
rect -3440 11350 -3350 11590
rect -3110 11350 -3020 11590
rect -2780 11350 -2690 11590
rect -2450 11350 -2360 11590
rect -2120 11350 -2030 11590
rect -1790 11350 -1700 11590
rect -1460 11350 -1370 11590
rect -1130 11350 -1040 11590
rect -800 11350 -710 11590
rect -470 11350 -380 11590
rect -140 11350 -50 11590
rect 190 11350 280 11590
rect 520 11350 610 11590
rect 850 11350 940 11590
rect 1180 11350 1270 11590
rect 1510 11350 1600 11590
rect 1840 11350 1930 11590
rect 2170 11350 2260 11590
rect 2500 11350 2590 11590
rect 2830 11350 2920 11590
rect 3160 11350 3250 11590
rect 3490 11350 3580 11590
rect 3820 11350 3910 11590
rect 4150 11350 4240 11590
rect 4480 11350 4570 11590
rect 4810 11350 4900 11590
rect 5140 11350 5230 11590
rect 5470 11350 5560 11590
rect 5800 11350 5890 11590
rect 6130 11350 6220 11590
rect 6460 11350 6550 11590
rect 6790 11350 6880 11590
rect 7120 11350 7290 11590
rect -5020 11260 7290 11350
rect -5020 11020 -4670 11260
rect -4430 11020 -4340 11260
rect -4100 11020 -4010 11260
rect -3770 11020 -3680 11260
rect -3440 11020 -3350 11260
rect -3110 11020 -3020 11260
rect -2780 11020 -2690 11260
rect -2450 11020 -2360 11260
rect -2120 11020 -2030 11260
rect -1790 11020 -1700 11260
rect -1460 11020 -1370 11260
rect -1130 11020 -1040 11260
rect -800 11020 -710 11260
rect -470 11020 -380 11260
rect -140 11020 -50 11260
rect 190 11020 280 11260
rect 520 11020 610 11260
rect 850 11020 940 11260
rect 1180 11020 1270 11260
rect 1510 11020 1600 11260
rect 1840 11020 1930 11260
rect 2170 11020 2260 11260
rect 2500 11020 2590 11260
rect 2830 11020 2920 11260
rect 3160 11020 3250 11260
rect 3490 11020 3580 11260
rect 3820 11020 3910 11260
rect 4150 11020 4240 11260
rect 4480 11020 4570 11260
rect 4810 11020 4900 11260
rect 5140 11020 5230 11260
rect 5470 11020 5560 11260
rect 5800 11020 5890 11260
rect 6130 11020 6220 11260
rect 6460 11020 6550 11260
rect 6790 11020 6880 11260
rect 7120 11020 7290 11260
rect -5020 10930 7290 11020
rect -5020 10690 -4670 10930
rect -4430 10690 -4340 10930
rect -4100 10690 -4010 10930
rect -3770 10690 -3680 10930
rect -3440 10690 -3350 10930
rect -3110 10690 -3020 10930
rect -2780 10690 -2690 10930
rect -2450 10690 -2360 10930
rect -2120 10690 -2030 10930
rect -1790 10690 -1700 10930
rect -1460 10690 -1370 10930
rect -1130 10690 -1040 10930
rect -800 10690 -710 10930
rect -470 10690 -380 10930
rect -140 10690 -50 10930
rect 190 10690 280 10930
rect 520 10690 610 10930
rect 850 10690 940 10930
rect 1180 10690 1270 10930
rect 1510 10690 1600 10930
rect 1840 10690 1930 10930
rect 2170 10690 2260 10930
rect 2500 10690 2590 10930
rect 2830 10690 2920 10930
rect 3160 10690 3250 10930
rect 3490 10690 3580 10930
rect 3820 10690 3910 10930
rect 4150 10690 4240 10930
rect 4480 10690 4570 10930
rect 4810 10690 4900 10930
rect 5140 10690 5230 10930
rect 5470 10690 5560 10930
rect 5800 10690 5890 10930
rect 6130 10690 6220 10930
rect 6460 10690 6550 10930
rect 6790 10690 6880 10930
rect 7120 10690 7290 10930
rect -5020 10600 7290 10690
rect -5020 10360 -4670 10600
rect -4430 10360 -4340 10600
rect -4100 10360 -4010 10600
rect -3770 10360 -3680 10600
rect -3440 10360 -3350 10600
rect -3110 10360 -3020 10600
rect -2780 10360 -2690 10600
rect -2450 10360 -2360 10600
rect -2120 10360 -2030 10600
rect -1790 10360 -1700 10600
rect -1460 10360 -1370 10600
rect -1130 10360 -1040 10600
rect -800 10360 -710 10600
rect -470 10360 -380 10600
rect -140 10360 -50 10600
rect 190 10360 280 10600
rect 520 10360 610 10600
rect 850 10360 940 10600
rect 1180 10360 1270 10600
rect 1510 10360 1600 10600
rect 1840 10360 1930 10600
rect 2170 10360 2260 10600
rect 2500 10360 2590 10600
rect 2830 10360 2920 10600
rect 3160 10360 3250 10600
rect 3490 10360 3580 10600
rect 3820 10360 3910 10600
rect 4150 10360 4240 10600
rect 4480 10360 4570 10600
rect 4810 10360 4900 10600
rect 5140 10360 5230 10600
rect 5470 10360 5560 10600
rect 5800 10360 5890 10600
rect 6130 10360 6220 10600
rect 6460 10360 6550 10600
rect 6790 10360 6880 10600
rect 7120 10360 7290 10600
rect -5020 10270 7290 10360
rect -5020 10030 -4670 10270
rect -4430 10030 -4340 10270
rect -4100 10030 -4010 10270
rect -3770 10030 -3680 10270
rect -3440 10030 -3350 10270
rect -3110 10030 -3020 10270
rect -2780 10030 -2690 10270
rect -2450 10030 -2360 10270
rect -2120 10030 -2030 10270
rect -1790 10030 -1700 10270
rect -1460 10030 -1370 10270
rect -1130 10030 -1040 10270
rect -800 10030 -710 10270
rect -470 10030 -380 10270
rect -140 10030 -50 10270
rect 190 10030 280 10270
rect 520 10030 610 10270
rect 850 10030 940 10270
rect 1180 10030 1270 10270
rect 1510 10030 1600 10270
rect 1840 10030 1930 10270
rect 2170 10030 2260 10270
rect 2500 10030 2590 10270
rect 2830 10030 2920 10270
rect 3160 10030 3250 10270
rect 3490 10030 3580 10270
rect 3820 10030 3910 10270
rect 4150 10030 4240 10270
rect 4480 10030 4570 10270
rect 4810 10030 4900 10270
rect 5140 10030 5230 10270
rect 5470 10030 5560 10270
rect 5800 10030 5890 10270
rect 6130 10030 6220 10270
rect 6460 10030 6550 10270
rect 6790 10030 6880 10270
rect 7120 10030 7290 10270
rect -5020 9940 7290 10030
rect -5020 9700 -4670 9940
rect -4430 9700 -4340 9940
rect -4100 9700 -4010 9940
rect -3770 9700 -3680 9940
rect -3440 9700 -3350 9940
rect -3110 9700 -3020 9940
rect -2780 9700 -2690 9940
rect -2450 9700 -2360 9940
rect -2120 9700 -2030 9940
rect -1790 9700 -1700 9940
rect -1460 9700 -1370 9940
rect -1130 9700 -1040 9940
rect -800 9700 -710 9940
rect -470 9700 -380 9940
rect -140 9700 -50 9940
rect 190 9700 280 9940
rect 520 9700 610 9940
rect 850 9700 940 9940
rect 1180 9700 1270 9940
rect 1510 9700 1600 9940
rect 1840 9700 1930 9940
rect 2170 9700 2260 9940
rect 2500 9700 2590 9940
rect 2830 9700 2920 9940
rect 3160 9700 3250 9940
rect 3490 9700 3580 9940
rect 3820 9700 3910 9940
rect 4150 9700 4240 9940
rect 4480 9700 4570 9940
rect 4810 9700 4900 9940
rect 5140 9700 5230 9940
rect 5470 9700 5560 9940
rect 5800 9700 5890 9940
rect 6130 9700 6220 9940
rect 6460 9700 6550 9940
rect 6790 9700 6880 9940
rect 7120 9700 7290 9940
rect -5020 9610 7290 9700
rect -5020 9370 -4670 9610
rect -4430 9370 -4340 9610
rect -4100 9370 -4010 9610
rect -3770 9370 -3680 9610
rect -3440 9370 -3350 9610
rect -3110 9370 -3020 9610
rect -2780 9370 -2690 9610
rect -2450 9370 -2360 9610
rect -2120 9370 -2030 9610
rect -1790 9370 -1700 9610
rect -1460 9370 -1370 9610
rect -1130 9370 -1040 9610
rect -800 9370 -710 9610
rect -470 9370 -380 9610
rect -140 9370 -50 9610
rect 190 9370 280 9610
rect 520 9370 610 9610
rect 850 9370 940 9610
rect 1180 9370 1270 9610
rect 1510 9370 1600 9610
rect 1840 9370 1930 9610
rect 2170 9370 2260 9610
rect 2500 9370 2590 9610
rect 2830 9370 2920 9610
rect 3160 9370 3250 9610
rect 3490 9370 3580 9610
rect 3820 9370 3910 9610
rect 4150 9370 4240 9610
rect 4480 9370 4570 9610
rect 4810 9370 4900 9610
rect 5140 9370 5230 9610
rect 5470 9370 5560 9610
rect 5800 9370 5890 9610
rect 6130 9370 6220 9610
rect 6460 9370 6550 9610
rect 6790 9370 6880 9610
rect 7120 9370 7290 9610
rect -5020 9280 7290 9370
rect -5020 9040 -4670 9280
rect -4430 9040 -4340 9280
rect -4100 9040 -4010 9280
rect -3770 9040 -3680 9280
rect -3440 9040 -3350 9280
rect -3110 9040 -3020 9280
rect -2780 9040 -2690 9280
rect -2450 9040 -2360 9280
rect -2120 9040 -2030 9280
rect -1790 9040 -1700 9280
rect -1460 9040 -1370 9280
rect -1130 9040 -1040 9280
rect -800 9040 -710 9280
rect -470 9040 -380 9280
rect -140 9040 -50 9280
rect 190 9040 280 9280
rect 520 9040 610 9280
rect 850 9040 940 9280
rect 1180 9040 1270 9280
rect 1510 9040 1600 9280
rect 1840 9040 1930 9280
rect 2170 9040 2260 9280
rect 2500 9040 2590 9280
rect 2830 9040 2920 9280
rect 3160 9040 3250 9280
rect 3490 9040 3580 9280
rect 3820 9040 3910 9280
rect 4150 9040 4240 9280
rect 4480 9040 4570 9280
rect 4810 9040 4900 9280
rect 5140 9040 5230 9280
rect 5470 9040 5560 9280
rect 5800 9040 5890 9280
rect 6130 9040 6220 9280
rect 6460 9040 6550 9280
rect 6790 9040 6880 9280
rect 7120 9040 7290 9280
rect -5020 8690 7290 9040
rect 7610 21610 19920 21640
rect 7610 21370 7640 21610
rect 7880 21370 7970 21610
rect 8210 21370 8300 21610
rect 8540 21370 8630 21610
rect 8870 21370 8960 21610
rect 9200 21370 9290 21610
rect 9530 21370 9620 21610
rect 9860 21370 9950 21610
rect 10190 21370 10280 21610
rect 10520 21370 10650 21610
rect 10890 21370 10980 21610
rect 11220 21370 11310 21610
rect 11550 21370 11640 21610
rect 11880 21370 11970 21610
rect 12210 21370 12300 21610
rect 12540 21370 12630 21610
rect 12870 21370 12960 21610
rect 13200 21370 13290 21610
rect 13530 21370 13660 21610
rect 13900 21370 13990 21610
rect 14230 21370 14320 21610
rect 14560 21370 14650 21610
rect 14890 21370 14980 21610
rect 15220 21370 15310 21610
rect 15550 21370 15640 21610
rect 15880 21370 15970 21610
rect 16210 21370 16300 21610
rect 16540 21370 16670 21610
rect 16910 21370 17000 21610
rect 17240 21370 17330 21610
rect 17570 21370 17660 21610
rect 17900 21370 17990 21610
rect 18230 21370 18320 21610
rect 18560 21370 18650 21610
rect 18890 21370 18980 21610
rect 19220 21370 19310 21610
rect 19550 21370 19920 21610
rect 7610 20830 19920 21370
rect 7610 20590 7780 20830
rect 8020 20590 8110 20830
rect 8350 20590 8440 20830
rect 8680 20590 8770 20830
rect 9010 20590 9100 20830
rect 9340 20590 9430 20830
rect 9670 20590 9760 20830
rect 10000 20590 10090 20830
rect 10330 20590 10420 20830
rect 10660 20590 10750 20830
rect 10990 20590 11080 20830
rect 11320 20590 11410 20830
rect 11650 20590 11740 20830
rect 11980 20590 12070 20830
rect 12310 20590 12400 20830
rect 12640 20590 12730 20830
rect 12970 20590 13060 20830
rect 13300 20590 13390 20830
rect 13630 20590 13720 20830
rect 13960 20590 14050 20830
rect 14290 20590 14380 20830
rect 14620 20590 14710 20830
rect 14950 20590 15040 20830
rect 15280 20590 15370 20830
rect 15610 20590 15700 20830
rect 15940 20590 16030 20830
rect 16270 20590 16360 20830
rect 16600 20590 16690 20830
rect 16930 20590 17020 20830
rect 17260 20590 17350 20830
rect 17590 20590 17680 20830
rect 17920 20590 18010 20830
rect 18250 20590 18340 20830
rect 18580 20590 18670 20830
rect 18910 20590 19000 20830
rect 19240 20590 19330 20830
rect 19570 20590 19920 20830
rect 7610 20500 19920 20590
rect 7610 20260 7780 20500
rect 8020 20260 8110 20500
rect 8350 20260 8440 20500
rect 8680 20260 8770 20500
rect 9010 20260 9100 20500
rect 9340 20260 9430 20500
rect 9670 20260 9760 20500
rect 10000 20260 10090 20500
rect 10330 20260 10420 20500
rect 10660 20260 10750 20500
rect 10990 20260 11080 20500
rect 11320 20260 11410 20500
rect 11650 20260 11740 20500
rect 11980 20260 12070 20500
rect 12310 20260 12400 20500
rect 12640 20260 12730 20500
rect 12970 20260 13060 20500
rect 13300 20260 13390 20500
rect 13630 20260 13720 20500
rect 13960 20260 14050 20500
rect 14290 20260 14380 20500
rect 14620 20260 14710 20500
rect 14950 20260 15040 20500
rect 15280 20260 15370 20500
rect 15610 20260 15700 20500
rect 15940 20260 16030 20500
rect 16270 20260 16360 20500
rect 16600 20260 16690 20500
rect 16930 20260 17020 20500
rect 17260 20260 17350 20500
rect 17590 20260 17680 20500
rect 17920 20260 18010 20500
rect 18250 20260 18340 20500
rect 18580 20260 18670 20500
rect 18910 20260 19000 20500
rect 19240 20260 19330 20500
rect 19570 20260 19920 20500
rect 7610 20170 19920 20260
rect 7610 19930 7780 20170
rect 8020 19930 8110 20170
rect 8350 19930 8440 20170
rect 8680 19930 8770 20170
rect 9010 19930 9100 20170
rect 9340 19930 9430 20170
rect 9670 19930 9760 20170
rect 10000 19930 10090 20170
rect 10330 19930 10420 20170
rect 10660 19930 10750 20170
rect 10990 19930 11080 20170
rect 11320 19930 11410 20170
rect 11650 19930 11740 20170
rect 11980 19930 12070 20170
rect 12310 19930 12400 20170
rect 12640 19930 12730 20170
rect 12970 19930 13060 20170
rect 13300 19930 13390 20170
rect 13630 19930 13720 20170
rect 13960 19930 14050 20170
rect 14290 19930 14380 20170
rect 14620 19930 14710 20170
rect 14950 19930 15040 20170
rect 15280 19930 15370 20170
rect 15610 19930 15700 20170
rect 15940 19930 16030 20170
rect 16270 19930 16360 20170
rect 16600 19930 16690 20170
rect 16930 19930 17020 20170
rect 17260 19930 17350 20170
rect 17590 19930 17680 20170
rect 17920 19930 18010 20170
rect 18250 19930 18340 20170
rect 18580 19930 18670 20170
rect 18910 19930 19000 20170
rect 19240 19930 19330 20170
rect 19570 19930 19920 20170
rect 7610 19840 19920 19930
rect 7610 19600 7780 19840
rect 8020 19600 8110 19840
rect 8350 19600 8440 19840
rect 8680 19600 8770 19840
rect 9010 19600 9100 19840
rect 9340 19600 9430 19840
rect 9670 19600 9760 19840
rect 10000 19600 10090 19840
rect 10330 19600 10420 19840
rect 10660 19600 10750 19840
rect 10990 19600 11080 19840
rect 11320 19600 11410 19840
rect 11650 19600 11740 19840
rect 11980 19600 12070 19840
rect 12310 19600 12400 19840
rect 12640 19600 12730 19840
rect 12970 19600 13060 19840
rect 13300 19600 13390 19840
rect 13630 19600 13720 19840
rect 13960 19600 14050 19840
rect 14290 19600 14380 19840
rect 14620 19600 14710 19840
rect 14950 19600 15040 19840
rect 15280 19600 15370 19840
rect 15610 19600 15700 19840
rect 15940 19600 16030 19840
rect 16270 19600 16360 19840
rect 16600 19600 16690 19840
rect 16930 19600 17020 19840
rect 17260 19600 17350 19840
rect 17590 19600 17680 19840
rect 17920 19600 18010 19840
rect 18250 19600 18340 19840
rect 18580 19600 18670 19840
rect 18910 19600 19000 19840
rect 19240 19600 19330 19840
rect 19570 19600 19920 19840
rect 7610 19510 19920 19600
rect 7610 19270 7780 19510
rect 8020 19270 8110 19510
rect 8350 19270 8440 19510
rect 8680 19270 8770 19510
rect 9010 19270 9100 19510
rect 9340 19270 9430 19510
rect 9670 19270 9760 19510
rect 10000 19270 10090 19510
rect 10330 19270 10420 19510
rect 10660 19270 10750 19510
rect 10990 19270 11080 19510
rect 11320 19270 11410 19510
rect 11650 19270 11740 19510
rect 11980 19270 12070 19510
rect 12310 19270 12400 19510
rect 12640 19270 12730 19510
rect 12970 19270 13060 19510
rect 13300 19270 13390 19510
rect 13630 19270 13720 19510
rect 13960 19270 14050 19510
rect 14290 19270 14380 19510
rect 14620 19270 14710 19510
rect 14950 19270 15040 19510
rect 15280 19270 15370 19510
rect 15610 19270 15700 19510
rect 15940 19270 16030 19510
rect 16270 19270 16360 19510
rect 16600 19270 16690 19510
rect 16930 19270 17020 19510
rect 17260 19270 17350 19510
rect 17590 19270 17680 19510
rect 17920 19270 18010 19510
rect 18250 19270 18340 19510
rect 18580 19270 18670 19510
rect 18910 19270 19000 19510
rect 19240 19270 19330 19510
rect 19570 19270 19920 19510
rect 7610 19180 19920 19270
rect 7610 18940 7780 19180
rect 8020 18940 8110 19180
rect 8350 18940 8440 19180
rect 8680 18940 8770 19180
rect 9010 18940 9100 19180
rect 9340 18940 9430 19180
rect 9670 18940 9760 19180
rect 10000 18940 10090 19180
rect 10330 18940 10420 19180
rect 10660 18940 10750 19180
rect 10990 18940 11080 19180
rect 11320 18940 11410 19180
rect 11650 18940 11740 19180
rect 11980 18940 12070 19180
rect 12310 18940 12400 19180
rect 12640 18940 12730 19180
rect 12970 18940 13060 19180
rect 13300 18940 13390 19180
rect 13630 18940 13720 19180
rect 13960 18940 14050 19180
rect 14290 18940 14380 19180
rect 14620 18940 14710 19180
rect 14950 18940 15040 19180
rect 15280 18940 15370 19180
rect 15610 18940 15700 19180
rect 15940 18940 16030 19180
rect 16270 18940 16360 19180
rect 16600 18940 16690 19180
rect 16930 18940 17020 19180
rect 17260 18940 17350 19180
rect 17590 18940 17680 19180
rect 17920 18940 18010 19180
rect 18250 18940 18340 19180
rect 18580 18940 18670 19180
rect 18910 18940 19000 19180
rect 19240 18940 19330 19180
rect 19570 18940 19920 19180
rect 7610 18850 19920 18940
rect 7610 18610 7780 18850
rect 8020 18610 8110 18850
rect 8350 18610 8440 18850
rect 8680 18610 8770 18850
rect 9010 18610 9100 18850
rect 9340 18610 9430 18850
rect 9670 18610 9760 18850
rect 10000 18610 10090 18850
rect 10330 18610 10420 18850
rect 10660 18610 10750 18850
rect 10990 18610 11080 18850
rect 11320 18610 11410 18850
rect 11650 18610 11740 18850
rect 11980 18610 12070 18850
rect 12310 18610 12400 18850
rect 12640 18610 12730 18850
rect 12970 18610 13060 18850
rect 13300 18610 13390 18850
rect 13630 18610 13720 18850
rect 13960 18610 14050 18850
rect 14290 18610 14380 18850
rect 14620 18610 14710 18850
rect 14950 18610 15040 18850
rect 15280 18610 15370 18850
rect 15610 18610 15700 18850
rect 15940 18610 16030 18850
rect 16270 18610 16360 18850
rect 16600 18610 16690 18850
rect 16930 18610 17020 18850
rect 17260 18610 17350 18850
rect 17590 18610 17680 18850
rect 17920 18610 18010 18850
rect 18250 18610 18340 18850
rect 18580 18610 18670 18850
rect 18910 18610 19000 18850
rect 19240 18610 19330 18850
rect 19570 18610 19920 18850
rect 7610 18520 19920 18610
rect 7610 18280 7780 18520
rect 8020 18280 8110 18520
rect 8350 18280 8440 18520
rect 8680 18280 8770 18520
rect 9010 18280 9100 18520
rect 9340 18280 9430 18520
rect 9670 18280 9760 18520
rect 10000 18280 10090 18520
rect 10330 18280 10420 18520
rect 10660 18280 10750 18520
rect 10990 18280 11080 18520
rect 11320 18280 11410 18520
rect 11650 18280 11740 18520
rect 11980 18280 12070 18520
rect 12310 18280 12400 18520
rect 12640 18280 12730 18520
rect 12970 18280 13060 18520
rect 13300 18280 13390 18520
rect 13630 18280 13720 18520
rect 13960 18280 14050 18520
rect 14290 18280 14380 18520
rect 14620 18280 14710 18520
rect 14950 18280 15040 18520
rect 15280 18280 15370 18520
rect 15610 18280 15700 18520
rect 15940 18280 16030 18520
rect 16270 18280 16360 18520
rect 16600 18280 16690 18520
rect 16930 18280 17020 18520
rect 17260 18280 17350 18520
rect 17590 18280 17680 18520
rect 17920 18280 18010 18520
rect 18250 18280 18340 18520
rect 18580 18280 18670 18520
rect 18910 18280 19000 18520
rect 19240 18280 19330 18520
rect 19570 18280 19920 18520
rect 7610 18190 19920 18280
rect 7610 17950 7780 18190
rect 8020 17950 8110 18190
rect 8350 17950 8440 18190
rect 8680 17950 8770 18190
rect 9010 17950 9100 18190
rect 9340 17950 9430 18190
rect 9670 17950 9760 18190
rect 10000 17950 10090 18190
rect 10330 17950 10420 18190
rect 10660 17950 10750 18190
rect 10990 17950 11080 18190
rect 11320 17950 11410 18190
rect 11650 17950 11740 18190
rect 11980 17950 12070 18190
rect 12310 17950 12400 18190
rect 12640 17950 12730 18190
rect 12970 17950 13060 18190
rect 13300 17950 13390 18190
rect 13630 17950 13720 18190
rect 13960 17950 14050 18190
rect 14290 17950 14380 18190
rect 14620 17950 14710 18190
rect 14950 17950 15040 18190
rect 15280 17950 15370 18190
rect 15610 17950 15700 18190
rect 15940 17950 16030 18190
rect 16270 17950 16360 18190
rect 16600 17950 16690 18190
rect 16930 17950 17020 18190
rect 17260 17950 17350 18190
rect 17590 17950 17680 18190
rect 17920 17950 18010 18190
rect 18250 17950 18340 18190
rect 18580 17950 18670 18190
rect 18910 17950 19000 18190
rect 19240 17950 19330 18190
rect 19570 17950 19920 18190
rect 7610 17860 19920 17950
rect 7610 17620 7780 17860
rect 8020 17620 8110 17860
rect 8350 17620 8440 17860
rect 8680 17620 8770 17860
rect 9010 17620 9100 17860
rect 9340 17620 9430 17860
rect 9670 17620 9760 17860
rect 10000 17620 10090 17860
rect 10330 17620 10420 17860
rect 10660 17620 10750 17860
rect 10990 17620 11080 17860
rect 11320 17620 11410 17860
rect 11650 17620 11740 17860
rect 11980 17620 12070 17860
rect 12310 17620 12400 17860
rect 12640 17620 12730 17860
rect 12970 17620 13060 17860
rect 13300 17620 13390 17860
rect 13630 17620 13720 17860
rect 13960 17620 14050 17860
rect 14290 17620 14380 17860
rect 14620 17620 14710 17860
rect 14950 17620 15040 17860
rect 15280 17620 15370 17860
rect 15610 17620 15700 17860
rect 15940 17620 16030 17860
rect 16270 17620 16360 17860
rect 16600 17620 16690 17860
rect 16930 17620 17020 17860
rect 17260 17620 17350 17860
rect 17590 17620 17680 17860
rect 17920 17620 18010 17860
rect 18250 17620 18340 17860
rect 18580 17620 18670 17860
rect 18910 17620 19000 17860
rect 19240 17620 19330 17860
rect 19570 17620 19920 17860
rect 7610 17530 19920 17620
rect 7610 17290 7780 17530
rect 8020 17290 8110 17530
rect 8350 17290 8440 17530
rect 8680 17290 8770 17530
rect 9010 17290 9100 17530
rect 9340 17290 9430 17530
rect 9670 17290 9760 17530
rect 10000 17290 10090 17530
rect 10330 17290 10420 17530
rect 10660 17290 10750 17530
rect 10990 17290 11080 17530
rect 11320 17290 11410 17530
rect 11650 17290 11740 17530
rect 11980 17290 12070 17530
rect 12310 17290 12400 17530
rect 12640 17290 12730 17530
rect 12970 17290 13060 17530
rect 13300 17290 13390 17530
rect 13630 17290 13720 17530
rect 13960 17290 14050 17530
rect 14290 17290 14380 17530
rect 14620 17290 14710 17530
rect 14950 17290 15040 17530
rect 15280 17290 15370 17530
rect 15610 17290 15700 17530
rect 15940 17290 16030 17530
rect 16270 17290 16360 17530
rect 16600 17290 16690 17530
rect 16930 17290 17020 17530
rect 17260 17290 17350 17530
rect 17590 17290 17680 17530
rect 17920 17290 18010 17530
rect 18250 17290 18340 17530
rect 18580 17290 18670 17530
rect 18910 17290 19000 17530
rect 19240 17290 19330 17530
rect 19570 17290 19920 17530
rect 7610 17200 19920 17290
rect 7610 16960 7780 17200
rect 8020 16960 8110 17200
rect 8350 16960 8440 17200
rect 8680 16960 8770 17200
rect 9010 16960 9100 17200
rect 9340 16960 9430 17200
rect 9670 16960 9760 17200
rect 10000 16960 10090 17200
rect 10330 16960 10420 17200
rect 10660 16960 10750 17200
rect 10990 16960 11080 17200
rect 11320 16960 11410 17200
rect 11650 16960 11740 17200
rect 11980 16960 12070 17200
rect 12310 16960 12400 17200
rect 12640 16960 12730 17200
rect 12970 16960 13060 17200
rect 13300 16960 13390 17200
rect 13630 16960 13720 17200
rect 13960 16960 14050 17200
rect 14290 16960 14380 17200
rect 14620 16960 14710 17200
rect 14950 16960 15040 17200
rect 15280 16960 15370 17200
rect 15610 16960 15700 17200
rect 15940 16960 16030 17200
rect 16270 16960 16360 17200
rect 16600 16960 16690 17200
rect 16930 16960 17020 17200
rect 17260 16960 17350 17200
rect 17590 16960 17680 17200
rect 17920 16960 18010 17200
rect 18250 16960 18340 17200
rect 18580 16960 18670 17200
rect 18910 16960 19000 17200
rect 19240 16960 19330 17200
rect 19570 16960 19920 17200
rect 7610 16870 19920 16960
rect 7610 16630 7780 16870
rect 8020 16630 8110 16870
rect 8350 16630 8440 16870
rect 8680 16630 8770 16870
rect 9010 16630 9100 16870
rect 9340 16630 9430 16870
rect 9670 16630 9760 16870
rect 10000 16630 10090 16870
rect 10330 16630 10420 16870
rect 10660 16630 10750 16870
rect 10990 16630 11080 16870
rect 11320 16630 11410 16870
rect 11650 16630 11740 16870
rect 11980 16630 12070 16870
rect 12310 16630 12400 16870
rect 12640 16630 12730 16870
rect 12970 16630 13060 16870
rect 13300 16630 13390 16870
rect 13630 16630 13720 16870
rect 13960 16630 14050 16870
rect 14290 16630 14380 16870
rect 14620 16630 14710 16870
rect 14950 16630 15040 16870
rect 15280 16630 15370 16870
rect 15610 16630 15700 16870
rect 15940 16630 16030 16870
rect 16270 16630 16360 16870
rect 16600 16630 16690 16870
rect 16930 16630 17020 16870
rect 17260 16630 17350 16870
rect 17590 16630 17680 16870
rect 17920 16630 18010 16870
rect 18250 16630 18340 16870
rect 18580 16630 18670 16870
rect 18910 16630 19000 16870
rect 19240 16630 19330 16870
rect 19570 16630 19920 16870
rect 7610 16540 19920 16630
rect 7610 16300 7780 16540
rect 8020 16300 8110 16540
rect 8350 16300 8440 16540
rect 8680 16300 8770 16540
rect 9010 16300 9100 16540
rect 9340 16300 9430 16540
rect 9670 16300 9760 16540
rect 10000 16300 10090 16540
rect 10330 16300 10420 16540
rect 10660 16300 10750 16540
rect 10990 16300 11080 16540
rect 11320 16300 11410 16540
rect 11650 16300 11740 16540
rect 11980 16300 12070 16540
rect 12310 16300 12400 16540
rect 12640 16300 12730 16540
rect 12970 16300 13060 16540
rect 13300 16300 13390 16540
rect 13630 16300 13720 16540
rect 13960 16300 14050 16540
rect 14290 16300 14380 16540
rect 14620 16300 14710 16540
rect 14950 16300 15040 16540
rect 15280 16300 15370 16540
rect 15610 16300 15700 16540
rect 15940 16300 16030 16540
rect 16270 16300 16360 16540
rect 16600 16300 16690 16540
rect 16930 16300 17020 16540
rect 17260 16300 17350 16540
rect 17590 16300 17680 16540
rect 17920 16300 18010 16540
rect 18250 16300 18340 16540
rect 18580 16300 18670 16540
rect 18910 16300 19000 16540
rect 19240 16300 19330 16540
rect 19570 16300 19920 16540
rect 7610 16210 19920 16300
rect 7610 15970 7780 16210
rect 8020 15970 8110 16210
rect 8350 15970 8440 16210
rect 8680 15970 8770 16210
rect 9010 15970 9100 16210
rect 9340 15970 9430 16210
rect 9670 15970 9760 16210
rect 10000 15970 10090 16210
rect 10330 15970 10420 16210
rect 10660 15970 10750 16210
rect 10990 15970 11080 16210
rect 11320 15970 11410 16210
rect 11650 15970 11740 16210
rect 11980 15970 12070 16210
rect 12310 15970 12400 16210
rect 12640 15970 12730 16210
rect 12970 15970 13060 16210
rect 13300 15970 13390 16210
rect 13630 15970 13720 16210
rect 13960 15970 14050 16210
rect 14290 15970 14380 16210
rect 14620 15970 14710 16210
rect 14950 15970 15040 16210
rect 15280 15970 15370 16210
rect 15610 15970 15700 16210
rect 15940 15970 16030 16210
rect 16270 15970 16360 16210
rect 16600 15970 16690 16210
rect 16930 15970 17020 16210
rect 17260 15970 17350 16210
rect 17590 15970 17680 16210
rect 17920 15970 18010 16210
rect 18250 15970 18340 16210
rect 18580 15970 18670 16210
rect 18910 15970 19000 16210
rect 19240 15970 19330 16210
rect 19570 15970 19920 16210
rect 7610 15880 19920 15970
rect 7610 15640 7780 15880
rect 8020 15640 8110 15880
rect 8350 15640 8440 15880
rect 8680 15640 8770 15880
rect 9010 15640 9100 15880
rect 9340 15640 9430 15880
rect 9670 15640 9760 15880
rect 10000 15640 10090 15880
rect 10330 15640 10420 15880
rect 10660 15640 10750 15880
rect 10990 15640 11080 15880
rect 11320 15640 11410 15880
rect 11650 15640 11740 15880
rect 11980 15640 12070 15880
rect 12310 15640 12400 15880
rect 12640 15640 12730 15880
rect 12970 15640 13060 15880
rect 13300 15640 13390 15880
rect 13630 15640 13720 15880
rect 13960 15640 14050 15880
rect 14290 15640 14380 15880
rect 14620 15640 14710 15880
rect 14950 15640 15040 15880
rect 15280 15640 15370 15880
rect 15610 15640 15700 15880
rect 15940 15640 16030 15880
rect 16270 15640 16360 15880
rect 16600 15640 16690 15880
rect 16930 15640 17020 15880
rect 17260 15640 17350 15880
rect 17590 15640 17680 15880
rect 17920 15640 18010 15880
rect 18250 15640 18340 15880
rect 18580 15640 18670 15880
rect 18910 15640 19000 15880
rect 19240 15640 19330 15880
rect 19570 15640 19920 15880
rect 7610 15550 19920 15640
rect 7610 15310 7780 15550
rect 8020 15310 8110 15550
rect 8350 15310 8440 15550
rect 8680 15310 8770 15550
rect 9010 15310 9100 15550
rect 9340 15310 9430 15550
rect 9670 15310 9760 15550
rect 10000 15310 10090 15550
rect 10330 15310 10420 15550
rect 10660 15310 10750 15550
rect 10990 15310 11080 15550
rect 11320 15310 11410 15550
rect 11650 15310 11740 15550
rect 11980 15310 12070 15550
rect 12310 15310 12400 15550
rect 12640 15310 12730 15550
rect 12970 15310 13060 15550
rect 13300 15310 13390 15550
rect 13630 15310 13720 15550
rect 13960 15310 14050 15550
rect 14290 15310 14380 15550
rect 14620 15310 14710 15550
rect 14950 15310 15040 15550
rect 15280 15310 15370 15550
rect 15610 15310 15700 15550
rect 15940 15310 16030 15550
rect 16270 15310 16360 15550
rect 16600 15310 16690 15550
rect 16930 15310 17020 15550
rect 17260 15310 17350 15550
rect 17590 15310 17680 15550
rect 17920 15310 18010 15550
rect 18250 15310 18340 15550
rect 18580 15310 18670 15550
rect 18910 15310 19000 15550
rect 19240 15310 19330 15550
rect 19570 15310 19920 15550
rect 7610 15220 19920 15310
rect 7610 14980 7780 15220
rect 8020 14980 8110 15220
rect 8350 14980 8440 15220
rect 8680 14980 8770 15220
rect 9010 14980 9100 15220
rect 9340 14980 9430 15220
rect 9670 14980 9760 15220
rect 10000 14980 10090 15220
rect 10330 14980 10420 15220
rect 10660 14980 10750 15220
rect 10990 14980 11080 15220
rect 11320 14980 11410 15220
rect 11650 14980 11740 15220
rect 11980 14980 12070 15220
rect 12310 14980 12400 15220
rect 12640 14980 12730 15220
rect 12970 14980 13060 15220
rect 13300 14980 13390 15220
rect 13630 14980 13720 15220
rect 13960 14980 14050 15220
rect 14290 14980 14380 15220
rect 14620 14980 14710 15220
rect 14950 14980 15040 15220
rect 15280 14980 15370 15220
rect 15610 14980 15700 15220
rect 15940 14980 16030 15220
rect 16270 14980 16360 15220
rect 16600 14980 16690 15220
rect 16930 14980 17020 15220
rect 17260 14980 17350 15220
rect 17590 14980 17680 15220
rect 17920 14980 18010 15220
rect 18250 14980 18340 15220
rect 18580 14980 18670 15220
rect 18910 14980 19000 15220
rect 19240 14980 19330 15220
rect 19570 14980 19920 15220
rect 7610 14890 19920 14980
rect 7610 14650 7780 14890
rect 8020 14650 8110 14890
rect 8350 14650 8440 14890
rect 8680 14650 8770 14890
rect 9010 14650 9100 14890
rect 9340 14650 9430 14890
rect 9670 14650 9760 14890
rect 10000 14650 10090 14890
rect 10330 14650 10420 14890
rect 10660 14650 10750 14890
rect 10990 14650 11080 14890
rect 11320 14650 11410 14890
rect 11650 14650 11740 14890
rect 11980 14650 12070 14890
rect 12310 14650 12400 14890
rect 12640 14650 12730 14890
rect 12970 14650 13060 14890
rect 13300 14650 13390 14890
rect 13630 14650 13720 14890
rect 13960 14650 14050 14890
rect 14290 14650 14380 14890
rect 14620 14650 14710 14890
rect 14950 14650 15040 14890
rect 15280 14650 15370 14890
rect 15610 14650 15700 14890
rect 15940 14650 16030 14890
rect 16270 14650 16360 14890
rect 16600 14650 16690 14890
rect 16930 14650 17020 14890
rect 17260 14650 17350 14890
rect 17590 14650 17680 14890
rect 17920 14650 18010 14890
rect 18250 14650 18340 14890
rect 18580 14650 18670 14890
rect 18910 14650 19000 14890
rect 19240 14650 19330 14890
rect 19570 14650 19920 14890
rect 7610 14560 19920 14650
rect 7610 14320 7780 14560
rect 8020 14320 8110 14560
rect 8350 14320 8440 14560
rect 8680 14320 8770 14560
rect 9010 14320 9100 14560
rect 9340 14320 9430 14560
rect 9670 14320 9760 14560
rect 10000 14320 10090 14560
rect 10330 14320 10420 14560
rect 10660 14320 10750 14560
rect 10990 14320 11080 14560
rect 11320 14320 11410 14560
rect 11650 14320 11740 14560
rect 11980 14320 12070 14560
rect 12310 14320 12400 14560
rect 12640 14320 12730 14560
rect 12970 14320 13060 14560
rect 13300 14320 13390 14560
rect 13630 14320 13720 14560
rect 13960 14320 14050 14560
rect 14290 14320 14380 14560
rect 14620 14320 14710 14560
rect 14950 14320 15040 14560
rect 15280 14320 15370 14560
rect 15610 14320 15700 14560
rect 15940 14320 16030 14560
rect 16270 14320 16360 14560
rect 16600 14320 16690 14560
rect 16930 14320 17020 14560
rect 17260 14320 17350 14560
rect 17590 14320 17680 14560
rect 17920 14320 18010 14560
rect 18250 14320 18340 14560
rect 18580 14320 18670 14560
rect 18910 14320 19000 14560
rect 19240 14320 19330 14560
rect 19570 14320 19920 14560
rect 7610 14230 19920 14320
rect 7610 13990 7780 14230
rect 8020 13990 8110 14230
rect 8350 13990 8440 14230
rect 8680 13990 8770 14230
rect 9010 13990 9100 14230
rect 9340 13990 9430 14230
rect 9670 13990 9760 14230
rect 10000 13990 10090 14230
rect 10330 13990 10420 14230
rect 10660 13990 10750 14230
rect 10990 13990 11080 14230
rect 11320 13990 11410 14230
rect 11650 13990 11740 14230
rect 11980 13990 12070 14230
rect 12310 13990 12400 14230
rect 12640 13990 12730 14230
rect 12970 13990 13060 14230
rect 13300 13990 13390 14230
rect 13630 13990 13720 14230
rect 13960 13990 14050 14230
rect 14290 13990 14380 14230
rect 14620 13990 14710 14230
rect 14950 13990 15040 14230
rect 15280 13990 15370 14230
rect 15610 13990 15700 14230
rect 15940 13990 16030 14230
rect 16270 13990 16360 14230
rect 16600 13990 16690 14230
rect 16930 13990 17020 14230
rect 17260 13990 17350 14230
rect 17590 13990 17680 14230
rect 17920 13990 18010 14230
rect 18250 13990 18340 14230
rect 18580 13990 18670 14230
rect 18910 13990 19000 14230
rect 19240 13990 19330 14230
rect 19570 13990 19920 14230
rect 7610 13900 19920 13990
rect 7610 13660 7780 13900
rect 8020 13660 8110 13900
rect 8350 13660 8440 13900
rect 8680 13660 8770 13900
rect 9010 13660 9100 13900
rect 9340 13660 9430 13900
rect 9670 13660 9760 13900
rect 10000 13660 10090 13900
rect 10330 13660 10420 13900
rect 10660 13660 10750 13900
rect 10990 13660 11080 13900
rect 11320 13660 11410 13900
rect 11650 13660 11740 13900
rect 11980 13660 12070 13900
rect 12310 13660 12400 13900
rect 12640 13660 12730 13900
rect 12970 13660 13060 13900
rect 13300 13660 13390 13900
rect 13630 13660 13720 13900
rect 13960 13660 14050 13900
rect 14290 13660 14380 13900
rect 14620 13660 14710 13900
rect 14950 13660 15040 13900
rect 15280 13660 15370 13900
rect 15610 13660 15700 13900
rect 15940 13660 16030 13900
rect 16270 13660 16360 13900
rect 16600 13660 16690 13900
rect 16930 13660 17020 13900
rect 17260 13660 17350 13900
rect 17590 13660 17680 13900
rect 17920 13660 18010 13900
rect 18250 13660 18340 13900
rect 18580 13660 18670 13900
rect 18910 13660 19000 13900
rect 19240 13660 19330 13900
rect 19570 13660 19920 13900
rect 7610 13570 19920 13660
rect 7610 13330 7780 13570
rect 8020 13330 8110 13570
rect 8350 13330 8440 13570
rect 8680 13330 8770 13570
rect 9010 13330 9100 13570
rect 9340 13330 9430 13570
rect 9670 13330 9760 13570
rect 10000 13330 10090 13570
rect 10330 13330 10420 13570
rect 10660 13330 10750 13570
rect 10990 13330 11080 13570
rect 11320 13330 11410 13570
rect 11650 13330 11740 13570
rect 11980 13330 12070 13570
rect 12310 13330 12400 13570
rect 12640 13330 12730 13570
rect 12970 13330 13060 13570
rect 13300 13330 13390 13570
rect 13630 13330 13720 13570
rect 13960 13330 14050 13570
rect 14290 13330 14380 13570
rect 14620 13330 14710 13570
rect 14950 13330 15040 13570
rect 15280 13330 15370 13570
rect 15610 13330 15700 13570
rect 15940 13330 16030 13570
rect 16270 13330 16360 13570
rect 16600 13330 16690 13570
rect 16930 13330 17020 13570
rect 17260 13330 17350 13570
rect 17590 13330 17680 13570
rect 17920 13330 18010 13570
rect 18250 13330 18340 13570
rect 18580 13330 18670 13570
rect 18910 13330 19000 13570
rect 19240 13330 19330 13570
rect 19570 13330 19920 13570
rect 7610 13240 19920 13330
rect 7610 13000 7780 13240
rect 8020 13000 8110 13240
rect 8350 13000 8440 13240
rect 8680 13000 8770 13240
rect 9010 13000 9100 13240
rect 9340 13000 9430 13240
rect 9670 13000 9760 13240
rect 10000 13000 10090 13240
rect 10330 13000 10420 13240
rect 10660 13000 10750 13240
rect 10990 13000 11080 13240
rect 11320 13000 11410 13240
rect 11650 13000 11740 13240
rect 11980 13000 12070 13240
rect 12310 13000 12400 13240
rect 12640 13000 12730 13240
rect 12970 13000 13060 13240
rect 13300 13000 13390 13240
rect 13630 13000 13720 13240
rect 13960 13000 14050 13240
rect 14290 13000 14380 13240
rect 14620 13000 14710 13240
rect 14950 13000 15040 13240
rect 15280 13000 15370 13240
rect 15610 13000 15700 13240
rect 15940 13000 16030 13240
rect 16270 13000 16360 13240
rect 16600 13000 16690 13240
rect 16930 13000 17020 13240
rect 17260 13000 17350 13240
rect 17590 13000 17680 13240
rect 17920 13000 18010 13240
rect 18250 13000 18340 13240
rect 18580 13000 18670 13240
rect 18910 13000 19000 13240
rect 19240 13000 19330 13240
rect 19570 13000 19920 13240
rect 7610 12910 19920 13000
rect 7610 12670 7780 12910
rect 8020 12670 8110 12910
rect 8350 12670 8440 12910
rect 8680 12670 8770 12910
rect 9010 12670 9100 12910
rect 9340 12670 9430 12910
rect 9670 12670 9760 12910
rect 10000 12670 10090 12910
rect 10330 12670 10420 12910
rect 10660 12670 10750 12910
rect 10990 12670 11080 12910
rect 11320 12670 11410 12910
rect 11650 12670 11740 12910
rect 11980 12670 12070 12910
rect 12310 12670 12400 12910
rect 12640 12670 12730 12910
rect 12970 12670 13060 12910
rect 13300 12670 13390 12910
rect 13630 12670 13720 12910
rect 13960 12670 14050 12910
rect 14290 12670 14380 12910
rect 14620 12670 14710 12910
rect 14950 12670 15040 12910
rect 15280 12670 15370 12910
rect 15610 12670 15700 12910
rect 15940 12670 16030 12910
rect 16270 12670 16360 12910
rect 16600 12670 16690 12910
rect 16930 12670 17020 12910
rect 17260 12670 17350 12910
rect 17590 12670 17680 12910
rect 17920 12670 18010 12910
rect 18250 12670 18340 12910
rect 18580 12670 18670 12910
rect 18910 12670 19000 12910
rect 19240 12670 19330 12910
rect 19570 12670 19920 12910
rect 7610 12580 19920 12670
rect 7610 12340 7780 12580
rect 8020 12340 8110 12580
rect 8350 12340 8440 12580
rect 8680 12340 8770 12580
rect 9010 12340 9100 12580
rect 9340 12340 9430 12580
rect 9670 12340 9760 12580
rect 10000 12340 10090 12580
rect 10330 12340 10420 12580
rect 10660 12340 10750 12580
rect 10990 12340 11080 12580
rect 11320 12340 11410 12580
rect 11650 12340 11740 12580
rect 11980 12340 12070 12580
rect 12310 12340 12400 12580
rect 12640 12340 12730 12580
rect 12970 12340 13060 12580
rect 13300 12340 13390 12580
rect 13630 12340 13720 12580
rect 13960 12340 14050 12580
rect 14290 12340 14380 12580
rect 14620 12340 14710 12580
rect 14950 12340 15040 12580
rect 15280 12340 15370 12580
rect 15610 12340 15700 12580
rect 15940 12340 16030 12580
rect 16270 12340 16360 12580
rect 16600 12340 16690 12580
rect 16930 12340 17020 12580
rect 17260 12340 17350 12580
rect 17590 12340 17680 12580
rect 17920 12340 18010 12580
rect 18250 12340 18340 12580
rect 18580 12340 18670 12580
rect 18910 12340 19000 12580
rect 19240 12340 19330 12580
rect 19570 12340 19920 12580
rect 7610 12250 19920 12340
rect 7610 12010 7780 12250
rect 8020 12010 8110 12250
rect 8350 12010 8440 12250
rect 8680 12010 8770 12250
rect 9010 12010 9100 12250
rect 9340 12010 9430 12250
rect 9670 12010 9760 12250
rect 10000 12010 10090 12250
rect 10330 12010 10420 12250
rect 10660 12010 10750 12250
rect 10990 12010 11080 12250
rect 11320 12010 11410 12250
rect 11650 12010 11740 12250
rect 11980 12010 12070 12250
rect 12310 12010 12400 12250
rect 12640 12010 12730 12250
rect 12970 12010 13060 12250
rect 13300 12010 13390 12250
rect 13630 12010 13720 12250
rect 13960 12010 14050 12250
rect 14290 12010 14380 12250
rect 14620 12010 14710 12250
rect 14950 12010 15040 12250
rect 15280 12010 15370 12250
rect 15610 12010 15700 12250
rect 15940 12010 16030 12250
rect 16270 12010 16360 12250
rect 16600 12010 16690 12250
rect 16930 12010 17020 12250
rect 17260 12010 17350 12250
rect 17590 12010 17680 12250
rect 17920 12010 18010 12250
rect 18250 12010 18340 12250
rect 18580 12010 18670 12250
rect 18910 12010 19000 12250
rect 19240 12010 19330 12250
rect 19570 12010 19920 12250
rect 7610 11920 19920 12010
rect 7610 11680 7780 11920
rect 8020 11680 8110 11920
rect 8350 11680 8440 11920
rect 8680 11680 8770 11920
rect 9010 11680 9100 11920
rect 9340 11680 9430 11920
rect 9670 11680 9760 11920
rect 10000 11680 10090 11920
rect 10330 11680 10420 11920
rect 10660 11680 10750 11920
rect 10990 11680 11080 11920
rect 11320 11680 11410 11920
rect 11650 11680 11740 11920
rect 11980 11680 12070 11920
rect 12310 11680 12400 11920
rect 12640 11680 12730 11920
rect 12970 11680 13060 11920
rect 13300 11680 13390 11920
rect 13630 11680 13720 11920
rect 13960 11680 14050 11920
rect 14290 11680 14380 11920
rect 14620 11680 14710 11920
rect 14950 11680 15040 11920
rect 15280 11680 15370 11920
rect 15610 11680 15700 11920
rect 15940 11680 16030 11920
rect 16270 11680 16360 11920
rect 16600 11680 16690 11920
rect 16930 11680 17020 11920
rect 17260 11680 17350 11920
rect 17590 11680 17680 11920
rect 17920 11680 18010 11920
rect 18250 11680 18340 11920
rect 18580 11680 18670 11920
rect 18910 11680 19000 11920
rect 19240 11680 19330 11920
rect 19570 11680 19920 11920
rect 7610 11590 19920 11680
rect 7610 11350 7780 11590
rect 8020 11350 8110 11590
rect 8350 11350 8440 11590
rect 8680 11350 8770 11590
rect 9010 11350 9100 11590
rect 9340 11350 9430 11590
rect 9670 11350 9760 11590
rect 10000 11350 10090 11590
rect 10330 11350 10420 11590
rect 10660 11350 10750 11590
rect 10990 11350 11080 11590
rect 11320 11350 11410 11590
rect 11650 11350 11740 11590
rect 11980 11350 12070 11590
rect 12310 11350 12400 11590
rect 12640 11350 12730 11590
rect 12970 11350 13060 11590
rect 13300 11350 13390 11590
rect 13630 11350 13720 11590
rect 13960 11350 14050 11590
rect 14290 11350 14380 11590
rect 14620 11350 14710 11590
rect 14950 11350 15040 11590
rect 15280 11350 15370 11590
rect 15610 11350 15700 11590
rect 15940 11350 16030 11590
rect 16270 11350 16360 11590
rect 16600 11350 16690 11590
rect 16930 11350 17020 11590
rect 17260 11350 17350 11590
rect 17590 11350 17680 11590
rect 17920 11350 18010 11590
rect 18250 11350 18340 11590
rect 18580 11350 18670 11590
rect 18910 11350 19000 11590
rect 19240 11350 19330 11590
rect 19570 11350 19920 11590
rect 7610 11260 19920 11350
rect 7610 11020 7780 11260
rect 8020 11020 8110 11260
rect 8350 11020 8440 11260
rect 8680 11020 8770 11260
rect 9010 11020 9100 11260
rect 9340 11020 9430 11260
rect 9670 11020 9760 11260
rect 10000 11020 10090 11260
rect 10330 11020 10420 11260
rect 10660 11020 10750 11260
rect 10990 11020 11080 11260
rect 11320 11020 11410 11260
rect 11650 11020 11740 11260
rect 11980 11020 12070 11260
rect 12310 11020 12400 11260
rect 12640 11020 12730 11260
rect 12970 11020 13060 11260
rect 13300 11020 13390 11260
rect 13630 11020 13720 11260
rect 13960 11020 14050 11260
rect 14290 11020 14380 11260
rect 14620 11020 14710 11260
rect 14950 11020 15040 11260
rect 15280 11020 15370 11260
rect 15610 11020 15700 11260
rect 15940 11020 16030 11260
rect 16270 11020 16360 11260
rect 16600 11020 16690 11260
rect 16930 11020 17020 11260
rect 17260 11020 17350 11260
rect 17590 11020 17680 11260
rect 17920 11020 18010 11260
rect 18250 11020 18340 11260
rect 18580 11020 18670 11260
rect 18910 11020 19000 11260
rect 19240 11020 19330 11260
rect 19570 11020 19920 11260
rect 7610 10930 19920 11020
rect 7610 10690 7780 10930
rect 8020 10690 8110 10930
rect 8350 10690 8440 10930
rect 8680 10690 8770 10930
rect 9010 10690 9100 10930
rect 9340 10690 9430 10930
rect 9670 10690 9760 10930
rect 10000 10690 10090 10930
rect 10330 10690 10420 10930
rect 10660 10690 10750 10930
rect 10990 10690 11080 10930
rect 11320 10690 11410 10930
rect 11650 10690 11740 10930
rect 11980 10690 12070 10930
rect 12310 10690 12400 10930
rect 12640 10690 12730 10930
rect 12970 10690 13060 10930
rect 13300 10690 13390 10930
rect 13630 10690 13720 10930
rect 13960 10690 14050 10930
rect 14290 10690 14380 10930
rect 14620 10690 14710 10930
rect 14950 10690 15040 10930
rect 15280 10690 15370 10930
rect 15610 10690 15700 10930
rect 15940 10690 16030 10930
rect 16270 10690 16360 10930
rect 16600 10690 16690 10930
rect 16930 10690 17020 10930
rect 17260 10690 17350 10930
rect 17590 10690 17680 10930
rect 17920 10690 18010 10930
rect 18250 10690 18340 10930
rect 18580 10690 18670 10930
rect 18910 10690 19000 10930
rect 19240 10690 19330 10930
rect 19570 10690 19920 10930
rect 7610 10600 19920 10690
rect 7610 10360 7780 10600
rect 8020 10360 8110 10600
rect 8350 10360 8440 10600
rect 8680 10360 8770 10600
rect 9010 10360 9100 10600
rect 9340 10360 9430 10600
rect 9670 10360 9760 10600
rect 10000 10360 10090 10600
rect 10330 10360 10420 10600
rect 10660 10360 10750 10600
rect 10990 10360 11080 10600
rect 11320 10360 11410 10600
rect 11650 10360 11740 10600
rect 11980 10360 12070 10600
rect 12310 10360 12400 10600
rect 12640 10360 12730 10600
rect 12970 10360 13060 10600
rect 13300 10360 13390 10600
rect 13630 10360 13720 10600
rect 13960 10360 14050 10600
rect 14290 10360 14380 10600
rect 14620 10360 14710 10600
rect 14950 10360 15040 10600
rect 15280 10360 15370 10600
rect 15610 10360 15700 10600
rect 15940 10360 16030 10600
rect 16270 10360 16360 10600
rect 16600 10360 16690 10600
rect 16930 10360 17020 10600
rect 17260 10360 17350 10600
rect 17590 10360 17680 10600
rect 17920 10360 18010 10600
rect 18250 10360 18340 10600
rect 18580 10360 18670 10600
rect 18910 10360 19000 10600
rect 19240 10360 19330 10600
rect 19570 10360 19920 10600
rect 7610 10270 19920 10360
rect 7610 10030 7780 10270
rect 8020 10030 8110 10270
rect 8350 10030 8440 10270
rect 8680 10030 8770 10270
rect 9010 10030 9100 10270
rect 9340 10030 9430 10270
rect 9670 10030 9760 10270
rect 10000 10030 10090 10270
rect 10330 10030 10420 10270
rect 10660 10030 10750 10270
rect 10990 10030 11080 10270
rect 11320 10030 11410 10270
rect 11650 10030 11740 10270
rect 11980 10030 12070 10270
rect 12310 10030 12400 10270
rect 12640 10030 12730 10270
rect 12970 10030 13060 10270
rect 13300 10030 13390 10270
rect 13630 10030 13720 10270
rect 13960 10030 14050 10270
rect 14290 10030 14380 10270
rect 14620 10030 14710 10270
rect 14950 10030 15040 10270
rect 15280 10030 15370 10270
rect 15610 10030 15700 10270
rect 15940 10030 16030 10270
rect 16270 10030 16360 10270
rect 16600 10030 16690 10270
rect 16930 10030 17020 10270
rect 17260 10030 17350 10270
rect 17590 10030 17680 10270
rect 17920 10030 18010 10270
rect 18250 10030 18340 10270
rect 18580 10030 18670 10270
rect 18910 10030 19000 10270
rect 19240 10030 19330 10270
rect 19570 10030 19920 10270
rect 7610 9940 19920 10030
rect 7610 9700 7780 9940
rect 8020 9700 8110 9940
rect 8350 9700 8440 9940
rect 8680 9700 8770 9940
rect 9010 9700 9100 9940
rect 9340 9700 9430 9940
rect 9670 9700 9760 9940
rect 10000 9700 10090 9940
rect 10330 9700 10420 9940
rect 10660 9700 10750 9940
rect 10990 9700 11080 9940
rect 11320 9700 11410 9940
rect 11650 9700 11740 9940
rect 11980 9700 12070 9940
rect 12310 9700 12400 9940
rect 12640 9700 12730 9940
rect 12970 9700 13060 9940
rect 13300 9700 13390 9940
rect 13630 9700 13720 9940
rect 13960 9700 14050 9940
rect 14290 9700 14380 9940
rect 14620 9700 14710 9940
rect 14950 9700 15040 9940
rect 15280 9700 15370 9940
rect 15610 9700 15700 9940
rect 15940 9700 16030 9940
rect 16270 9700 16360 9940
rect 16600 9700 16690 9940
rect 16930 9700 17020 9940
rect 17260 9700 17350 9940
rect 17590 9700 17680 9940
rect 17920 9700 18010 9940
rect 18250 9700 18340 9940
rect 18580 9700 18670 9940
rect 18910 9700 19000 9940
rect 19240 9700 19330 9940
rect 19570 9700 19920 9940
rect 7610 9610 19920 9700
rect 7610 9370 7780 9610
rect 8020 9370 8110 9610
rect 8350 9370 8440 9610
rect 8680 9370 8770 9610
rect 9010 9370 9100 9610
rect 9340 9370 9430 9610
rect 9670 9370 9760 9610
rect 10000 9370 10090 9610
rect 10330 9370 10420 9610
rect 10660 9370 10750 9610
rect 10990 9370 11080 9610
rect 11320 9370 11410 9610
rect 11650 9370 11740 9610
rect 11980 9370 12070 9610
rect 12310 9370 12400 9610
rect 12640 9370 12730 9610
rect 12970 9370 13060 9610
rect 13300 9370 13390 9610
rect 13630 9370 13720 9610
rect 13960 9370 14050 9610
rect 14290 9370 14380 9610
rect 14620 9370 14710 9610
rect 14950 9370 15040 9610
rect 15280 9370 15370 9610
rect 15610 9370 15700 9610
rect 15940 9370 16030 9610
rect 16270 9370 16360 9610
rect 16600 9370 16690 9610
rect 16930 9370 17020 9610
rect 17260 9370 17350 9610
rect 17590 9370 17680 9610
rect 17920 9370 18010 9610
rect 18250 9370 18340 9610
rect 18580 9370 18670 9610
rect 18910 9370 19000 9610
rect 19240 9370 19330 9610
rect 19570 9370 19920 9610
rect 7610 9280 19920 9370
rect 7610 9040 7780 9280
rect 8020 9040 8110 9280
rect 8350 9040 8440 9280
rect 8680 9040 8770 9280
rect 9010 9040 9100 9280
rect 9340 9040 9430 9280
rect 9670 9040 9760 9280
rect 10000 9040 10090 9280
rect 10330 9040 10420 9280
rect 10660 9040 10750 9280
rect 10990 9040 11080 9280
rect 11320 9040 11410 9280
rect 11650 9040 11740 9280
rect 11980 9040 12070 9280
rect 12310 9040 12400 9280
rect 12640 9040 12730 9280
rect 12970 9040 13060 9280
rect 13300 9040 13390 9280
rect 13630 9040 13720 9280
rect 13960 9040 14050 9280
rect 14290 9040 14380 9280
rect 14620 9040 14710 9280
rect 14950 9040 15040 9280
rect 15280 9040 15370 9280
rect 15610 9040 15700 9280
rect 15940 9040 16030 9280
rect 16270 9040 16360 9280
rect 16600 9040 16690 9280
rect 16930 9040 17020 9280
rect 17260 9040 17350 9280
rect 17590 9040 17680 9280
rect 17920 9040 18010 9280
rect 18250 9040 18340 9280
rect 18580 9040 18670 9280
rect 18910 9040 19000 9280
rect 19240 9040 19330 9280
rect 19570 9040 19920 9280
rect 7610 8690 19920 9040
rect -6530 7270 29270 8130
rect -6530 7100 23510 7270
rect -6530 -2160 -2530 7100
rect 1540 6910 3140 7100
rect 1540 6670 1720 6910
rect 1960 6670 2050 6910
rect 2290 6670 2390 6910
rect 2630 6670 2720 6910
rect 2960 6670 3140 6910
rect 11760 6940 13360 7100
rect 23460 7030 23510 7100
rect 23880 7100 25910 7270
rect 23880 7030 23940 7100
rect 23460 7000 23940 7030
rect 25860 7030 25910 7100
rect 26280 7100 29270 7270
rect 26280 7030 26340 7100
rect 25860 7000 26340 7030
rect 11760 6700 11940 6940
rect 12180 6700 12270 6940
rect 12510 6700 12610 6940
rect 12850 6700 12940 6940
rect 13180 6700 13360 6940
rect 11760 6670 13360 6700
rect 1540 6640 3140 6670
rect 17610 2500 21610 6760
rect 22420 2600 22900 2630
rect 22420 2500 22480 2600
rect 17610 2360 22480 2500
rect 22850 2500 22900 2600
rect 26900 2600 27380 2630
rect 26900 2500 26960 2600
rect 22850 2360 26960 2500
rect 27330 2360 27380 2600
rect 17610 2100 27380 2360
rect 1080 -790 2680 -760
rect 1080 -1030 1260 -790
rect 1500 -1030 1590 -790
rect 1830 -1030 1930 -790
rect 2170 -1030 2260 -790
rect 2500 -1030 2680 -790
rect 1080 -1040 2680 -1030
rect 12220 -790 13820 -760
rect 12220 -1030 12400 -790
rect 12640 -1030 12730 -790
rect 12970 -1030 13070 -790
rect 13310 -1030 13400 -790
rect 13640 -1030 13820 -790
rect 12220 -1040 13820 -1030
rect 17610 -1040 21610 2100
rect 28580 1440 29270 7100
rect 22080 1040 29270 1440
rect 31100 7830 38500 7910
rect 31100 7590 31180 7830
rect 31420 7590 31510 7830
rect 31750 7590 31840 7830
rect 32080 7590 32170 7830
rect 32410 7590 32500 7830
rect 32740 7590 32830 7830
rect 33070 7590 33160 7830
rect 33400 7590 33490 7830
rect 33730 7590 33820 7830
rect 34060 7590 34150 7830
rect 34390 7590 34480 7830
rect 34720 7590 34810 7830
rect 35050 7590 35140 7830
rect 35380 7590 35470 7830
rect 35710 7590 35800 7830
rect 36040 7590 36130 7830
rect 36370 7590 36460 7830
rect 36700 7590 36790 7830
rect 37030 7590 37120 7830
rect 37360 7590 37450 7830
rect 37690 7770 38500 7830
rect 37690 7590 38230 7770
rect 31100 7530 38230 7590
rect 38470 7530 38500 7770
rect 31100 7500 38500 7530
rect 31100 7260 31180 7500
rect 31420 7260 31510 7500
rect 31750 7260 31840 7500
rect 32080 7260 32170 7500
rect 32410 7260 32500 7500
rect 32740 7260 32830 7500
rect 33070 7260 33160 7500
rect 33400 7260 33490 7500
rect 33730 7260 33820 7500
rect 34060 7260 34150 7500
rect 34390 7260 34480 7500
rect 34720 7260 34810 7500
rect 35050 7260 35140 7500
rect 35380 7260 35470 7500
rect 35710 7260 35800 7500
rect 36040 7260 36130 7500
rect 36370 7260 36460 7500
rect 36700 7260 36790 7500
rect 37030 7260 37120 7500
rect 37360 7260 37450 7500
rect 37690 7440 38500 7500
rect 37690 7260 38230 7440
rect 31100 7200 38230 7260
rect 38470 7200 38500 7440
rect 31100 7170 38500 7200
rect 31100 6930 31180 7170
rect 31420 6930 31510 7170
rect 31750 6930 31840 7170
rect 32080 6930 32170 7170
rect 32410 6930 32500 7170
rect 32740 6930 32830 7170
rect 33070 6930 33160 7170
rect 33400 6930 33490 7170
rect 33730 6930 33820 7170
rect 34060 6930 34150 7170
rect 34390 6930 34480 7170
rect 34720 6930 34810 7170
rect 35050 6930 35140 7170
rect 35380 6930 35470 7170
rect 35710 6930 35800 7170
rect 36040 6930 36130 7170
rect 36370 6930 36460 7170
rect 36700 6930 36790 7170
rect 37030 6930 37120 7170
rect 37360 6930 37450 7170
rect 37690 7070 38500 7170
rect 37690 6930 38230 7070
rect 31100 6840 38230 6930
rect 31100 6600 31180 6840
rect 31420 6600 31510 6840
rect 31750 6600 31840 6840
rect 32080 6600 32170 6840
rect 32410 6600 32500 6840
rect 32740 6600 32830 6840
rect 33070 6600 33160 6840
rect 33400 6600 33490 6840
rect 33730 6600 33820 6840
rect 34060 6600 34150 6840
rect 34390 6600 34480 6840
rect 34720 6600 34810 6840
rect 35050 6600 35140 6840
rect 35380 6600 35470 6840
rect 35710 6600 35800 6840
rect 36040 6600 36130 6840
rect 36370 6600 36460 6840
rect 36700 6600 36790 6840
rect 37030 6600 37120 6840
rect 37360 6600 37450 6840
rect 37690 6830 38230 6840
rect 38470 6830 38500 7070
rect 37690 6740 38500 6830
rect 37690 6600 38230 6740
rect 31100 6510 38230 6600
rect 31100 6270 31180 6510
rect 31420 6270 31510 6510
rect 31750 6270 31840 6510
rect 32080 6270 32170 6510
rect 32410 6270 32500 6510
rect 32740 6270 32830 6510
rect 33070 6270 33160 6510
rect 33400 6270 33490 6510
rect 33730 6270 33820 6510
rect 34060 6270 34150 6510
rect 34390 6270 34480 6510
rect 34720 6270 34810 6510
rect 35050 6270 35140 6510
rect 35380 6270 35470 6510
rect 35710 6270 35800 6510
rect 36040 6270 36130 6510
rect 36370 6270 36460 6510
rect 36700 6270 36790 6510
rect 37030 6270 37120 6510
rect 37360 6270 37450 6510
rect 37690 6500 38230 6510
rect 38470 6500 38500 6740
rect 37690 6410 38500 6500
rect 37690 6270 38230 6410
rect 31100 6180 38230 6270
rect 31100 5940 31180 6180
rect 31420 5940 31510 6180
rect 31750 5940 31840 6180
rect 32080 5940 32170 6180
rect 32410 5940 32500 6180
rect 32740 5940 32830 6180
rect 33070 5940 33160 6180
rect 33400 5940 33490 6180
rect 33730 5940 33820 6180
rect 34060 5940 34150 6180
rect 34390 5940 34480 6180
rect 34720 5940 34810 6180
rect 35050 5940 35140 6180
rect 35380 5940 35470 6180
rect 35710 5940 35800 6180
rect 36040 5940 36130 6180
rect 36370 5940 36460 6180
rect 36700 5940 36790 6180
rect 37030 5940 37120 6180
rect 37360 5940 37450 6180
rect 37690 6170 38230 6180
rect 38470 6170 38500 6410
rect 37690 6080 38500 6170
rect 37690 5940 38230 6080
rect 31100 5850 38230 5940
rect 31100 5610 31180 5850
rect 31420 5610 31510 5850
rect 31750 5610 31840 5850
rect 32080 5610 32170 5850
rect 32410 5610 32500 5850
rect 32740 5610 32830 5850
rect 33070 5610 33160 5850
rect 33400 5610 33490 5850
rect 33730 5610 33820 5850
rect 34060 5610 34150 5850
rect 34390 5610 34480 5850
rect 34720 5610 34810 5850
rect 35050 5610 35140 5850
rect 35380 5610 35470 5850
rect 35710 5610 35800 5850
rect 36040 5610 36130 5850
rect 36370 5610 36460 5850
rect 36700 5610 36790 5850
rect 37030 5610 37120 5850
rect 37360 5610 37450 5850
rect 37690 5840 38230 5850
rect 38470 5840 38500 6080
rect 37690 5750 38500 5840
rect 37690 5610 38230 5750
rect 31100 5520 38230 5610
rect 31100 5280 31180 5520
rect 31420 5280 31510 5520
rect 31750 5280 31840 5520
rect 32080 5280 32170 5520
rect 32410 5280 32500 5520
rect 32740 5280 32830 5520
rect 33070 5280 33160 5520
rect 33400 5280 33490 5520
rect 33730 5280 33820 5520
rect 34060 5280 34150 5520
rect 34390 5280 34480 5520
rect 34720 5280 34810 5520
rect 35050 5280 35140 5520
rect 35380 5280 35470 5520
rect 35710 5280 35800 5520
rect 36040 5280 36130 5520
rect 36370 5280 36460 5520
rect 36700 5280 36790 5520
rect 37030 5280 37120 5520
rect 37360 5280 37450 5520
rect 37690 5510 38230 5520
rect 38470 5510 38500 5750
rect 37690 5420 38500 5510
rect 37690 5280 38230 5420
rect 31100 5190 38230 5280
rect 31100 4950 31180 5190
rect 31420 4950 31510 5190
rect 31750 4950 31840 5190
rect 32080 4950 32170 5190
rect 32410 4950 32500 5190
rect 32740 4950 32830 5190
rect 33070 4950 33160 5190
rect 33400 4950 33490 5190
rect 33730 4950 33820 5190
rect 34060 4950 34150 5190
rect 34390 4950 34480 5190
rect 34720 4950 34810 5190
rect 35050 4950 35140 5190
rect 35380 4950 35470 5190
rect 35710 4950 35800 5190
rect 36040 4950 36130 5190
rect 36370 4950 36460 5190
rect 36700 4950 36790 5190
rect 37030 4950 37120 5190
rect 37360 4950 37450 5190
rect 37690 5180 38230 5190
rect 38470 5180 38500 5420
rect 37690 5090 38500 5180
rect 37690 4950 38230 5090
rect 31100 4860 38230 4950
rect 31100 4620 31180 4860
rect 31420 4620 31510 4860
rect 31750 4620 31840 4860
rect 32080 4620 32170 4860
rect 32410 4620 32500 4860
rect 32740 4620 32830 4860
rect 33070 4620 33160 4860
rect 33400 4620 33490 4860
rect 33730 4620 33820 4860
rect 34060 4620 34150 4860
rect 34390 4620 34480 4860
rect 34720 4620 34810 4860
rect 35050 4620 35140 4860
rect 35380 4620 35470 4860
rect 35710 4620 35800 4860
rect 36040 4620 36130 4860
rect 36370 4620 36460 4860
rect 36700 4620 36790 4860
rect 37030 4620 37120 4860
rect 37360 4620 37450 4860
rect 37690 4850 38230 4860
rect 38470 4850 38500 5090
rect 37690 4760 38500 4850
rect 37690 4620 38230 4760
rect 31100 4530 38230 4620
rect 31100 4290 31180 4530
rect 31420 4290 31510 4530
rect 31750 4290 31840 4530
rect 32080 4290 32170 4530
rect 32410 4290 32500 4530
rect 32740 4290 32830 4530
rect 33070 4290 33160 4530
rect 33400 4290 33490 4530
rect 33730 4290 33820 4530
rect 34060 4290 34150 4530
rect 34390 4290 34480 4530
rect 34720 4290 34810 4530
rect 35050 4290 35140 4530
rect 35380 4290 35470 4530
rect 35710 4290 35800 4530
rect 36040 4290 36130 4530
rect 36370 4290 36460 4530
rect 36700 4290 36790 4530
rect 37030 4290 37120 4530
rect 37360 4290 37450 4530
rect 37690 4520 38230 4530
rect 38470 4520 38500 4760
rect 37690 4430 38500 4520
rect 37690 4290 38230 4430
rect 31100 4200 38230 4290
rect 31100 3960 31180 4200
rect 31420 3960 31510 4200
rect 31750 3960 31840 4200
rect 32080 3960 32170 4200
rect 32410 3960 32500 4200
rect 32740 3960 32830 4200
rect 33070 3960 33160 4200
rect 33400 3960 33490 4200
rect 33730 3960 33820 4200
rect 34060 3960 34150 4200
rect 34390 3960 34480 4200
rect 34720 3960 34810 4200
rect 35050 3960 35140 4200
rect 35380 3960 35470 4200
rect 35710 3960 35800 4200
rect 36040 3960 36130 4200
rect 36370 3960 36460 4200
rect 36700 3960 36790 4200
rect 37030 3960 37120 4200
rect 37360 3960 37450 4200
rect 37690 4190 38230 4200
rect 38470 4190 38500 4430
rect 37690 4060 38500 4190
rect 37690 3960 38230 4060
rect 31100 3870 38230 3960
rect 31100 3630 31180 3870
rect 31420 3630 31510 3870
rect 31750 3630 31840 3870
rect 32080 3630 32170 3870
rect 32410 3630 32500 3870
rect 32740 3630 32830 3870
rect 33070 3630 33160 3870
rect 33400 3630 33490 3870
rect 33730 3630 33820 3870
rect 34060 3630 34150 3870
rect 34390 3630 34480 3870
rect 34720 3630 34810 3870
rect 35050 3630 35140 3870
rect 35380 3630 35470 3870
rect 35710 3630 35800 3870
rect 36040 3630 36130 3870
rect 36370 3630 36460 3870
rect 36700 3630 36790 3870
rect 37030 3630 37120 3870
rect 37360 3630 37450 3870
rect 37690 3820 38230 3870
rect 38470 3820 38500 4060
rect 37690 3730 38500 3820
rect 37690 3630 38230 3730
rect 31100 3540 38230 3630
rect 31100 3300 31180 3540
rect 31420 3300 31510 3540
rect 31750 3300 31840 3540
rect 32080 3300 32170 3540
rect 32410 3300 32500 3540
rect 32740 3300 32830 3540
rect 33070 3300 33160 3540
rect 33400 3300 33490 3540
rect 33730 3300 33820 3540
rect 34060 3300 34150 3540
rect 34390 3300 34480 3540
rect 34720 3300 34810 3540
rect 35050 3300 35140 3540
rect 35380 3300 35470 3540
rect 35710 3300 35800 3540
rect 36040 3300 36130 3540
rect 36370 3300 36460 3540
rect 36700 3300 36790 3540
rect 37030 3300 37120 3540
rect 37360 3300 37450 3540
rect 37690 3490 38230 3540
rect 38470 3490 38500 3730
rect 37690 3400 38500 3490
rect 37690 3300 38230 3400
rect 31100 3210 38230 3300
rect 31100 2970 31180 3210
rect 31420 2970 31510 3210
rect 31750 2970 31840 3210
rect 32080 2970 32170 3210
rect 32410 2970 32500 3210
rect 32740 2970 32830 3210
rect 33070 2970 33160 3210
rect 33400 2970 33490 3210
rect 33730 2970 33820 3210
rect 34060 2970 34150 3210
rect 34390 2970 34480 3210
rect 34720 2970 34810 3210
rect 35050 2970 35140 3210
rect 35380 2970 35470 3210
rect 35710 2970 35800 3210
rect 36040 2970 36130 3210
rect 36370 2970 36460 3210
rect 36700 2970 36790 3210
rect 37030 2970 37120 3210
rect 37360 2970 37450 3210
rect 37690 3160 38230 3210
rect 38470 3160 38500 3400
rect 37690 3070 38500 3160
rect 37690 2970 38230 3070
rect 31100 2880 38230 2970
rect 31100 2640 31180 2880
rect 31420 2640 31510 2880
rect 31750 2640 31840 2880
rect 32080 2640 32170 2880
rect 32410 2640 32500 2880
rect 32740 2640 32830 2880
rect 33070 2640 33160 2880
rect 33400 2640 33490 2880
rect 33730 2640 33820 2880
rect 34060 2640 34150 2880
rect 34390 2640 34480 2880
rect 34720 2640 34810 2880
rect 35050 2640 35140 2880
rect 35380 2640 35470 2880
rect 35710 2640 35800 2880
rect 36040 2640 36130 2880
rect 36370 2640 36460 2880
rect 36700 2640 36790 2880
rect 37030 2640 37120 2880
rect 37360 2640 37450 2880
rect 37690 2830 38230 2880
rect 38470 2830 38500 3070
rect 37690 2740 38500 2830
rect 37690 2640 38230 2740
rect 31100 2550 38230 2640
rect 31100 2310 31180 2550
rect 31420 2310 31510 2550
rect 31750 2310 31840 2550
rect 32080 2310 32170 2550
rect 32410 2310 32500 2550
rect 32740 2310 32830 2550
rect 33070 2310 33160 2550
rect 33400 2310 33490 2550
rect 33730 2310 33820 2550
rect 34060 2310 34150 2550
rect 34390 2310 34480 2550
rect 34720 2310 34810 2550
rect 35050 2310 35140 2550
rect 35380 2310 35470 2550
rect 35710 2310 35800 2550
rect 36040 2310 36130 2550
rect 36370 2310 36460 2550
rect 36700 2310 36790 2550
rect 37030 2310 37120 2550
rect 37360 2310 37450 2550
rect 37690 2500 38230 2550
rect 38470 2500 38500 2740
rect 37690 2410 38500 2500
rect 37690 2310 38230 2410
rect 31100 2220 38230 2310
rect 31100 1980 31180 2220
rect 31420 1980 31510 2220
rect 31750 1980 31840 2220
rect 32080 1980 32170 2220
rect 32410 1980 32500 2220
rect 32740 1980 32830 2220
rect 33070 1980 33160 2220
rect 33400 1980 33490 2220
rect 33730 1980 33820 2220
rect 34060 1980 34150 2220
rect 34390 1980 34480 2220
rect 34720 1980 34810 2220
rect 35050 1980 35140 2220
rect 35380 1980 35470 2220
rect 35710 1980 35800 2220
rect 36040 1980 36130 2220
rect 36370 1980 36460 2220
rect 36700 1980 36790 2220
rect 37030 1980 37120 2220
rect 37360 1980 37450 2220
rect 37690 2170 38230 2220
rect 38470 2170 38500 2410
rect 37690 2080 38500 2170
rect 37690 1980 38230 2080
rect 31100 1890 38230 1980
rect 31100 1650 31180 1890
rect 31420 1650 31510 1890
rect 31750 1650 31840 1890
rect 32080 1650 32170 1890
rect 32410 1650 32500 1890
rect 32740 1650 32830 1890
rect 33070 1650 33160 1890
rect 33400 1650 33490 1890
rect 33730 1650 33820 1890
rect 34060 1650 34150 1890
rect 34390 1650 34480 1890
rect 34720 1650 34810 1890
rect 35050 1650 35140 1890
rect 35380 1650 35470 1890
rect 35710 1650 35800 1890
rect 36040 1650 36130 1890
rect 36370 1650 36460 1890
rect 36700 1650 36790 1890
rect 37030 1650 37120 1890
rect 37360 1650 37450 1890
rect 37690 1840 38230 1890
rect 38470 1840 38500 2080
rect 37690 1750 38500 1840
rect 37690 1650 38230 1750
rect 31100 1560 38230 1650
rect 31100 1320 31180 1560
rect 31420 1320 31510 1560
rect 31750 1320 31840 1560
rect 32080 1320 32170 1560
rect 32410 1320 32500 1560
rect 32740 1320 32830 1560
rect 33070 1320 33160 1560
rect 33400 1320 33490 1560
rect 33730 1320 33820 1560
rect 34060 1320 34150 1560
rect 34390 1320 34480 1560
rect 34720 1320 34810 1560
rect 35050 1320 35140 1560
rect 35380 1320 35470 1560
rect 35710 1320 35800 1560
rect 36040 1320 36130 1560
rect 36370 1320 36460 1560
rect 36700 1320 36790 1560
rect 37030 1320 37120 1560
rect 37360 1320 37450 1560
rect 37690 1510 38230 1560
rect 38470 1510 38500 1750
rect 37690 1420 38500 1510
rect 37690 1320 38230 1420
rect 31100 1180 38230 1320
rect 38470 1180 38500 1420
rect 23460 980 23940 1040
rect 23460 740 23510 980
rect 23880 740 23940 980
rect 23460 710 23940 740
rect 25860 980 26340 1040
rect 25860 740 25910 980
rect 26280 740 26340 980
rect 25860 710 26340 740
rect -170 -1840 21610 -1040
rect -6530 -2720 14530 -2160
rect -6530 -2960 1720 -2720
rect 1960 -2960 2050 -2720
rect 2290 -2960 2390 -2720
rect 2630 -2960 2720 -2720
rect 2960 -2960 11940 -2720
rect 12180 -2960 12270 -2720
rect 12510 -2960 12610 -2720
rect 12850 -2960 12940 -2720
rect 13180 -2960 14530 -2720
rect -6530 -11680 -2530 -2960
rect 1540 -2990 3140 -2960
rect 11760 -2990 13360 -2960
rect 17610 -3840 21610 -1840
rect 31100 230 38500 1180
rect 31100 -10 31180 230
rect 31420 -10 31510 230
rect 31750 -10 31840 230
rect 32080 -10 32170 230
rect 32410 -10 32500 230
rect 32740 -10 32830 230
rect 33070 -10 33160 230
rect 33400 -10 33490 230
rect 33730 -10 33820 230
rect 34060 -10 34150 230
rect 34390 -10 34480 230
rect 34720 -10 34810 230
rect 35050 -10 35140 230
rect 35380 -10 35470 230
rect 35710 -10 35800 230
rect 36040 -10 36130 230
rect 36370 -10 36460 230
rect 36700 -10 36790 230
rect 37030 -10 37120 230
rect 37360 -10 37450 230
rect 37690 170 38500 230
rect 37690 -10 38230 170
rect 31100 -70 38230 -10
rect 38470 -70 38500 170
rect 31100 -100 38500 -70
rect 31100 -340 31180 -100
rect 31420 -340 31510 -100
rect 31750 -340 31840 -100
rect 32080 -340 32170 -100
rect 32410 -340 32500 -100
rect 32740 -340 32830 -100
rect 33070 -340 33160 -100
rect 33400 -340 33490 -100
rect 33730 -340 33820 -100
rect 34060 -340 34150 -100
rect 34390 -340 34480 -100
rect 34720 -340 34810 -100
rect 35050 -340 35140 -100
rect 35380 -340 35470 -100
rect 35710 -340 35800 -100
rect 36040 -340 36130 -100
rect 36370 -340 36460 -100
rect 36700 -340 36790 -100
rect 37030 -340 37120 -100
rect 37360 -340 37450 -100
rect 37690 -160 38500 -100
rect 37690 -340 38230 -160
rect 31100 -400 38230 -340
rect 38470 -400 38500 -160
rect 31100 -430 38500 -400
rect 31100 -670 31180 -430
rect 31420 -670 31510 -430
rect 31750 -670 31840 -430
rect 32080 -670 32170 -430
rect 32410 -670 32500 -430
rect 32740 -670 32830 -430
rect 33070 -670 33160 -430
rect 33400 -670 33490 -430
rect 33730 -670 33820 -430
rect 34060 -670 34150 -430
rect 34390 -670 34480 -430
rect 34720 -670 34810 -430
rect 35050 -670 35140 -430
rect 35380 -670 35470 -430
rect 35710 -670 35800 -430
rect 36040 -670 36130 -430
rect 36370 -670 36460 -430
rect 36700 -670 36790 -430
rect 37030 -670 37120 -430
rect 37360 -670 37450 -430
rect 37690 -530 38500 -430
rect 37690 -670 38230 -530
rect 31100 -760 38230 -670
rect 31100 -1000 31180 -760
rect 31420 -1000 31510 -760
rect 31750 -1000 31840 -760
rect 32080 -1000 32170 -760
rect 32410 -1000 32500 -760
rect 32740 -1000 32830 -760
rect 33070 -1000 33160 -760
rect 33400 -1000 33490 -760
rect 33730 -1000 33820 -760
rect 34060 -1000 34150 -760
rect 34390 -1000 34480 -760
rect 34720 -1000 34810 -760
rect 35050 -1000 35140 -760
rect 35380 -1000 35470 -760
rect 35710 -1000 35800 -760
rect 36040 -1000 36130 -760
rect 36370 -1000 36460 -760
rect 36700 -1000 36790 -760
rect 37030 -1000 37120 -760
rect 37360 -1000 37450 -760
rect 37690 -770 38230 -760
rect 38470 -770 38500 -530
rect 37690 -860 38500 -770
rect 37690 -1000 38230 -860
rect 31100 -1090 38230 -1000
rect 31100 -1330 31180 -1090
rect 31420 -1330 31510 -1090
rect 31750 -1330 31840 -1090
rect 32080 -1330 32170 -1090
rect 32410 -1330 32500 -1090
rect 32740 -1330 32830 -1090
rect 33070 -1330 33160 -1090
rect 33400 -1330 33490 -1090
rect 33730 -1330 33820 -1090
rect 34060 -1330 34150 -1090
rect 34390 -1330 34480 -1090
rect 34720 -1330 34810 -1090
rect 35050 -1330 35140 -1090
rect 35380 -1330 35470 -1090
rect 35710 -1330 35800 -1090
rect 36040 -1330 36130 -1090
rect 36370 -1330 36460 -1090
rect 36700 -1330 36790 -1090
rect 37030 -1330 37120 -1090
rect 37360 -1330 37450 -1090
rect 37690 -1100 38230 -1090
rect 38470 -1100 38500 -860
rect 37690 -1190 38500 -1100
rect 37690 -1330 38230 -1190
rect 31100 -1420 38230 -1330
rect 31100 -1660 31180 -1420
rect 31420 -1660 31510 -1420
rect 31750 -1660 31840 -1420
rect 32080 -1660 32170 -1420
rect 32410 -1660 32500 -1420
rect 32740 -1660 32830 -1420
rect 33070 -1660 33160 -1420
rect 33400 -1660 33490 -1420
rect 33730 -1660 33820 -1420
rect 34060 -1660 34150 -1420
rect 34390 -1660 34480 -1420
rect 34720 -1660 34810 -1420
rect 35050 -1660 35140 -1420
rect 35380 -1660 35470 -1420
rect 35710 -1660 35800 -1420
rect 36040 -1660 36130 -1420
rect 36370 -1660 36460 -1420
rect 36700 -1660 36790 -1420
rect 37030 -1660 37120 -1420
rect 37360 -1660 37450 -1420
rect 37690 -1430 38230 -1420
rect 38470 -1430 38500 -1190
rect 37690 -1520 38500 -1430
rect 37690 -1660 38230 -1520
rect 31100 -1750 38230 -1660
rect 31100 -1990 31180 -1750
rect 31420 -1990 31510 -1750
rect 31750 -1990 31840 -1750
rect 32080 -1990 32170 -1750
rect 32410 -1990 32500 -1750
rect 32740 -1990 32830 -1750
rect 33070 -1990 33160 -1750
rect 33400 -1990 33490 -1750
rect 33730 -1990 33820 -1750
rect 34060 -1990 34150 -1750
rect 34390 -1990 34480 -1750
rect 34720 -1990 34810 -1750
rect 35050 -1990 35140 -1750
rect 35380 -1990 35470 -1750
rect 35710 -1990 35800 -1750
rect 36040 -1990 36130 -1750
rect 36370 -1990 36460 -1750
rect 36700 -1990 36790 -1750
rect 37030 -1990 37120 -1750
rect 37360 -1990 37450 -1750
rect 37690 -1760 38230 -1750
rect 38470 -1760 38500 -1520
rect 37690 -1850 38500 -1760
rect 37690 -1990 38230 -1850
rect 31100 -2080 38230 -1990
rect 31100 -2320 31180 -2080
rect 31420 -2320 31510 -2080
rect 31750 -2320 31840 -2080
rect 32080 -2320 32170 -2080
rect 32410 -2320 32500 -2080
rect 32740 -2320 32830 -2080
rect 33070 -2320 33160 -2080
rect 33400 -2320 33490 -2080
rect 33730 -2320 33820 -2080
rect 34060 -2320 34150 -2080
rect 34390 -2320 34480 -2080
rect 34720 -2320 34810 -2080
rect 35050 -2320 35140 -2080
rect 35380 -2320 35470 -2080
rect 35710 -2320 35800 -2080
rect 36040 -2320 36130 -2080
rect 36370 -2320 36460 -2080
rect 36700 -2320 36790 -2080
rect 37030 -2320 37120 -2080
rect 37360 -2320 37450 -2080
rect 37690 -2090 38230 -2080
rect 38470 -2090 38500 -1850
rect 37690 -2180 38500 -2090
rect 37690 -2320 38230 -2180
rect 31100 -2410 38230 -2320
rect 31100 -2650 31180 -2410
rect 31420 -2650 31510 -2410
rect 31750 -2650 31840 -2410
rect 32080 -2650 32170 -2410
rect 32410 -2650 32500 -2410
rect 32740 -2650 32830 -2410
rect 33070 -2650 33160 -2410
rect 33400 -2650 33490 -2410
rect 33730 -2650 33820 -2410
rect 34060 -2650 34150 -2410
rect 34390 -2650 34480 -2410
rect 34720 -2650 34810 -2410
rect 35050 -2650 35140 -2410
rect 35380 -2650 35470 -2410
rect 35710 -2650 35800 -2410
rect 36040 -2650 36130 -2410
rect 36370 -2650 36460 -2410
rect 36700 -2650 36790 -2410
rect 37030 -2650 37120 -2410
rect 37360 -2650 37450 -2410
rect 37690 -2420 38230 -2410
rect 38470 -2420 38500 -2180
rect 37690 -2510 38500 -2420
rect 37690 -2650 38230 -2510
rect 31100 -2740 38230 -2650
rect 31100 -2980 31180 -2740
rect 31420 -2980 31510 -2740
rect 31750 -2980 31840 -2740
rect 32080 -2980 32170 -2740
rect 32410 -2980 32500 -2740
rect 32740 -2980 32830 -2740
rect 33070 -2980 33160 -2740
rect 33400 -2980 33490 -2740
rect 33730 -2980 33820 -2740
rect 34060 -2980 34150 -2740
rect 34390 -2980 34480 -2740
rect 34720 -2980 34810 -2740
rect 35050 -2980 35140 -2740
rect 35380 -2980 35470 -2740
rect 35710 -2980 35800 -2740
rect 36040 -2980 36130 -2740
rect 36370 -2980 36460 -2740
rect 36700 -2980 36790 -2740
rect 37030 -2980 37120 -2740
rect 37360 -2980 37450 -2740
rect 37690 -2750 38230 -2740
rect 38470 -2750 38500 -2510
rect 37690 -2840 38500 -2750
rect 37690 -2980 38230 -2840
rect 31100 -3070 38230 -2980
rect 31100 -3310 31180 -3070
rect 31420 -3310 31510 -3070
rect 31750 -3310 31840 -3070
rect 32080 -3310 32170 -3070
rect 32410 -3310 32500 -3070
rect 32740 -3310 32830 -3070
rect 33070 -3310 33160 -3070
rect 33400 -3310 33490 -3070
rect 33730 -3310 33820 -3070
rect 34060 -3310 34150 -3070
rect 34390 -3310 34480 -3070
rect 34720 -3310 34810 -3070
rect 35050 -3310 35140 -3070
rect 35380 -3310 35470 -3070
rect 35710 -3310 35800 -3070
rect 36040 -3310 36130 -3070
rect 36370 -3310 36460 -3070
rect 36700 -3310 36790 -3070
rect 37030 -3310 37120 -3070
rect 37360 -3310 37450 -3070
rect 37690 -3080 38230 -3070
rect 38470 -3080 38500 -2840
rect 37690 -3170 38500 -3080
rect 37690 -3310 38230 -3170
rect 31100 -3400 38230 -3310
rect 31100 -3640 31180 -3400
rect 31420 -3640 31510 -3400
rect 31750 -3640 31840 -3400
rect 32080 -3640 32170 -3400
rect 32410 -3640 32500 -3400
rect 32740 -3640 32830 -3400
rect 33070 -3640 33160 -3400
rect 33400 -3640 33490 -3400
rect 33730 -3640 33820 -3400
rect 34060 -3640 34150 -3400
rect 34390 -3640 34480 -3400
rect 34720 -3640 34810 -3400
rect 35050 -3640 35140 -3400
rect 35380 -3640 35470 -3400
rect 35710 -3640 35800 -3400
rect 36040 -3640 36130 -3400
rect 36370 -3640 36460 -3400
rect 36700 -3640 36790 -3400
rect 37030 -3640 37120 -3400
rect 37360 -3640 37450 -3400
rect 37690 -3410 38230 -3400
rect 38470 -3410 38500 -3170
rect 37690 -3540 38500 -3410
rect 37690 -3640 38230 -3540
rect 22420 -3690 22900 -3660
rect 22420 -3840 22480 -3690
rect 17610 -3930 22480 -3840
rect 22850 -3840 22900 -3690
rect 26900 -3690 27380 -3660
rect 26900 -3840 26960 -3690
rect 22850 -3930 26960 -3840
rect 27330 -3840 27380 -3690
rect 31100 -3730 38230 -3640
rect 31100 -3840 31180 -3730
rect 27330 -3850 29220 -3840
rect 30380 -3850 31180 -3840
rect 27330 -3930 31180 -3850
rect 17610 -3970 31180 -3930
rect 31420 -3970 31510 -3730
rect 31750 -3970 31840 -3730
rect 32080 -3970 32170 -3730
rect 32410 -3970 32500 -3730
rect 32740 -3970 32830 -3730
rect 33070 -3970 33160 -3730
rect 33400 -3970 33490 -3730
rect 33730 -3970 33820 -3730
rect 34060 -3970 34150 -3730
rect 34390 -3970 34480 -3730
rect 34720 -3970 34810 -3730
rect 35050 -3970 35140 -3730
rect 35380 -3970 35470 -3730
rect 35710 -3970 35800 -3730
rect 36040 -3970 36130 -3730
rect 36370 -3970 36460 -3730
rect 36700 -3970 36790 -3730
rect 37030 -3970 37120 -3730
rect 37360 -3970 37450 -3730
rect 37690 -3780 38230 -3730
rect 38470 -3780 38500 -3540
rect 37690 -3870 38500 -3780
rect 37690 -3970 38230 -3870
rect 17610 -4060 38230 -3970
rect 17610 -4240 31180 -4060
rect -1350 -4840 260 -4630
rect -1350 -5080 -1180 -4840
rect -940 -5080 -850 -4840
rect -610 -5080 -520 -4840
rect -280 -5080 -190 -4840
rect 50 -5080 260 -4840
rect -1350 -5170 260 -5080
rect -1350 -5410 -1180 -5170
rect -940 -5410 -850 -5170
rect -610 -5410 -520 -5170
rect -280 -5410 -190 -5170
rect 50 -5410 260 -5170
rect -1350 -5500 260 -5410
rect -1350 -5740 -1180 -5500
rect -940 -5740 -850 -5500
rect -610 -5740 -520 -5500
rect -280 -5740 -190 -5500
rect 50 -5740 260 -5500
rect -1350 -5830 260 -5740
rect -1350 -6070 -1180 -5830
rect -940 -6070 -850 -5830
rect -610 -6070 -520 -5830
rect -280 -6070 -190 -5830
rect 50 -6070 260 -5830
rect -1350 -6370 260 -6070
rect -1350 -6610 -1170 -6370
rect -930 -6610 -840 -6370
rect -600 -6610 -510 -6370
rect -270 -6610 -180 -6370
rect 60 -6610 260 -6370
rect -1350 -6640 260 -6610
rect 14520 -4840 16130 -4630
rect 14520 -5080 14730 -4840
rect 14970 -5080 15060 -4840
rect 15300 -5080 15390 -4840
rect 15630 -5080 15720 -4840
rect 15960 -5080 16130 -4840
rect 14520 -5170 16130 -5080
rect 14520 -5410 14730 -5170
rect 14970 -5410 15060 -5170
rect 15300 -5410 15390 -5170
rect 15630 -5410 15720 -5170
rect 15960 -5410 16130 -5170
rect 14520 -5500 16130 -5410
rect 14520 -5740 14730 -5500
rect 14970 -5740 15060 -5500
rect 15300 -5740 15390 -5500
rect 15630 -5740 15720 -5500
rect 15960 -5740 16130 -5500
rect 14520 -5830 16130 -5740
rect 14520 -6070 14730 -5830
rect 14970 -6070 15060 -5830
rect 15300 -6070 15390 -5830
rect 15630 -6070 15720 -5830
rect 15960 -6070 16130 -5830
rect 14520 -6370 16130 -6070
rect 14520 -6610 14720 -6370
rect 14960 -6610 15050 -6370
rect 15290 -6610 15380 -6370
rect 15620 -6610 15710 -6370
rect 15950 -6610 16130 -6370
rect 14520 -6640 16130 -6610
rect 17610 -8330 21610 -4240
rect 29220 -4250 30380 -4240
rect 31100 -4300 31180 -4240
rect 31420 -4300 31510 -4060
rect 31750 -4300 31840 -4060
rect 32080 -4300 32170 -4060
rect 32410 -4300 32500 -4060
rect 32740 -4300 32830 -4060
rect 33070 -4300 33160 -4060
rect 33400 -4300 33490 -4060
rect 33730 -4300 33820 -4060
rect 34060 -4300 34150 -4060
rect 34390 -4300 34480 -4060
rect 34720 -4300 34810 -4060
rect 35050 -4300 35140 -4060
rect 35380 -4300 35470 -4060
rect 35710 -4300 35800 -4060
rect 36040 -4300 36130 -4060
rect 36370 -4300 36460 -4060
rect 36700 -4300 36790 -4060
rect 37030 -4300 37120 -4060
rect 37360 -4300 37450 -4060
rect 37690 -4110 38230 -4060
rect 38470 -4110 38500 -3870
rect 37690 -4200 38500 -4110
rect 37690 -4300 38230 -4200
rect 31100 -4390 38230 -4300
rect 31100 -4630 31180 -4390
rect 31420 -4630 31510 -4390
rect 31750 -4630 31840 -4390
rect 32080 -4630 32170 -4390
rect 32410 -4630 32500 -4390
rect 32740 -4630 32830 -4390
rect 33070 -4630 33160 -4390
rect 33400 -4630 33490 -4390
rect 33730 -4630 33820 -4390
rect 34060 -4630 34150 -4390
rect 34390 -4630 34480 -4390
rect 34720 -4630 34810 -4390
rect 35050 -4630 35140 -4390
rect 35380 -4630 35470 -4390
rect 35710 -4630 35800 -4390
rect 36040 -4630 36130 -4390
rect 36370 -4630 36460 -4390
rect 36700 -4630 36790 -4390
rect 37030 -4630 37120 -4390
rect 37360 -4630 37450 -4390
rect 37690 -4440 38230 -4390
rect 38470 -4440 38500 -4200
rect 37690 -4530 38500 -4440
rect 37690 -4630 38230 -4530
rect 31100 -4720 38230 -4630
rect 31100 -4960 31180 -4720
rect 31420 -4960 31510 -4720
rect 31750 -4960 31840 -4720
rect 32080 -4960 32170 -4720
rect 32410 -4960 32500 -4720
rect 32740 -4960 32830 -4720
rect 33070 -4960 33160 -4720
rect 33400 -4960 33490 -4720
rect 33730 -4960 33820 -4720
rect 34060 -4960 34150 -4720
rect 34390 -4960 34480 -4720
rect 34720 -4960 34810 -4720
rect 35050 -4960 35140 -4720
rect 35380 -4960 35470 -4720
rect 35710 -4960 35800 -4720
rect 36040 -4960 36130 -4720
rect 36370 -4960 36460 -4720
rect 36700 -4960 36790 -4720
rect 37030 -4960 37120 -4720
rect 37360 -4960 37450 -4720
rect 37690 -4770 38230 -4720
rect 38470 -4770 38500 -4530
rect 37690 -4860 38500 -4770
rect 37690 -4960 38230 -4860
rect 31100 -5050 38230 -4960
rect 31100 -5290 31180 -5050
rect 31420 -5290 31510 -5050
rect 31750 -5290 31840 -5050
rect 32080 -5290 32170 -5050
rect 32410 -5290 32500 -5050
rect 32740 -5290 32830 -5050
rect 33070 -5290 33160 -5050
rect 33400 -5290 33490 -5050
rect 33730 -5290 33820 -5050
rect 34060 -5290 34150 -5050
rect 34390 -5290 34480 -5050
rect 34720 -5290 34810 -5050
rect 35050 -5290 35140 -5050
rect 35380 -5290 35470 -5050
rect 35710 -5290 35800 -5050
rect 36040 -5290 36130 -5050
rect 36370 -5290 36460 -5050
rect 36700 -5290 36790 -5050
rect 37030 -5290 37120 -5050
rect 37360 -5290 37450 -5050
rect 37690 -5100 38230 -5050
rect 38470 -5100 38500 -4860
rect 37690 -5190 38500 -5100
rect 37690 -5290 38230 -5190
rect 31100 -5380 38230 -5290
rect 31100 -5620 31180 -5380
rect 31420 -5620 31510 -5380
rect 31750 -5620 31840 -5380
rect 32080 -5620 32170 -5380
rect 32410 -5620 32500 -5380
rect 32740 -5620 32830 -5380
rect 33070 -5620 33160 -5380
rect 33400 -5620 33490 -5380
rect 33730 -5620 33820 -5380
rect 34060 -5620 34150 -5380
rect 34390 -5620 34480 -5380
rect 34720 -5620 34810 -5380
rect 35050 -5620 35140 -5380
rect 35380 -5620 35470 -5380
rect 35710 -5620 35800 -5380
rect 36040 -5620 36130 -5380
rect 36370 -5620 36460 -5380
rect 36700 -5620 36790 -5380
rect 37030 -5620 37120 -5380
rect 37360 -5620 37450 -5380
rect 37690 -5430 38230 -5380
rect 38470 -5430 38500 -5190
rect 37690 -5520 38500 -5430
rect 37690 -5620 38230 -5520
rect 31100 -5710 38230 -5620
rect 31100 -5950 31180 -5710
rect 31420 -5950 31510 -5710
rect 31750 -5950 31840 -5710
rect 32080 -5950 32170 -5710
rect 32410 -5950 32500 -5710
rect 32740 -5950 32830 -5710
rect 33070 -5950 33160 -5710
rect 33400 -5950 33490 -5710
rect 33730 -5950 33820 -5710
rect 34060 -5950 34150 -5710
rect 34390 -5950 34480 -5710
rect 34720 -5950 34810 -5710
rect 35050 -5950 35140 -5710
rect 35380 -5950 35470 -5710
rect 35710 -5950 35800 -5710
rect 36040 -5950 36130 -5710
rect 36370 -5950 36460 -5710
rect 36700 -5950 36790 -5710
rect 37030 -5950 37120 -5710
rect 37360 -5950 37450 -5710
rect 37690 -5760 38230 -5710
rect 38470 -5760 38500 -5520
rect 37690 -5850 38500 -5760
rect 37690 -5950 38230 -5850
rect 31100 -6040 38230 -5950
rect 31100 -6280 31180 -6040
rect 31420 -6280 31510 -6040
rect 31750 -6280 31840 -6040
rect 32080 -6280 32170 -6040
rect 32410 -6280 32500 -6040
rect 32740 -6280 32830 -6040
rect 33070 -6280 33160 -6040
rect 33400 -6280 33490 -6040
rect 33730 -6280 33820 -6040
rect 34060 -6280 34150 -6040
rect 34390 -6280 34480 -6040
rect 34720 -6280 34810 -6040
rect 35050 -6280 35140 -6040
rect 35380 -6280 35470 -6040
rect 35710 -6280 35800 -6040
rect 36040 -6280 36130 -6040
rect 36370 -6280 36460 -6040
rect 36700 -6280 36790 -6040
rect 37030 -6280 37120 -6040
rect 37360 -6280 37450 -6040
rect 37690 -6090 38230 -6040
rect 38470 -6090 38500 -5850
rect 37690 -6180 38500 -6090
rect 37690 -6280 38230 -6180
rect 31100 -6420 38230 -6280
rect 38470 -6420 38500 -6180
rect 31100 -6450 38500 -6420
rect 17610 -8370 21930 -8330
rect 17610 -8610 21650 -8370
rect 21890 -8610 21930 -8370
rect 17610 -8650 21930 -8610
rect 17610 -9970 21610 -8650
rect 26880 -9970 30100 -9600
rect 1080 -10340 2680 -10310
rect 1080 -10560 1260 -10340
rect 40 -10580 1260 -10560
rect 1500 -10580 1590 -10340
rect 1830 -10580 1930 -10340
rect 2170 -10580 2260 -10340
rect 2500 -10560 2680 -10340
rect 12220 -10370 13820 -10340
rect 12220 -10560 12400 -10370
rect 2500 -10580 12400 -10560
rect 40 -10610 12400 -10580
rect 12640 -10610 12730 -10370
rect 12970 -10610 13070 -10370
rect 13310 -10610 13400 -10370
rect 13640 -10560 13820 -10370
rect 17610 -10370 30100 -9970
rect 17610 -10560 21610 -10370
rect 13640 -10610 21610 -10560
rect 40 -11360 21610 -10610
rect -6530 -12240 13070 -11680
rect -6530 -12480 2390 -12240
rect 2630 -12480 2720 -12240
rect 2960 -12480 3060 -12240
rect 3300 -12480 3390 -12240
rect 3630 -12480 11270 -12240
rect 11510 -12480 11600 -12240
rect 11840 -12480 11940 -12240
rect 12180 -12480 12270 -12240
rect 12510 -12480 13070 -12240
rect 2210 -12510 3810 -12480
rect 11090 -12510 12690 -12480
rect 17610 -13990 21610 -11360
rect 17610 -14030 21930 -13990
rect 17610 -14270 21650 -14030
rect 21890 -14270 21930 -14030
rect 17610 -14310 21930 -14270
rect 17610 -15860 21610 -14310
rect 27160 -15860 30380 -15460
rect 17610 -16260 30380 -15860
rect 17610 -20070 21610 -16260
rect 17610 -20110 21930 -20070
rect 17610 -20350 21650 -20110
rect 21890 -20350 21930 -20110
rect 17610 -20390 21930 -20350
rect 17610 -21680 21610 -20390
rect 26960 -21680 30180 -21340
rect 17610 -22080 30180 -21680
rect 2210 -22660 3810 -22630
rect 2210 -22670 2390 -22660
rect -6530 -22900 2390 -22670
rect 2630 -22900 2720 -22660
rect 2960 -22900 3060 -22660
rect 3300 -22900 3390 -22660
rect 3630 -22670 3810 -22660
rect 11090 -22660 12690 -22630
rect 11090 -22670 11270 -22660
rect 3630 -22900 11270 -22670
rect 11510 -22900 11600 -22660
rect 11840 -22900 11940 -22660
rect 12180 -22900 12270 -22660
rect 12510 -22670 12690 -22660
rect 17610 -22670 21610 -22080
rect 12510 -22900 21610 -22670
rect -6530 -23700 21610 -22900
use core  core_0
timestamp 1636213402
transform 1 0 7320 0 1 2520
box -7010 -2490 7580 4060
use core  core_1
timestamp 1636213402
transform 1 0 7320 0 1 -7060
box -7010 -2490 7580 4060
use sf  sf_0
timestamp 1634767319
transform 1 0 12590 0 1 -29850
box -10660 7260 380 17300
use cmfb  cmfb_0
timestamp 1634684585
transform 1 0 25700 0 1 2690
box -3910 -30 2310 4270
use cmfb  cmfb_1
timestamp 1634684585
transform 1 0 25700 0 1 -3610
box -3910 -30 2310 4270
use mirror_1  mirror_1_0
timestamp 1635749472
transform 1 0 20860 0 1 -9070
box 840 -570 9240 3290
use mirror_4  mirror_4_0
timestamp 1635749603
transform 1 0 20940 0 1 -20790
box 760 -570 9240 3290
use mirror_3  mirror_3_0
timestamp 1635750117
transform 1 0 21140 0 1 -14930
box 560 -570 9240 3290
<< labels >>
rlabel metal1 13060 40 13060 40 1 GND
port 7 n
rlabel metal5 -2700 7440 -2700 7440 1 VDD
port 1 n
rlabel metal3 9730 -23610 9730 -23610 1 Vout_n
port 17 n
rlabel metal3 5150 -23580 5150 -23580 1 Vout_p
port 18 n
rlabel metal3 8330 2730 8330 2730 1 Vop
rlabel metal3 6540 2730 6540 2730 1 Von
rlabel metal2 7400 360 7400 360 1 Vcm1
rlabel metal3 8870 -6850 8870 -6850 1 pre_Vout_n
rlabel metal3 6040 -6890 6040 -6890 1 pre_Vout_p
rlabel metal2 7420 -9350 7420 -9350 1 Vcm2
rlabel metal2 7620 -3520 7620 -3520 1 Vcmfb2
rlabel metal2 7470 6130 7470 6130 1 Vcmfb1
rlabel metal5 29100 7420 29100 7420 1 VDD
port 1 n
rlabel metal4 7700 8530 7700 8530 1 Vinn
rlabel metal4 7160 8530 7160 8530 1 Vinp
rlabel metal5 -6360 -23210 -6360 -23210 1 GND
port 7 n
rlabel metal4 39610 8360 39610 8360 1 Vb5
port 20 n
rlabel metal4 30970 -10670 30970 -10670 1 Vb1_
port 21 n
rlabel metal4 30890 -16530 30890 -16530 1 Vb3_
port 22 n
rlabel metal4 30660 -22400 30660 -22400 1 Vb4_
port 23 n
rlabel space 7450 21850 7450 21850 1 MIDDLE_TOP
rlabel metal4 21200 8860 21200 8860 1 Vb2
port 19 n
rlabel metal5 19910 21510 19910 21510 1 Iin_n
port 26 n
rlabel metal5 -5000 21540 -5000 21540 1 Iin_p
port 25 n
<< end >>
